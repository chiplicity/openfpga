magic
tech EFS8A
magscale 1 2
timestamp 1602269862
<< locali >>
rect 9723 11169 9758 11203
rect 7291 9129 7297 9163
rect 7291 9061 7325 9129
rect 10051 8041 10057 8075
rect 10051 7973 10085 8041
rect 18647 7905 18682 7939
rect 4445 7395 4479 7497
rect 12265 7327 12299 7497
rect 12265 7293 12518 7327
rect 2329 6817 2490 6851
rect 2329 6647 2363 6817
rect 13737 5695 13771 5797
rect 10701 5015 10735 5117
rect 7757 4471 7791 4709
rect 7849 4471 7883 4641
rect 5641 4131 5675 4233
rect 19441 3655 19475 3689
rect 19349 3621 19475 3655
rect 10793 3383 10827 3485
rect 16957 3383 16991 3485
rect 4813 2295 4847 2397
rect 6101 2295 6135 2533
rect 11897 2295 11931 2465
<< viali >>
rect 1593 18377 1627 18411
rect 4629 18377 4663 18411
rect 7665 18377 7699 18411
rect 1409 18173 1443 18207
rect 1961 18173 1995 18207
rect 4445 18173 4479 18207
rect 7481 18173 7515 18207
rect 5089 18037 5123 18071
rect 8125 18037 8159 18071
rect 1593 15657 1627 15691
rect 1409 15521 1443 15555
rect 1685 14773 1719 14807
rect 19073 13345 19107 13379
rect 19257 13209 19291 13243
rect 19073 12597 19107 12631
rect 19257 11305 19291 11339
rect 9689 11169 9723 11203
rect 19073 11169 19107 11203
rect 8217 11101 8251 11135
rect 6929 10965 6963 10999
rect 9827 10965 9861 10999
rect 10103 10761 10137 10795
rect 8401 10557 8435 10591
rect 8585 10557 8619 10591
rect 10000 10557 10034 10591
rect 10425 10557 10459 10591
rect 11012 10557 11046 10591
rect 11437 10557 11471 10591
rect 12516 10557 12550 10591
rect 6929 10489 6963 10523
rect 7021 10489 7055 10523
rect 7573 10489 7607 10523
rect 8309 10489 8343 10523
rect 6561 10421 6595 10455
rect 9781 10421 9815 10455
rect 11115 10421 11149 10455
rect 12587 10421 12621 10455
rect 12909 10421 12943 10455
rect 19073 10421 19107 10455
rect 7573 10217 7607 10251
rect 6653 10149 6687 10183
rect 7205 10149 7239 10183
rect 8125 10149 8159 10183
rect 8217 10149 8251 10183
rect 9781 10149 9815 10183
rect 9873 10149 9907 10183
rect 12357 10081 12391 10115
rect 6561 10013 6595 10047
rect 8401 10013 8435 10047
rect 10425 10013 10459 10047
rect 9229 9877 9263 9911
rect 12449 9877 12483 9911
rect 4859 9673 4893 9707
rect 7021 9673 7055 9707
rect 8585 9673 8619 9707
rect 10517 9673 10551 9707
rect 12265 9673 12299 9707
rect 16773 9673 16807 9707
rect 5273 9605 5307 9639
rect 5871 9605 5905 9639
rect 11161 9605 11195 9639
rect 7665 9537 7699 9571
rect 8309 9537 8343 9571
rect 9229 9537 9263 9571
rect 12541 9537 12575 9571
rect 13461 9537 13495 9571
rect 4788 9469 4822 9503
rect 5800 9469 5834 9503
rect 10977 9469 11011 9503
rect 11529 9469 11563 9503
rect 15612 9469 15646 9503
rect 16037 9469 16071 9503
rect 16589 9469 16623 9503
rect 17233 9469 17267 9503
rect 18128 9469 18162 9503
rect 18521 9469 18555 9503
rect 19140 9469 19174 9503
rect 19533 9469 19567 9503
rect 7481 9401 7515 9435
rect 7757 9401 7791 9435
rect 9321 9401 9355 9435
rect 9873 9401 9907 9435
rect 12633 9401 12667 9435
rect 13185 9401 13219 9435
rect 6285 9333 6319 9367
rect 6561 9333 6595 9367
rect 9045 9333 9079 9367
rect 10149 9333 10183 9367
rect 14197 9333 14231 9367
rect 15715 9333 15749 9367
rect 18199 9333 18233 9367
rect 19211 9333 19245 9367
rect 7297 9129 7331 9163
rect 7849 9129 7883 9163
rect 8125 9129 8159 9163
rect 10885 9129 10919 9163
rect 14105 9129 14139 9163
rect 19257 9129 19291 9163
rect 6101 9061 6135 9095
rect 11482 9061 11516 9095
rect 12541 9061 12575 9095
rect 13093 9061 13127 9095
rect 16497 9061 16531 9095
rect 16589 9061 16623 9095
rect 1536 8993 1570 9027
rect 6009 8993 6043 9027
rect 9724 8993 9758 9027
rect 12081 8993 12115 9027
rect 15428 8993 15462 9027
rect 18004 8993 18038 9027
rect 19073 8993 19107 9027
rect 6929 8925 6963 8959
rect 11161 8925 11195 8959
rect 13001 8925 13035 8959
rect 14381 8925 14415 8959
rect 17141 8925 17175 8959
rect 1639 8857 1673 8891
rect 8861 8857 8895 8891
rect 9827 8857 9861 8891
rect 13553 8857 13587 8891
rect 6469 8789 6503 8823
rect 6837 8789 6871 8823
rect 8493 8789 8527 8823
rect 9229 8789 9263 8823
rect 10149 8789 10183 8823
rect 10517 8789 10551 8823
rect 15531 8789 15565 8823
rect 16313 8789 16347 8823
rect 18107 8789 18141 8823
rect 1593 8585 1627 8619
rect 6193 8585 6227 8619
rect 7757 8585 7791 8619
rect 13461 8585 13495 8619
rect 15393 8585 15427 8619
rect 17417 8585 17451 8619
rect 8723 8517 8757 8551
rect 11299 8517 11333 8551
rect 13093 8517 13127 8551
rect 9413 8449 9447 8483
rect 9689 8449 9723 8483
rect 10333 8449 10367 8483
rect 12541 8449 12575 8483
rect 14381 8449 14415 8483
rect 15025 8449 15059 8483
rect 16497 8449 16531 8483
rect 18153 8449 18187 8483
rect 18429 8449 18463 8483
rect 4997 8381 5031 8415
rect 5181 8381 5215 8415
rect 6837 8381 6871 8415
rect 8652 8381 8686 8415
rect 9045 8381 9079 8415
rect 11196 8381 11230 8415
rect 11621 8381 11655 8415
rect 19676 8381 19710 8415
rect 20085 8381 20119 8415
rect 5089 8313 5123 8347
rect 7158 8313 7192 8347
rect 8033 8313 8067 8347
rect 9781 8313 9815 8347
rect 10609 8313 10643 8347
rect 12633 8313 12667 8347
rect 14105 8313 14139 8347
rect 14197 8313 14231 8347
rect 16313 8313 16347 8347
rect 16589 8313 16623 8347
rect 17141 8313 17175 8347
rect 17877 8313 17911 8347
rect 18245 8313 18279 8347
rect 19763 8313 19797 8347
rect 4077 8245 4111 8279
rect 6653 8245 6687 8279
rect 8493 8245 8527 8279
rect 11069 8245 11103 8279
rect 11989 8245 12023 8279
rect 13921 8245 13955 8279
rect 15945 8245 15979 8279
rect 19165 8245 19199 8279
rect 3893 8041 3927 8075
rect 8769 8041 8803 8075
rect 10057 8041 10091 8075
rect 16221 8041 16255 8075
rect 16865 8041 16899 8075
rect 18061 8041 18095 8075
rect 5911 7973 5945 8007
rect 8170 7973 8204 8007
rect 11942 7973 11976 8007
rect 13553 7973 13587 8007
rect 15663 7973 15697 8007
rect 17233 7973 17267 8007
rect 7849 7905 7883 7939
rect 12541 7905 12575 7939
rect 13185 7905 13219 7939
rect 18613 7905 18647 7939
rect 4537 7837 4571 7871
rect 5181 7837 5215 7871
rect 5549 7837 5583 7871
rect 9689 7837 9723 7871
rect 10885 7837 10919 7871
rect 11621 7837 11655 7871
rect 13461 7837 13495 7871
rect 13737 7837 13771 7871
rect 15301 7837 15335 7871
rect 17141 7837 17175 7871
rect 17417 7837 17451 7871
rect 19625 7837 19659 7871
rect 10609 7769 10643 7803
rect 12817 7769 12851 7803
rect 4445 7701 4479 7735
rect 6469 7701 6503 7735
rect 6929 7701 6963 7735
rect 7573 7701 7607 7735
rect 9045 7701 9079 7735
rect 9413 7701 9447 7735
rect 11529 7701 11563 7735
rect 14473 7701 14507 7735
rect 16497 7701 16531 7735
rect 18751 7701 18785 7735
rect 4445 7497 4479 7531
rect 10701 7497 10735 7531
rect 12265 7497 12299 7531
rect 13001 7497 13035 7531
rect 13645 7497 13679 7531
rect 17049 7497 17083 7531
rect 17325 7497 17359 7531
rect 18245 7497 18279 7531
rect 1685 7429 1719 7463
rect 6653 7429 6687 7463
rect 4353 7361 4387 7395
rect 4445 7361 4479 7395
rect 5273 7361 5307 7395
rect 5917 7361 5951 7395
rect 15301 7361 15335 7395
rect 16129 7361 16163 7395
rect 17785 7361 17819 7395
rect 3525 7293 3559 7327
rect 3709 7293 3743 7327
rect 7481 7293 7515 7327
rect 8217 7293 8251 7327
rect 8493 7293 8527 7327
rect 8677 7293 8711 7327
rect 9781 7293 9815 7327
rect 11621 7293 11655 7327
rect 12587 7293 12621 7327
rect 13829 7293 13863 7327
rect 14289 7293 14323 7327
rect 14657 7293 14691 7327
rect 15209 7293 15243 7327
rect 18061 7293 18095 7327
rect 19165 7293 19199 7327
rect 19717 7293 19751 7327
rect 4721 7225 4755 7259
rect 5365 7225 5399 7259
rect 6285 7225 6319 7259
rect 9229 7225 9263 7259
rect 9597 7225 9631 7259
rect 10102 7225 10136 7259
rect 11989 7225 12023 7259
rect 16450 7225 16484 7259
rect 18705 7225 18739 7259
rect 2053 7157 2087 7191
rect 2421 7157 2455 7191
rect 2697 7157 2731 7191
rect 3065 7157 3099 7191
rect 5089 7157 5123 7191
rect 7389 7157 7423 7191
rect 7757 7157 7791 7191
rect 10977 7157 11011 7191
rect 13277 7157 13311 7191
rect 15669 7157 15703 7191
rect 16037 7157 16071 7191
rect 19349 7157 19383 7191
rect 4537 6953 4571 6987
rect 5089 6953 5123 6987
rect 9781 6953 9815 6987
rect 12081 6953 12115 6987
rect 14657 6953 14691 6987
rect 15117 6953 15151 6987
rect 15393 6953 15427 6987
rect 17417 6953 17451 6987
rect 8769 6885 8803 6919
rect 13921 6885 13955 6919
rect 17785 6885 17819 6919
rect 18337 6885 18371 6919
rect 1476 6817 1510 6851
rect 5273 6817 5307 6851
rect 5733 6817 5767 6851
rect 6009 6817 6043 6851
rect 6193 6817 6227 6851
rect 7481 6817 7515 6851
rect 7941 6817 7975 6851
rect 8125 6817 8159 6851
rect 8493 6817 8527 6851
rect 9505 6817 9539 6851
rect 9965 6817 9999 6851
rect 10425 6817 10459 6851
rect 10701 6817 10735 6851
rect 10885 6817 10919 6851
rect 11897 6817 11931 6851
rect 12265 6817 12299 6851
rect 12725 6817 12759 6851
rect 12909 6817 12943 6851
rect 13185 6817 13219 6851
rect 14381 6817 14415 6851
rect 15485 6817 15519 6851
rect 15761 6817 15795 6851
rect 16129 6817 16163 6851
rect 16497 6817 16531 6851
rect 19165 6817 19199 6851
rect 11437 6749 11471 6783
rect 17693 6749 17727 6783
rect 2559 6681 2593 6715
rect 6837 6681 6871 6715
rect 19349 6681 19383 6715
rect 1547 6613 1581 6647
rect 2145 6613 2179 6647
rect 2329 6613 2363 6647
rect 2881 6613 2915 6647
rect 3341 6613 3375 6647
rect 3617 6613 3651 6647
rect 4905 6613 4939 6647
rect 9045 6613 9079 6647
rect 17049 6613 17083 6647
rect 18705 6613 18739 6647
rect 1593 6409 1627 6443
rect 6975 6409 7009 6443
rect 12587 6409 12621 6443
rect 16037 6409 16071 6443
rect 17141 6409 17175 6443
rect 17509 6409 17543 6443
rect 17785 6409 17819 6443
rect 19763 6409 19797 6443
rect 7113 6341 7147 6375
rect 9505 6341 9539 6375
rect 11437 6341 11471 6375
rect 7205 6273 7239 6307
rect 8585 6273 8619 6307
rect 12909 6273 12943 6307
rect 15393 6273 15427 6307
rect 16221 6273 16255 6307
rect 18153 6273 18187 6307
rect 18797 6273 18831 6307
rect 1409 6205 1443 6239
rect 1961 6205 1995 6239
rect 2329 6205 2363 6239
rect 2548 6205 2582 6239
rect 2973 6205 3007 6239
rect 3525 6205 3559 6239
rect 4261 6205 4295 6239
rect 5365 6205 5399 6239
rect 6837 6205 6871 6239
rect 10057 6205 10091 6239
rect 10517 6205 10551 6239
rect 11069 6205 11103 6239
rect 11253 6205 11287 6239
rect 12484 6205 12518 6239
rect 13277 6205 13311 6239
rect 14013 6205 14047 6239
rect 14381 6205 14415 6239
rect 14749 6205 14783 6239
rect 15117 6205 15151 6239
rect 19692 6205 19726 6239
rect 20085 6205 20119 6239
rect 4353 6137 4387 6171
rect 4721 6137 4755 6171
rect 5917 6137 5951 6171
rect 7573 6137 7607 6171
rect 8677 6137 8711 6171
rect 9229 6137 9263 6171
rect 16542 6137 16576 6171
rect 18245 6137 18279 6171
rect 2651 6069 2685 6103
rect 5089 6069 5123 6103
rect 6285 6069 6319 6103
rect 6561 6069 6595 6103
rect 7849 6069 7883 6103
rect 8309 6069 8343 6103
rect 9873 6069 9907 6103
rect 11989 6069 12023 6103
rect 13737 6069 13771 6103
rect 15669 6069 15703 6103
rect 19165 6069 19199 6103
rect 6837 5865 6871 5899
rect 9137 5865 9171 5899
rect 11713 5865 11747 5899
rect 14749 5865 14783 5899
rect 15117 5865 15151 5899
rect 15485 5865 15519 5899
rect 16589 5865 16623 5899
rect 18429 5865 18463 5899
rect 18797 5865 18831 5899
rect 8125 5797 8159 5831
rect 8217 5797 8251 5831
rect 10241 5797 10275 5831
rect 11529 5797 11563 5831
rect 13553 5797 13587 5831
rect 13737 5797 13771 5831
rect 14013 5797 14047 5831
rect 16031 5797 16065 5831
rect 16865 5797 16899 5831
rect 17601 5797 17635 5831
rect 2237 5729 2271 5763
rect 4077 5729 4111 5763
rect 5641 5729 5675 5763
rect 6377 5729 6411 5763
rect 6469 5729 6503 5763
rect 6929 5729 6963 5763
rect 11897 5729 11931 5763
rect 12081 5729 12115 5763
rect 12541 5729 12575 5763
rect 12817 5729 12851 5763
rect 14105 5729 14139 5763
rect 18153 5729 18187 5763
rect 19073 5729 19107 5763
rect 3801 5661 3835 5695
rect 4445 5661 4479 5695
rect 10149 5661 10183 5695
rect 10793 5661 10827 5695
rect 13737 5661 13771 5695
rect 15669 5661 15703 5695
rect 17325 5661 17359 5695
rect 17509 5661 17543 5695
rect 18981 5661 19015 5695
rect 5181 5593 5215 5627
rect 7757 5593 7791 5627
rect 8677 5593 8711 5627
rect 14289 5593 14323 5627
rect 1777 5525 1811 5559
rect 2421 5525 2455 5559
rect 3525 5525 3559 5559
rect 4215 5525 4249 5559
rect 4353 5525 4387 5559
rect 4721 5525 4755 5559
rect 7481 5525 7515 5559
rect 9413 5525 9447 5559
rect 9873 5525 9907 5559
rect 11161 5525 11195 5559
rect 2605 5321 2639 5355
rect 5273 5321 5307 5355
rect 7941 5321 7975 5355
rect 10885 5321 10919 5355
rect 11621 5321 11655 5355
rect 12265 5321 12299 5355
rect 17417 5321 17451 5355
rect 19073 5321 19107 5355
rect 4813 5253 4847 5287
rect 5162 5253 5196 5287
rect 8585 5253 8619 5287
rect 13553 5253 13587 5287
rect 18705 5253 18739 5287
rect 5365 5185 5399 5219
rect 5733 5185 5767 5219
rect 15209 5185 15243 5219
rect 18153 5185 18187 5219
rect 1593 5117 1627 5151
rect 3433 5117 3467 5151
rect 7021 5117 7055 5151
rect 8217 5117 8251 5151
rect 9045 5117 9079 5151
rect 9229 5117 9263 5151
rect 9597 5117 9631 5151
rect 10149 5117 10183 5151
rect 10701 5117 10735 5151
rect 11069 5117 11103 5151
rect 12449 5117 12483 5151
rect 13737 5117 13771 5151
rect 14197 5117 14231 5151
rect 14657 5117 14691 5151
rect 15117 5117 15151 5151
rect 16037 5117 16071 5151
rect 16957 5117 16991 5151
rect 17785 5117 17819 5151
rect 2145 5049 2179 5083
rect 4997 5049 5031 5083
rect 7342 5049 7376 5083
rect 13185 5049 13219 5083
rect 16358 5049 16392 5083
rect 18245 5049 18279 5083
rect 2973 4981 3007 5015
rect 3525 4981 3559 5015
rect 4077 4981 4111 5015
rect 4445 4981 4479 5015
rect 6009 4981 6043 5015
rect 6469 4981 6503 5015
rect 9045 4981 9079 5015
rect 10609 4981 10643 5015
rect 10701 4981 10735 5015
rect 11253 4981 11287 5015
rect 12633 4981 12667 5015
rect 15485 4981 15519 5015
rect 15853 4981 15887 5015
rect 19625 4981 19659 5015
rect 1593 4777 1627 4811
rect 2237 4777 2271 4811
rect 3433 4777 3467 4811
rect 4353 4777 4387 4811
rect 5641 4777 5675 4811
rect 6469 4777 6503 4811
rect 8309 4777 8343 4811
rect 9413 4777 9447 4811
rect 10885 4777 10919 4811
rect 12081 4777 12115 4811
rect 17141 4777 17175 4811
rect 18705 4777 18739 4811
rect 2513 4709 2547 4743
rect 3065 4709 3099 4743
rect 4813 4709 4847 4743
rect 6101 4709 6135 4743
rect 7757 4709 7791 4743
rect 11482 4709 11516 4743
rect 12357 4709 12391 4743
rect 14657 4709 14691 4743
rect 15939 4709 15973 4743
rect 17509 4709 17543 4743
rect 5365 4641 5399 4675
rect 6193 4641 6227 4675
rect 6653 4641 6687 4675
rect 7021 4641 7055 4675
rect 7573 4641 7607 4675
rect 2421 4573 2455 4607
rect 4721 4573 4755 4607
rect 3893 4505 3927 4539
rect 7757 4437 7791 4471
rect 7849 4641 7883 4675
rect 8620 4641 8654 4675
rect 9045 4641 9079 4675
rect 9689 4641 9723 4675
rect 9873 4641 9907 4675
rect 10517 4641 10551 4675
rect 11161 4641 11195 4675
rect 13185 4641 13219 4675
rect 13369 4641 13403 4675
rect 13829 4641 13863 4675
rect 14289 4641 14323 4675
rect 15117 4641 15151 4675
rect 16773 4641 16807 4675
rect 19073 4641 19107 4675
rect 10241 4573 10275 4607
rect 14381 4573 14415 4607
rect 15577 4573 15611 4607
rect 17417 4573 17451 4607
rect 17693 4573 17727 4607
rect 18889 4573 18923 4607
rect 12817 4505 12851 4539
rect 16497 4505 16531 4539
rect 18337 4505 18371 4539
rect 7849 4437 7883 4471
rect 8033 4437 8067 4471
rect 8723 4437 8757 4471
rect 2697 4233 2731 4267
rect 3065 4233 3099 4267
rect 5641 4233 5675 4267
rect 6561 4233 6595 4267
rect 12633 4233 12667 4267
rect 17233 4233 17267 4267
rect 17877 4233 17911 4267
rect 19073 4233 19107 4267
rect 5825 4165 5859 4199
rect 7665 4165 7699 4199
rect 11805 4165 11839 4199
rect 13093 4165 13127 4199
rect 13369 4165 13403 4199
rect 15301 4165 15335 4199
rect 1777 4097 1811 4131
rect 5549 4097 5583 4131
rect 5641 4097 5675 4131
rect 7205 4097 7239 4131
rect 12173 4097 12207 4131
rect 16037 4097 16071 4131
rect 16957 4097 16991 4131
rect 18153 4097 18187 4131
rect 18797 4097 18831 4131
rect 4721 4029 4755 4063
rect 5457 4029 5491 4063
rect 7849 4029 7883 4063
rect 8217 4029 8251 4063
rect 8585 4029 8619 4063
rect 9137 4029 9171 4063
rect 10057 4029 10091 4063
rect 10977 4029 11011 4063
rect 12449 4029 12483 4063
rect 13921 4029 13955 4063
rect 14381 4029 14415 4063
rect 14841 4029 14875 4063
rect 15117 4029 15151 4063
rect 19676 4029 19710 4063
rect 20085 4029 20119 4063
rect 1869 3961 1903 3995
rect 2421 3961 2455 3995
rect 3341 3961 3375 3995
rect 3433 3961 3467 3995
rect 3985 3961 4019 3995
rect 4353 3961 4387 3995
rect 10378 3961 10412 3995
rect 16313 3961 16347 3995
rect 16405 3961 16439 3995
rect 18245 3961 18279 3995
rect 19763 3961 19797 3995
rect 6193 3893 6227 3927
rect 7849 3893 7883 3927
rect 9505 3893 9539 3927
rect 9873 3893 9907 3927
rect 11253 3893 11287 3927
rect 13829 3893 13863 3927
rect 15669 3893 15703 3927
rect 19441 3893 19475 3927
rect 2881 3689 2915 3723
rect 3433 3689 3467 3723
rect 3893 3689 3927 3723
rect 4905 3689 4939 3723
rect 5089 3689 5123 3723
rect 7389 3689 7423 3723
rect 14289 3689 14323 3723
rect 14657 3689 14691 3723
rect 14933 3689 14967 3723
rect 16405 3689 16439 3723
rect 16681 3689 16715 3723
rect 19441 3689 19475 3723
rect 2323 3621 2357 3655
rect 9045 3621 9079 3655
rect 9505 3621 9539 3655
rect 13369 3621 13403 3655
rect 15485 3621 15519 3655
rect 17233 3621 17267 3655
rect 18797 3621 18831 3655
rect 5273 3553 5307 3587
rect 5457 3553 5491 3587
rect 6009 3553 6043 3587
rect 6377 3553 6411 3587
rect 6837 3553 6871 3587
rect 7297 3553 7331 3587
rect 7757 3553 7791 3587
rect 8125 3553 8159 3587
rect 8677 3553 8711 3587
rect 9781 3553 9815 3587
rect 11161 3553 11195 3587
rect 11345 3553 11379 3587
rect 11713 3553 11747 3587
rect 12265 3553 12299 3587
rect 12817 3553 12851 3587
rect 1961 3485 1995 3519
rect 7113 3485 7147 3519
rect 10793 3485 10827 3519
rect 12357 3485 12391 3519
rect 13277 3485 13311 3519
rect 13553 3485 13587 3519
rect 15393 3485 15427 3519
rect 15669 3485 15703 3519
rect 16957 3485 16991 3519
rect 17141 3485 17175 3519
rect 18705 3485 18739 3519
rect 9965 3417 9999 3451
rect 1777 3349 1811 3383
rect 4537 3349 4571 3383
rect 10609 3349 10643 3383
rect 10793 3349 10827 3383
rect 17693 3417 17727 3451
rect 18429 3417 18463 3451
rect 16957 3349 16991 3383
rect 18061 3349 18095 3383
rect 19625 3349 19659 3383
rect 2145 3145 2179 3179
rect 3617 3145 3651 3179
rect 4261 3145 4295 3179
rect 7113 3145 7147 3179
rect 7757 3145 7791 3179
rect 8125 3145 8159 3179
rect 10057 3145 10091 3179
rect 10517 3145 10551 3179
rect 11805 3145 11839 3179
rect 12173 3145 12207 3179
rect 15025 3145 15059 3179
rect 17141 3145 17175 3179
rect 17509 3145 17543 3179
rect 1823 3077 1857 3111
rect 6193 3077 6227 3111
rect 20085 3077 20119 3111
rect 10609 3009 10643 3043
rect 14197 3009 14231 3043
rect 1752 2941 1786 2975
rect 2697 2941 2731 2975
rect 3985 2941 4019 2975
rect 4721 2941 4755 2975
rect 4997 2941 5031 2975
rect 5457 2941 5491 2975
rect 5641 2941 5675 2975
rect 6653 2941 6687 2975
rect 7021 2941 7055 2975
rect 8309 2941 8343 2975
rect 8769 2941 8803 2975
rect 9321 2941 9355 2975
rect 9505 2941 9539 2975
rect 11529 2941 11563 2975
rect 13001 2941 13035 2975
rect 13185 2941 13219 2975
rect 13737 2941 13771 2975
rect 14105 2941 14139 2975
rect 14473 2941 14507 2975
rect 15577 2941 15611 2975
rect 19073 2941 19107 2975
rect 19676 2941 19710 2975
rect 20453 2941 20487 2975
rect 3018 2873 3052 2907
rect 6837 2873 6871 2907
rect 9781 2873 9815 2907
rect 10930 2873 10964 2907
rect 15393 2873 15427 2907
rect 15898 2873 15932 2907
rect 18153 2873 18187 2907
rect 18245 2873 18279 2907
rect 18797 2873 18831 2907
rect 19763 2873 19797 2907
rect 2513 2805 2547 2839
rect 4537 2805 4571 2839
rect 16497 2805 16531 2839
rect 17785 2805 17819 2839
rect 19441 2805 19475 2839
rect 1409 2601 1443 2635
rect 3525 2601 3559 2635
rect 3893 2601 3927 2635
rect 4629 2601 4663 2635
rect 6377 2601 6411 2635
rect 8309 2601 8343 2635
rect 11667 2601 11701 2635
rect 15623 2601 15657 2635
rect 19717 2601 19751 2635
rect 2513 2533 2547 2567
rect 2605 2533 2639 2567
rect 5410 2533 5444 2567
rect 6101 2533 6135 2567
rect 6653 2533 6687 2567
rect 9045 2533 9079 2567
rect 10102 2533 10136 2567
rect 12357 2533 12391 2567
rect 12909 2533 12943 2567
rect 13915 2533 13949 2567
rect 14841 2533 14875 2567
rect 16681 2533 16715 2567
rect 17233 2533 17267 2567
rect 18153 2533 18187 2567
rect 18521 2533 18555 2567
rect 19349 2533 19383 2567
rect 3157 2465 3191 2499
rect 4112 2465 4146 2499
rect 4905 2465 4939 2499
rect 5089 2465 5123 2499
rect 4813 2397 4847 2431
rect 4215 2329 4249 2363
rect 6929 2465 6963 2499
rect 7389 2465 7423 2499
rect 7757 2465 7791 2499
rect 8125 2465 8159 2499
rect 10701 2465 10735 2499
rect 11596 2465 11630 2499
rect 11897 2465 11931 2499
rect 13369 2465 13403 2499
rect 13553 2465 13587 2499
rect 14473 2465 14507 2499
rect 15552 2465 15586 2499
rect 16037 2465 16071 2499
rect 17509 2465 17543 2499
rect 8677 2397 8711 2431
rect 9781 2397 9815 2431
rect 11069 2397 11103 2431
rect 11437 2397 11471 2431
rect 16313 2397 16347 2431
rect 16589 2397 16623 2431
rect 18429 2397 18463 2431
rect 18705 2397 18739 2431
rect 20453 2397 20487 2431
rect 15117 2329 15151 2363
rect 20085 2329 20119 2363
rect 1961 2261 1995 2295
rect 4813 2261 4847 2295
rect 6009 2261 6043 2295
rect 6101 2261 6135 2295
rect 9505 2261 9539 2295
rect 11897 2261 11931 2295
rect 12081 2261 12115 2295
<< metal1 >>
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 17218 21536 17224 21548
rect 16632 21508 17224 21536
rect 16632 21496 16638 21508
rect 17218 21496 17224 21508
rect 17276 21496 17282 21548
rect 1104 19610 20884 19632
rect 1104 19558 4648 19610
rect 4700 19558 4712 19610
rect 4764 19558 4776 19610
rect 4828 19558 4840 19610
rect 4892 19558 11982 19610
rect 12034 19558 12046 19610
rect 12098 19558 12110 19610
rect 12162 19558 12174 19610
rect 12226 19558 19315 19610
rect 19367 19558 19379 19610
rect 19431 19558 19443 19610
rect 19495 19558 19507 19610
rect 19559 19558 20884 19610
rect 1104 19536 20884 19558
rect 1104 19066 20884 19088
rect 1104 19014 8315 19066
rect 8367 19014 8379 19066
rect 8431 19014 8443 19066
rect 8495 19014 8507 19066
rect 8559 19014 15648 19066
rect 15700 19014 15712 19066
rect 15764 19014 15776 19066
rect 15828 19014 15840 19066
rect 15892 19014 20884 19066
rect 1104 18992 20884 19014
rect 1104 18522 20884 18544
rect 1104 18470 4648 18522
rect 4700 18470 4712 18522
rect 4764 18470 4776 18522
rect 4828 18470 4840 18522
rect 4892 18470 11982 18522
rect 12034 18470 12046 18522
rect 12098 18470 12110 18522
rect 12162 18470 12174 18522
rect 12226 18470 19315 18522
rect 19367 18470 19379 18522
rect 19431 18470 19443 18522
rect 19495 18470 19507 18522
rect 19559 18470 20884 18522
rect 1104 18448 20884 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 4522 18368 4528 18420
rect 4580 18408 4586 18420
rect 4617 18411 4675 18417
rect 4617 18408 4629 18411
rect 4580 18380 4629 18408
rect 4580 18368 4586 18380
rect 4617 18377 4629 18380
rect 4663 18377 4675 18411
rect 7650 18408 7656 18420
rect 7611 18380 7656 18408
rect 4617 18371 4675 18377
rect 7650 18368 7656 18380
rect 7708 18368 7714 18420
rect 1302 18164 1308 18216
rect 1360 18204 1366 18216
rect 1397 18207 1455 18213
rect 1397 18204 1409 18207
rect 1360 18176 1409 18204
rect 1360 18164 1366 18176
rect 1397 18173 1409 18176
rect 1443 18204 1455 18207
rect 1949 18207 2007 18213
rect 1949 18204 1961 18207
rect 1443 18176 1961 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 1949 18173 1961 18176
rect 1995 18173 2007 18207
rect 1949 18167 2007 18173
rect 4433 18207 4491 18213
rect 4433 18173 4445 18207
rect 4479 18204 4491 18207
rect 7469 18207 7527 18213
rect 4479 18176 5120 18204
rect 4479 18173 4491 18176
rect 4433 18167 4491 18173
rect 5092 18077 5120 18176
rect 7469 18173 7481 18207
rect 7515 18204 7527 18207
rect 7515 18176 8156 18204
rect 7515 18173 7527 18176
rect 7469 18167 7527 18173
rect 5077 18071 5135 18077
rect 5077 18037 5089 18071
rect 5123 18068 5135 18071
rect 5258 18068 5264 18080
rect 5123 18040 5264 18068
rect 5123 18037 5135 18040
rect 5077 18031 5135 18037
rect 5258 18028 5264 18040
rect 5316 18028 5322 18080
rect 8128 18077 8156 18176
rect 8113 18071 8171 18077
rect 8113 18037 8125 18071
rect 8159 18068 8171 18071
rect 10226 18068 10232 18080
rect 8159 18040 10232 18068
rect 8159 18037 8171 18040
rect 8113 18031 8171 18037
rect 10226 18028 10232 18040
rect 10284 18028 10290 18080
rect 1104 17978 20884 18000
rect 1104 17926 8315 17978
rect 8367 17926 8379 17978
rect 8431 17926 8443 17978
rect 8495 17926 8507 17978
rect 8559 17926 15648 17978
rect 15700 17926 15712 17978
rect 15764 17926 15776 17978
rect 15828 17926 15840 17978
rect 15892 17926 20884 17978
rect 1104 17904 20884 17926
rect 1104 17434 20884 17456
rect 1104 17382 4648 17434
rect 4700 17382 4712 17434
rect 4764 17382 4776 17434
rect 4828 17382 4840 17434
rect 4892 17382 11982 17434
rect 12034 17382 12046 17434
rect 12098 17382 12110 17434
rect 12162 17382 12174 17434
rect 12226 17382 19315 17434
rect 19367 17382 19379 17434
rect 19431 17382 19443 17434
rect 19495 17382 19507 17434
rect 19559 17382 20884 17434
rect 1104 17360 20884 17382
rect 1104 16890 20884 16912
rect 1104 16838 8315 16890
rect 8367 16838 8379 16890
rect 8431 16838 8443 16890
rect 8495 16838 8507 16890
rect 8559 16838 15648 16890
rect 15700 16838 15712 16890
rect 15764 16838 15776 16890
rect 15828 16838 15840 16890
rect 15892 16838 20884 16890
rect 1104 16816 20884 16838
rect 1104 16346 20884 16368
rect 1104 16294 4648 16346
rect 4700 16294 4712 16346
rect 4764 16294 4776 16346
rect 4828 16294 4840 16346
rect 4892 16294 11982 16346
rect 12034 16294 12046 16346
rect 12098 16294 12110 16346
rect 12162 16294 12174 16346
rect 12226 16294 19315 16346
rect 19367 16294 19379 16346
rect 19431 16294 19443 16346
rect 19495 16294 19507 16346
rect 19559 16294 20884 16346
rect 1104 16272 20884 16294
rect 1104 15802 20884 15824
rect 1104 15750 8315 15802
rect 8367 15750 8379 15802
rect 8431 15750 8443 15802
rect 8495 15750 8507 15802
rect 8559 15750 15648 15802
rect 15700 15750 15712 15802
rect 15764 15750 15776 15802
rect 15828 15750 15840 15802
rect 15892 15750 20884 15802
rect 1104 15728 20884 15750
rect 1578 15688 1584 15700
rect 1539 15660 1584 15688
rect 1578 15648 1584 15660
rect 1636 15648 1642 15700
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 1104 15258 20884 15280
rect 1104 15206 4648 15258
rect 4700 15206 4712 15258
rect 4764 15206 4776 15258
rect 4828 15206 4840 15258
rect 4892 15206 11982 15258
rect 12034 15206 12046 15258
rect 12098 15206 12110 15258
rect 12162 15206 12174 15258
rect 12226 15206 19315 15258
rect 19367 15206 19379 15258
rect 19431 15206 19443 15258
rect 19495 15206 19507 15258
rect 19559 15206 20884 15258
rect 1104 15184 20884 15206
rect 1394 14764 1400 14816
rect 1452 14804 1458 14816
rect 1673 14807 1731 14813
rect 1673 14804 1685 14807
rect 1452 14776 1685 14804
rect 1452 14764 1458 14776
rect 1673 14773 1685 14776
rect 1719 14804 1731 14807
rect 5350 14804 5356 14816
rect 1719 14776 5356 14804
rect 1719 14773 1731 14776
rect 1673 14767 1731 14773
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 1104 14714 20884 14736
rect 1104 14662 8315 14714
rect 8367 14662 8379 14714
rect 8431 14662 8443 14714
rect 8495 14662 8507 14714
rect 8559 14662 15648 14714
rect 15700 14662 15712 14714
rect 15764 14662 15776 14714
rect 15828 14662 15840 14714
rect 15892 14662 20884 14714
rect 1104 14640 20884 14662
rect 1104 14170 20884 14192
rect 1104 14118 4648 14170
rect 4700 14118 4712 14170
rect 4764 14118 4776 14170
rect 4828 14118 4840 14170
rect 4892 14118 11982 14170
rect 12034 14118 12046 14170
rect 12098 14118 12110 14170
rect 12162 14118 12174 14170
rect 12226 14118 19315 14170
rect 19367 14118 19379 14170
rect 19431 14118 19443 14170
rect 19495 14118 19507 14170
rect 19559 14118 20884 14170
rect 1104 14096 20884 14118
rect 1104 13626 20884 13648
rect 1104 13574 8315 13626
rect 8367 13574 8379 13626
rect 8431 13574 8443 13626
rect 8495 13574 8507 13626
rect 8559 13574 15648 13626
rect 15700 13574 15712 13626
rect 15764 13574 15776 13626
rect 15828 13574 15840 13626
rect 15892 13574 20884 13626
rect 1104 13552 20884 13574
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 13814 13376 13820 13388
rect 13044 13348 13820 13376
rect 13044 13336 13050 13348
rect 13814 13336 13820 13348
rect 13872 13336 13878 13388
rect 19058 13376 19064 13388
rect 19019 13348 19064 13376
rect 19058 13336 19064 13348
rect 19116 13336 19122 13388
rect 19242 13240 19248 13252
rect 19203 13212 19248 13240
rect 19242 13200 19248 13212
rect 19300 13200 19306 13252
rect 1104 13082 20884 13104
rect 1104 13030 4648 13082
rect 4700 13030 4712 13082
rect 4764 13030 4776 13082
rect 4828 13030 4840 13082
rect 4892 13030 11982 13082
rect 12034 13030 12046 13082
rect 12098 13030 12110 13082
rect 12162 13030 12174 13082
rect 12226 13030 19315 13082
rect 19367 13030 19379 13082
rect 19431 13030 19443 13082
rect 19495 13030 19507 13082
rect 19559 13030 20884 13082
rect 1104 13008 20884 13030
rect 18506 12588 18512 12640
rect 18564 12628 18570 12640
rect 19058 12628 19064 12640
rect 18564 12600 19064 12628
rect 18564 12588 18570 12600
rect 19058 12588 19064 12600
rect 19116 12588 19122 12640
rect 1104 12538 20884 12560
rect 1104 12486 8315 12538
rect 8367 12486 8379 12538
rect 8431 12486 8443 12538
rect 8495 12486 8507 12538
rect 8559 12486 15648 12538
rect 15700 12486 15712 12538
rect 15764 12486 15776 12538
rect 15828 12486 15840 12538
rect 15892 12486 20884 12538
rect 1104 12464 20884 12486
rect 1104 11994 20884 12016
rect 1104 11942 4648 11994
rect 4700 11942 4712 11994
rect 4764 11942 4776 11994
rect 4828 11942 4840 11994
rect 4892 11942 11982 11994
rect 12034 11942 12046 11994
rect 12098 11942 12110 11994
rect 12162 11942 12174 11994
rect 12226 11942 19315 11994
rect 19367 11942 19379 11994
rect 19431 11942 19443 11994
rect 19495 11942 19507 11994
rect 19559 11942 20884 11994
rect 1104 11920 20884 11942
rect 1104 11450 20884 11472
rect 1104 11398 8315 11450
rect 8367 11398 8379 11450
rect 8431 11398 8443 11450
rect 8495 11398 8507 11450
rect 8559 11398 15648 11450
rect 15700 11398 15712 11450
rect 15764 11398 15776 11450
rect 15828 11398 15840 11450
rect 15892 11398 20884 11450
rect 1104 11376 20884 11398
rect 19245 11339 19303 11345
rect 19245 11305 19257 11339
rect 19291 11336 19303 11339
rect 19334 11336 19340 11348
rect 19291 11308 19340 11336
rect 19291 11305 19303 11308
rect 19245 11299 19303 11305
rect 19334 11296 19340 11308
rect 19392 11296 19398 11348
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11200 9735 11203
rect 9766 11200 9772 11212
rect 9723 11172 9772 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 19058 11200 19064 11212
rect 19019 11172 19064 11200
rect 19058 11160 19064 11172
rect 19116 11160 19122 11212
rect 8110 11092 8116 11144
rect 8168 11132 8174 11144
rect 8205 11135 8263 11141
rect 8205 11132 8217 11135
rect 8168 11104 8217 11132
rect 8168 11092 8174 11104
rect 8205 11101 8217 11104
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 6914 10996 6920 11008
rect 6875 10968 6920 10996
rect 6914 10956 6920 10968
rect 6972 10956 6978 11008
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 9815 10999 9873 11005
rect 9815 10996 9827 10999
rect 9732 10968 9827 10996
rect 9732 10956 9738 10968
rect 9815 10965 9827 10968
rect 9861 10965 9873 10999
rect 9815 10959 9873 10965
rect 1104 10906 20884 10928
rect 1104 10854 4648 10906
rect 4700 10854 4712 10906
rect 4764 10854 4776 10906
rect 4828 10854 4840 10906
rect 4892 10854 11982 10906
rect 12034 10854 12046 10906
rect 12098 10854 12110 10906
rect 12162 10854 12174 10906
rect 12226 10854 19315 10906
rect 19367 10854 19379 10906
rect 19431 10854 19443 10906
rect 19495 10854 19507 10906
rect 19559 10854 20884 10906
rect 1104 10832 20884 10854
rect 10091 10795 10149 10801
rect 10091 10761 10103 10795
rect 10137 10792 10149 10795
rect 10318 10792 10324 10804
rect 10137 10764 10324 10792
rect 10137 10761 10149 10764
rect 10091 10755 10149 10761
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 8389 10591 8447 10597
rect 8389 10588 8401 10591
rect 8260 10560 8401 10588
rect 8260 10548 8266 10560
rect 8389 10557 8401 10560
rect 8435 10557 8447 10591
rect 8389 10551 8447 10557
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 6914 10520 6920 10532
rect 6875 10492 6920 10520
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 7009 10523 7067 10529
rect 7009 10489 7021 10523
rect 7055 10489 7067 10523
rect 7558 10520 7564 10532
rect 7519 10492 7564 10520
rect 7009 10483 7067 10489
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 6052 10424 6561 10452
rect 6052 10412 6058 10424
rect 6549 10421 6561 10424
rect 6595 10452 6607 10455
rect 7024 10452 7052 10483
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 7742 10480 7748 10532
rect 7800 10520 7806 10532
rect 8297 10523 8355 10529
rect 8297 10520 8309 10523
rect 7800 10492 8309 10520
rect 7800 10480 7806 10492
rect 8297 10489 8309 10492
rect 8343 10520 8355 10523
rect 8588 10520 8616 10551
rect 9582 10548 9588 10600
rect 9640 10588 9646 10600
rect 9988 10591 10046 10597
rect 9988 10588 10000 10591
rect 9640 10560 10000 10588
rect 9640 10548 9646 10560
rect 9988 10557 10000 10560
rect 10034 10588 10046 10591
rect 10413 10591 10471 10597
rect 10413 10588 10425 10591
rect 10034 10560 10425 10588
rect 10034 10557 10046 10560
rect 9988 10551 10046 10557
rect 10413 10557 10425 10560
rect 10459 10557 10471 10591
rect 10413 10551 10471 10557
rect 10870 10548 10876 10600
rect 10928 10588 10934 10600
rect 11000 10591 11058 10597
rect 11000 10588 11012 10591
rect 10928 10560 11012 10588
rect 10928 10548 10934 10560
rect 11000 10557 11012 10560
rect 11046 10588 11058 10591
rect 11425 10591 11483 10597
rect 11425 10588 11437 10591
rect 11046 10560 11437 10588
rect 11046 10557 11058 10560
rect 11000 10551 11058 10557
rect 11425 10557 11437 10560
rect 11471 10557 11483 10591
rect 11425 10551 11483 10557
rect 12504 10591 12562 10597
rect 12504 10557 12516 10591
rect 12550 10588 12562 10591
rect 12550 10560 12940 10588
rect 12550 10557 12562 10560
rect 12504 10551 12562 10557
rect 8343 10492 8616 10520
rect 8343 10489 8355 10492
rect 8297 10483 8355 10489
rect 12912 10464 12940 10560
rect 9766 10452 9772 10464
rect 6595 10424 7052 10452
rect 9679 10424 9772 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 9766 10412 9772 10424
rect 9824 10452 9830 10464
rect 10778 10452 10784 10464
rect 9824 10424 10784 10452
rect 9824 10412 9830 10424
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 11103 10455 11161 10461
rect 11103 10421 11115 10455
rect 11149 10452 11161 10455
rect 11330 10452 11336 10464
rect 11149 10424 11336 10452
rect 11149 10421 11161 10424
rect 11103 10415 11161 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12575 10455 12633 10461
rect 12575 10421 12587 10455
rect 12621 10452 12633 10455
rect 12710 10452 12716 10464
rect 12621 10424 12716 10452
rect 12621 10421 12633 10424
rect 12575 10415 12633 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 12894 10452 12900 10464
rect 12855 10424 12900 10452
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 15378 10412 15384 10464
rect 15436 10452 15442 10464
rect 19058 10452 19064 10464
rect 15436 10424 19064 10452
rect 15436 10412 15442 10424
rect 19058 10412 19064 10424
rect 19116 10412 19122 10464
rect 1104 10362 20884 10384
rect 1104 10310 8315 10362
rect 8367 10310 8379 10362
rect 8431 10310 8443 10362
rect 8495 10310 8507 10362
rect 8559 10310 15648 10362
rect 15700 10310 15712 10362
rect 15764 10310 15776 10362
rect 15828 10310 15840 10362
rect 15892 10310 20884 10362
rect 1104 10288 20884 10310
rect 7558 10248 7564 10260
rect 7208 10220 7564 10248
rect 6546 10140 6552 10192
rect 6604 10180 6610 10192
rect 7208 10189 7236 10220
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 6641 10183 6699 10189
rect 6641 10180 6653 10183
rect 6604 10152 6653 10180
rect 6604 10140 6610 10152
rect 6641 10149 6653 10152
rect 6687 10149 6699 10183
rect 6641 10143 6699 10149
rect 7193 10183 7251 10189
rect 7193 10149 7205 10183
rect 7239 10149 7251 10183
rect 8110 10180 8116 10192
rect 8071 10152 8116 10180
rect 7193 10143 7251 10149
rect 8110 10140 8116 10152
rect 8168 10140 8174 10192
rect 8202 10140 8208 10192
rect 8260 10180 8266 10192
rect 9766 10180 9772 10192
rect 8260 10152 8305 10180
rect 9727 10152 9772 10180
rect 8260 10140 8266 10152
rect 9766 10140 9772 10152
rect 9824 10140 9830 10192
rect 9861 10183 9919 10189
rect 9861 10149 9873 10183
rect 9907 10180 9919 10183
rect 10134 10180 10140 10192
rect 9907 10152 10140 10180
rect 9907 10149 9919 10152
rect 9861 10143 9919 10149
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 12342 10112 12348 10124
rect 12303 10084 12348 10112
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 6362 10004 6368 10056
rect 6420 10044 6426 10056
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 6420 10016 6561 10044
rect 6420 10004 6426 10016
rect 6549 10013 6561 10016
rect 6595 10013 6607 10047
rect 8386 10044 8392 10056
rect 8347 10016 8392 10044
rect 6549 10007 6607 10013
rect 8386 10004 8392 10016
rect 8444 10044 8450 10056
rect 9582 10044 9588 10056
rect 8444 10016 9588 10044
rect 8444 10004 8450 10016
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 9766 10044 9772 10056
rect 9692 10016 9772 10044
rect 6270 9936 6276 9988
rect 6328 9976 6334 9988
rect 9692 9976 9720 10016
rect 9766 10004 9772 10016
rect 9824 10004 9830 10056
rect 10413 10047 10471 10053
rect 10413 10013 10425 10047
rect 10459 10044 10471 10047
rect 13538 10044 13544 10056
rect 10459 10016 13544 10044
rect 10459 10013 10471 10016
rect 10413 10007 10471 10013
rect 6328 9948 9720 9976
rect 6328 9936 6334 9948
rect 9214 9908 9220 9920
rect 9127 9880 9220 9908
rect 9214 9868 9220 9880
rect 9272 9908 9278 9920
rect 10428 9908 10456 10007
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 10778 9936 10784 9988
rect 10836 9976 10842 9988
rect 13722 9976 13728 9988
rect 10836 9948 13728 9976
rect 10836 9936 10842 9948
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 12434 9908 12440 9920
rect 9272 9880 10456 9908
rect 12395 9880 12440 9908
rect 9272 9868 9278 9880
rect 12434 9868 12440 9880
rect 12492 9868 12498 9920
rect 1104 9818 20884 9840
rect 1104 9766 4648 9818
rect 4700 9766 4712 9818
rect 4764 9766 4776 9818
rect 4828 9766 4840 9818
rect 4892 9766 11982 9818
rect 12034 9766 12046 9818
rect 12098 9766 12110 9818
rect 12162 9766 12174 9818
rect 12226 9766 19315 9818
rect 19367 9766 19379 9818
rect 19431 9766 19443 9818
rect 19495 9766 19507 9818
rect 19559 9766 20884 9818
rect 1104 9744 20884 9766
rect 4847 9707 4905 9713
rect 4847 9673 4859 9707
rect 4893 9704 4905 9707
rect 6362 9704 6368 9716
rect 4893 9676 6368 9704
rect 4893 9673 4905 9676
rect 4847 9667 4905 9673
rect 6362 9664 6368 9676
rect 6420 9704 6426 9716
rect 7009 9707 7067 9713
rect 7009 9704 7021 9707
rect 6420 9676 7021 9704
rect 6420 9664 6426 9676
rect 7009 9673 7021 9676
rect 7055 9673 7067 9707
rect 7009 9667 7067 9673
rect 8202 9664 8208 9716
rect 8260 9704 8266 9716
rect 8573 9707 8631 9713
rect 8573 9704 8585 9707
rect 8260 9676 8585 9704
rect 8260 9664 8266 9676
rect 8573 9673 8585 9676
rect 8619 9673 8631 9707
rect 8573 9667 8631 9673
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 10505 9707 10563 9713
rect 10505 9704 10517 9707
rect 9824 9676 10517 9704
rect 9824 9664 9830 9676
rect 10505 9673 10517 9676
rect 10551 9673 10563 9707
rect 10505 9667 10563 9673
rect 12253 9707 12311 9713
rect 12253 9673 12265 9707
rect 12299 9704 12311 9707
rect 12342 9704 12348 9716
rect 12299 9676 12348 9704
rect 12299 9673 12311 9676
rect 12253 9667 12311 9673
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 16761 9707 16819 9713
rect 16761 9704 16773 9707
rect 16632 9676 16773 9704
rect 16632 9664 16638 9676
rect 16761 9673 16773 9676
rect 16807 9673 16819 9707
rect 16761 9667 16819 9673
rect 5258 9636 5264 9648
rect 5219 9608 5264 9636
rect 5258 9596 5264 9608
rect 5316 9596 5322 9648
rect 5859 9639 5917 9645
rect 5859 9605 5871 9639
rect 5905 9636 5917 9639
rect 6914 9636 6920 9648
rect 5905 9608 6920 9636
rect 5905 9605 5917 9608
rect 5859 9599 5917 9605
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 7558 9596 7564 9648
rect 7616 9636 7622 9648
rect 11149 9639 11207 9645
rect 7616 9608 7696 9636
rect 7616 9596 7622 9608
rect 4776 9503 4834 9509
rect 4776 9469 4788 9503
rect 4822 9500 4834 9503
rect 5276 9500 5304 9596
rect 7668 9577 7696 9608
rect 11149 9605 11161 9639
rect 11195 9636 11207 9639
rect 21542 9636 21548 9648
rect 11195 9608 21548 9636
rect 11195 9605 11207 9608
rect 11149 9599 11207 9605
rect 21542 9596 21548 9608
rect 21600 9596 21606 9648
rect 7653 9571 7711 9577
rect 7653 9537 7665 9571
rect 7699 9537 7711 9571
rect 7653 9531 7711 9537
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8386 9568 8392 9580
rect 8343 9540 8392 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 9214 9568 9220 9580
rect 9175 9540 9220 9568
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9568 12587 9571
rect 12710 9568 12716 9580
rect 12575 9540 12716 9568
rect 12575 9537 12587 9540
rect 12529 9531 12587 9537
rect 12710 9528 12716 9540
rect 12768 9568 12774 9580
rect 13449 9571 13507 9577
rect 13449 9568 13461 9571
rect 12768 9540 13461 9568
rect 12768 9528 12774 9540
rect 13449 9537 13461 9540
rect 13495 9537 13507 9571
rect 13449 9531 13507 9537
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 17770 9568 17776 9580
rect 13780 9540 17776 9568
rect 13780 9528 13786 9540
rect 17770 9528 17776 9540
rect 17828 9568 17834 9580
rect 19702 9568 19708 9580
rect 17828 9540 19708 9568
rect 17828 9528 17834 9540
rect 19702 9528 19708 9540
rect 19760 9528 19766 9580
rect 4822 9472 5304 9500
rect 4822 9469 4834 9472
rect 4776 9463 4834 9469
rect 5350 9460 5356 9512
rect 5408 9500 5414 9512
rect 5788 9503 5846 9509
rect 5788 9500 5800 9503
rect 5408 9472 5800 9500
rect 5408 9460 5414 9472
rect 5788 9469 5800 9472
rect 5834 9500 5846 9503
rect 10962 9500 10968 9512
rect 5834 9472 6316 9500
rect 10923 9472 10968 9500
rect 5834 9469 5846 9472
rect 5788 9463 5846 9469
rect 6288 9373 6316 9472
rect 10962 9460 10968 9472
rect 11020 9500 11026 9512
rect 11517 9503 11575 9509
rect 11517 9500 11529 9503
rect 11020 9472 11529 9500
rect 11020 9460 11026 9472
rect 11517 9469 11529 9472
rect 11563 9500 11575 9503
rect 11790 9500 11796 9512
rect 11563 9472 11796 9500
rect 11563 9469 11575 9472
rect 11517 9463 11575 9469
rect 11790 9460 11796 9472
rect 11848 9460 11854 9512
rect 15600 9503 15658 9509
rect 15600 9500 15612 9503
rect 13786 9472 15612 9500
rect 7469 9435 7527 9441
rect 7469 9401 7481 9435
rect 7515 9432 7527 9435
rect 7742 9432 7748 9444
rect 7515 9404 7748 9432
rect 7515 9401 7527 9404
rect 7469 9395 7527 9401
rect 7742 9392 7748 9404
rect 7800 9392 7806 9444
rect 9306 9392 9312 9444
rect 9364 9432 9370 9444
rect 9858 9432 9864 9444
rect 9364 9404 9409 9432
rect 9771 9404 9864 9432
rect 9364 9392 9370 9404
rect 9858 9392 9864 9404
rect 9916 9432 9922 9444
rect 11422 9432 11428 9444
rect 9916 9404 11428 9432
rect 9916 9392 9922 9404
rect 11422 9392 11428 9404
rect 11480 9392 11486 9444
rect 12618 9432 12624 9444
rect 12579 9404 12624 9432
rect 12618 9392 12624 9404
rect 12676 9392 12682 9444
rect 13170 9432 13176 9444
rect 13131 9404 13176 9432
rect 13170 9392 13176 9404
rect 13228 9392 13234 9444
rect 6273 9367 6331 9373
rect 6273 9333 6285 9367
rect 6319 9364 6331 9367
rect 6362 9364 6368 9376
rect 6319 9336 6368 9364
rect 6319 9333 6331 9336
rect 6273 9327 6331 9333
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 6546 9364 6552 9376
rect 6507 9336 6552 9364
rect 6546 9324 6552 9336
rect 6604 9324 6610 9376
rect 9033 9367 9091 9373
rect 9033 9333 9045 9367
rect 9079 9364 9091 9367
rect 9324 9364 9352 9392
rect 10134 9364 10140 9376
rect 9079 9336 9352 9364
rect 10095 9336 10140 9364
rect 9079 9333 9091 9336
rect 9033 9327 9091 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 11146 9324 11152 9376
rect 11204 9364 11210 9376
rect 12894 9364 12900 9376
rect 11204 9336 12900 9364
rect 11204 9324 11210 9336
rect 12894 9324 12900 9336
rect 12952 9364 12958 9376
rect 13786 9364 13814 9472
rect 15600 9469 15612 9472
rect 15646 9500 15658 9503
rect 16025 9503 16083 9509
rect 16025 9500 16037 9503
rect 15646 9472 16037 9500
rect 15646 9469 15658 9472
rect 15600 9463 15658 9469
rect 16025 9469 16037 9472
rect 16071 9469 16083 9503
rect 16025 9463 16083 9469
rect 16577 9503 16635 9509
rect 16577 9469 16589 9503
rect 16623 9500 16635 9503
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 16623 9472 17233 9500
rect 16623 9469 16635 9472
rect 16577 9463 16635 9469
rect 17221 9469 17233 9472
rect 17267 9500 17279 9503
rect 17862 9500 17868 9512
rect 17267 9472 17868 9500
rect 17267 9469 17279 9472
rect 17221 9463 17279 9469
rect 16040 9432 16068 9463
rect 17862 9460 17868 9472
rect 17920 9460 17926 9512
rect 18116 9503 18174 9509
rect 18116 9469 18128 9503
rect 18162 9500 18174 9503
rect 18506 9500 18512 9512
rect 18162 9472 18512 9500
rect 18162 9469 18174 9472
rect 18116 9463 18174 9469
rect 18506 9460 18512 9472
rect 18564 9460 18570 9512
rect 19128 9503 19186 9509
rect 19128 9469 19140 9503
rect 19174 9500 19186 9503
rect 19242 9500 19248 9512
rect 19174 9472 19248 9500
rect 19174 9469 19186 9472
rect 19128 9463 19186 9469
rect 19242 9460 19248 9472
rect 19300 9500 19306 9512
rect 19521 9503 19579 9509
rect 19521 9500 19533 9503
rect 19300 9472 19533 9500
rect 19300 9460 19306 9472
rect 19521 9469 19533 9472
rect 19567 9469 19579 9503
rect 19521 9463 19579 9469
rect 17770 9432 17776 9444
rect 16040 9404 17776 9432
rect 17770 9392 17776 9404
rect 17828 9392 17834 9444
rect 12952 9336 13814 9364
rect 14185 9367 14243 9373
rect 12952 9324 12958 9336
rect 14185 9333 14197 9367
rect 14231 9364 14243 9367
rect 15194 9364 15200 9376
rect 14231 9336 15200 9364
rect 14231 9333 14243 9336
rect 14185 9327 14243 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 15703 9367 15761 9373
rect 15703 9333 15715 9367
rect 15749 9364 15761 9367
rect 15930 9364 15936 9376
rect 15749 9336 15936 9364
rect 15749 9333 15761 9336
rect 15703 9327 15761 9333
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 17218 9324 17224 9376
rect 17276 9364 17282 9376
rect 18187 9367 18245 9373
rect 18187 9364 18199 9367
rect 17276 9336 18199 9364
rect 17276 9324 17282 9336
rect 18187 9333 18199 9336
rect 18233 9333 18245 9367
rect 18187 9327 18245 9333
rect 18322 9324 18328 9376
rect 18380 9364 18386 9376
rect 19199 9367 19257 9373
rect 19199 9364 19211 9367
rect 18380 9336 19211 9364
rect 18380 9324 18386 9336
rect 19199 9333 19211 9336
rect 19245 9333 19257 9367
rect 19199 9327 19257 9333
rect 1104 9274 20884 9296
rect 1104 9222 8315 9274
rect 8367 9222 8379 9274
rect 8431 9222 8443 9274
rect 8495 9222 8507 9274
rect 8559 9222 15648 9274
rect 15700 9222 15712 9274
rect 15764 9222 15776 9274
rect 15828 9222 15840 9274
rect 15892 9222 20884 9274
rect 1104 9200 20884 9222
rect 7282 9160 7288 9172
rect 7243 9132 7288 9160
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 7837 9163 7895 9169
rect 7837 9160 7849 9163
rect 7800 9132 7849 9160
rect 7800 9120 7806 9132
rect 7837 9129 7849 9132
rect 7883 9129 7895 9163
rect 8110 9160 8116 9172
rect 8071 9132 8116 9160
rect 7837 9123 7895 9129
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 10873 9163 10931 9169
rect 10873 9160 10885 9163
rect 9732 9132 10885 9160
rect 9732 9120 9738 9132
rect 10873 9129 10885 9132
rect 10919 9129 10931 9163
rect 14090 9160 14096 9172
rect 14003 9132 14096 9160
rect 10873 9123 10931 9129
rect 14090 9120 14096 9132
rect 14148 9160 14154 9172
rect 18322 9160 18328 9172
rect 14148 9132 18328 9160
rect 14148 9120 14154 9132
rect 18322 9120 18328 9132
rect 18380 9120 18386 9172
rect 19150 9120 19156 9172
rect 19208 9160 19214 9172
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 19208 9132 19257 9160
rect 19208 9120 19214 9132
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 19245 9123 19303 9129
rect 6089 9095 6147 9101
rect 6089 9061 6101 9095
rect 6135 9092 6147 9095
rect 6546 9092 6552 9104
rect 6135 9064 6552 9092
rect 6135 9061 6147 9064
rect 6089 9055 6147 9061
rect 6546 9052 6552 9064
rect 6604 9052 6610 9104
rect 10042 9052 10048 9104
rect 10100 9092 10106 9104
rect 11470 9095 11528 9101
rect 11470 9092 11482 9095
rect 10100 9064 11482 9092
rect 10100 9052 10106 9064
rect 11470 9061 11482 9064
rect 11516 9061 11528 9095
rect 12529 9095 12587 9101
rect 12529 9092 12541 9095
rect 11470 9055 11528 9061
rect 12084 9064 12541 9092
rect 1302 8984 1308 9036
rect 1360 9024 1366 9036
rect 1524 9027 1582 9033
rect 1524 9024 1536 9027
rect 1360 8996 1536 9024
rect 1360 8984 1366 8996
rect 1524 8993 1536 8996
rect 1570 8993 1582 9027
rect 5994 9024 6000 9036
rect 5955 8996 6000 9024
rect 1524 8987 1582 8993
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 12084 9033 12112 9064
rect 12529 9061 12541 9064
rect 12575 9092 12587 9095
rect 12618 9092 12624 9104
rect 12575 9064 12624 9092
rect 12575 9061 12587 9064
rect 12529 9055 12587 9061
rect 12618 9052 12624 9064
rect 12676 9092 12682 9104
rect 13081 9095 13139 9101
rect 13081 9092 13093 9095
rect 12676 9064 13093 9092
rect 12676 9052 12682 9064
rect 13081 9061 13093 9064
rect 13127 9092 13139 9095
rect 13446 9092 13452 9104
rect 13127 9064 13452 9092
rect 13127 9061 13139 9064
rect 13081 9055 13139 9061
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 15930 9052 15936 9104
rect 15988 9092 15994 9104
rect 16298 9092 16304 9104
rect 15988 9064 16304 9092
rect 15988 9052 15994 9064
rect 16298 9052 16304 9064
rect 16356 9092 16362 9104
rect 16485 9095 16543 9101
rect 16485 9092 16497 9095
rect 16356 9064 16497 9092
rect 16356 9052 16362 9064
rect 16485 9061 16497 9064
rect 16531 9061 16543 9095
rect 16485 9055 16543 9061
rect 16574 9052 16580 9104
rect 16632 9092 16638 9104
rect 16632 9064 16677 9092
rect 16632 9052 16638 9064
rect 9712 9027 9770 9033
rect 9712 9024 9724 9027
rect 9548 8996 9724 9024
rect 9548 8984 9554 8996
rect 9712 8993 9724 8996
rect 9758 9024 9770 9027
rect 12069 9027 12127 9033
rect 9758 8996 11284 9024
rect 9758 8993 9770 8996
rect 9712 8987 9770 8993
rect 6917 8959 6975 8965
rect 6917 8956 6929 8959
rect 6472 8928 6929 8956
rect 1627 8891 1685 8897
rect 1627 8857 1639 8891
rect 1673 8888 1685 8891
rect 6270 8888 6276 8900
rect 1673 8860 6276 8888
rect 1673 8857 1685 8860
rect 1627 8851 1685 8857
rect 6270 8848 6276 8860
rect 6328 8848 6334 8900
rect 6472 8832 6500 8928
rect 6917 8925 6929 8928
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 11149 8959 11207 8965
rect 11149 8956 11161 8959
rect 11112 8928 11161 8956
rect 11112 8916 11118 8928
rect 11149 8925 11161 8928
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 8110 8848 8116 8900
rect 8168 8888 8174 8900
rect 8849 8891 8907 8897
rect 8849 8888 8861 8891
rect 8168 8860 8861 8888
rect 8168 8848 8174 8860
rect 8849 8857 8861 8860
rect 8895 8857 8907 8891
rect 8849 8851 8907 8857
rect 9815 8891 9873 8897
rect 9815 8857 9827 8891
rect 9861 8888 9873 8891
rect 10594 8888 10600 8900
rect 9861 8860 10600 8888
rect 9861 8857 9873 8860
rect 9815 8851 9873 8857
rect 10594 8848 10600 8860
rect 10652 8848 10658 8900
rect 6454 8820 6460 8832
rect 6415 8792 6460 8820
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 6822 8820 6828 8832
rect 6783 8792 6828 8820
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 7926 8780 7932 8832
rect 7984 8820 7990 8832
rect 8481 8823 8539 8829
rect 8481 8820 8493 8823
rect 7984 8792 8493 8820
rect 7984 8780 7990 8792
rect 8481 8789 8493 8792
rect 8527 8789 8539 8823
rect 9214 8820 9220 8832
rect 9175 8792 9220 8820
rect 8481 8783 8539 8789
rect 9214 8780 9220 8792
rect 9272 8780 9278 8832
rect 9950 8780 9956 8832
rect 10008 8820 10014 8832
rect 10137 8823 10195 8829
rect 10137 8820 10149 8823
rect 10008 8792 10149 8820
rect 10008 8780 10014 8792
rect 10137 8789 10149 8792
rect 10183 8789 10195 8823
rect 10502 8820 10508 8832
rect 10463 8792 10508 8820
rect 10137 8783 10195 8789
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 11256 8820 11284 8996
rect 12069 8993 12081 9027
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 15102 8984 15108 9036
rect 15160 9024 15166 9036
rect 15416 9027 15474 9033
rect 15416 9024 15428 9027
rect 15160 8996 15428 9024
rect 15160 8984 15166 8996
rect 15416 8993 15428 8996
rect 15462 8993 15474 9027
rect 15416 8987 15474 8993
rect 17862 8984 17868 9036
rect 17920 9024 17926 9036
rect 17992 9027 18050 9033
rect 17992 9024 18004 9027
rect 17920 8996 18004 9024
rect 17920 8984 17926 8996
rect 17992 8993 18004 8996
rect 18038 8993 18050 9027
rect 17992 8987 18050 8993
rect 19061 9027 19119 9033
rect 19061 8993 19073 9027
rect 19107 9024 19119 9027
rect 19150 9024 19156 9036
rect 19107 8996 19156 9024
rect 19107 8993 19119 8996
rect 19061 8987 19119 8993
rect 19150 8984 19156 8996
rect 19208 8984 19214 9036
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 11388 8928 13001 8956
rect 11388 8916 11394 8928
rect 12989 8925 13001 8928
rect 13035 8956 13047 8959
rect 14369 8959 14427 8965
rect 14369 8956 14381 8959
rect 13035 8928 14381 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 14369 8925 14381 8928
rect 14415 8925 14427 8959
rect 14369 8919 14427 8925
rect 17129 8959 17187 8965
rect 17129 8925 17141 8959
rect 17175 8956 17187 8959
rect 18414 8956 18420 8968
rect 17175 8928 18420 8956
rect 17175 8925 17187 8928
rect 17129 8919 17187 8925
rect 18414 8916 18420 8928
rect 18472 8916 18478 8968
rect 13538 8888 13544 8900
rect 13499 8860 13544 8888
rect 13538 8848 13544 8860
rect 13596 8848 13602 8900
rect 15378 8820 15384 8832
rect 11256 8792 15384 8820
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15519 8823 15577 8829
rect 15519 8789 15531 8823
rect 15565 8820 15577 8823
rect 16206 8820 16212 8832
rect 15565 8792 16212 8820
rect 15565 8789 15577 8792
rect 15519 8783 15577 8789
rect 16206 8780 16212 8792
rect 16264 8780 16270 8832
rect 16301 8823 16359 8829
rect 16301 8789 16313 8823
rect 16347 8820 16359 8823
rect 16482 8820 16488 8832
rect 16347 8792 16488 8820
rect 16347 8789 16359 8792
rect 16301 8783 16359 8789
rect 16482 8780 16488 8792
rect 16540 8820 16546 8832
rect 18095 8823 18153 8829
rect 18095 8820 18107 8823
rect 16540 8792 18107 8820
rect 16540 8780 16546 8792
rect 18095 8789 18107 8792
rect 18141 8789 18153 8823
rect 18095 8783 18153 8789
rect 1104 8730 20884 8752
rect 1104 8678 4648 8730
rect 4700 8678 4712 8730
rect 4764 8678 4776 8730
rect 4828 8678 4840 8730
rect 4892 8678 11982 8730
rect 12034 8678 12046 8730
rect 12098 8678 12110 8730
rect 12162 8678 12174 8730
rect 12226 8678 19315 8730
rect 19367 8678 19379 8730
rect 19431 8678 19443 8730
rect 19495 8678 19507 8730
rect 19559 8678 20884 8730
rect 1104 8656 20884 8678
rect 1302 8576 1308 8628
rect 1360 8616 1366 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1360 8588 1593 8616
rect 1360 8576 1366 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 1581 8579 1639 8585
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 6052 8588 6193 8616
rect 6052 8576 6058 8588
rect 6181 8585 6193 8588
rect 6227 8616 6239 8619
rect 7745 8619 7803 8625
rect 7745 8616 7757 8619
rect 6227 8588 7757 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 7745 8585 7757 8588
rect 7791 8585 7803 8619
rect 13446 8616 13452 8628
rect 13407 8588 13452 8616
rect 7745 8579 7803 8585
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 15102 8576 15108 8628
rect 15160 8616 15166 8628
rect 15381 8619 15439 8625
rect 15381 8616 15393 8619
rect 15160 8588 15393 8616
rect 15160 8576 15166 8588
rect 15381 8585 15393 8588
rect 15427 8585 15439 8619
rect 15381 8579 15439 8585
rect 16206 8576 16212 8628
rect 16264 8616 16270 8628
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 16264 8588 17417 8616
rect 16264 8576 16270 8588
rect 17405 8585 17417 8588
rect 17451 8585 17463 8619
rect 17405 8579 17463 8585
rect 3878 8508 3884 8560
rect 3936 8548 3942 8560
rect 4154 8548 4160 8560
rect 3936 8520 4160 8548
rect 3936 8508 3942 8520
rect 4154 8508 4160 8520
rect 4212 8548 4218 8560
rect 8711 8551 8769 8557
rect 8711 8548 8723 8551
rect 4212 8520 8723 8548
rect 4212 8508 4218 8520
rect 8711 8517 8723 8520
rect 8757 8517 8769 8551
rect 8711 8511 8769 8517
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 11287 8551 11345 8557
rect 11287 8548 11299 8551
rect 9272 8520 11299 8548
rect 9272 8508 9278 8520
rect 11287 8517 11299 8520
rect 11333 8517 11345 8551
rect 11287 8511 11345 8517
rect 11422 8508 11428 8560
rect 11480 8548 11486 8560
rect 13081 8551 13139 8557
rect 13081 8548 13093 8551
rect 11480 8520 13093 8548
rect 11480 8508 11486 8520
rect 13081 8517 13093 8520
rect 13127 8517 13139 8551
rect 13081 8511 13139 8517
rect 2038 8440 2044 8492
rect 2096 8480 2102 8492
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 2096 8452 9413 8480
rect 2096 8440 2102 8452
rect 9401 8449 9413 8452
rect 9447 8480 9459 8483
rect 9490 8480 9496 8492
rect 9447 8452 9496 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 9674 8480 9680 8492
rect 9635 8452 9680 8480
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8480 10379 8483
rect 12529 8483 12587 8489
rect 12529 8480 12541 8483
rect 10367 8452 12541 8480
rect 10367 8449 10379 8452
rect 10321 8443 10379 8449
rect 12529 8449 12541 8452
rect 12575 8480 12587 8483
rect 13170 8480 13176 8492
rect 12575 8452 13176 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 13170 8440 13176 8452
rect 13228 8480 13234 8492
rect 14369 8483 14427 8489
rect 14369 8480 14381 8483
rect 13228 8452 14381 8480
rect 13228 8440 13234 8452
rect 14369 8449 14381 8452
rect 14415 8480 14427 8483
rect 15013 8483 15071 8489
rect 15013 8480 15025 8483
rect 14415 8452 15025 8480
rect 14415 8449 14427 8452
rect 14369 8443 14427 8449
rect 15013 8449 15025 8452
rect 15059 8449 15071 8483
rect 16482 8480 16488 8492
rect 16443 8452 16488 8480
rect 15013 8443 15071 8449
rect 16482 8440 16488 8452
rect 16540 8440 16546 8492
rect 17420 8480 17448 8579
rect 18141 8483 18199 8489
rect 18141 8480 18153 8483
rect 17420 8452 18153 8480
rect 18141 8449 18153 8452
rect 18187 8449 18199 8483
rect 18414 8480 18420 8492
rect 18375 8452 18420 8480
rect 18141 8443 18199 8449
rect 18414 8440 18420 8452
rect 18472 8440 18478 8492
rect 4522 8372 4528 8424
rect 4580 8412 4586 8424
rect 4985 8415 5043 8421
rect 4985 8412 4997 8415
rect 4580 8384 4997 8412
rect 4580 8372 4586 8384
rect 4985 8381 4997 8384
rect 5031 8412 5043 8415
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 5031 8384 5181 8412
rect 5031 8381 5043 8384
rect 4985 8375 5043 8381
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 5169 8375 5227 8381
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 8640 8415 8698 8421
rect 8640 8381 8652 8415
rect 8686 8412 8698 8415
rect 9030 8412 9036 8424
rect 8686 8384 9036 8412
rect 8686 8381 8698 8384
rect 8640 8375 8698 8381
rect 9030 8372 9036 8384
rect 9088 8372 9094 8424
rect 10870 8372 10876 8424
rect 10928 8412 10934 8424
rect 11184 8415 11242 8421
rect 11184 8412 11196 8415
rect 10928 8384 11196 8412
rect 10928 8372 10934 8384
rect 11184 8381 11196 8384
rect 11230 8412 11242 8415
rect 11609 8415 11667 8421
rect 11609 8412 11621 8415
rect 11230 8384 11621 8412
rect 11230 8381 11242 8384
rect 11184 8375 11242 8381
rect 11609 8381 11621 8384
rect 11655 8381 11667 8415
rect 11609 8375 11667 8381
rect 18874 8372 18880 8424
rect 18932 8412 18938 8424
rect 19664 8415 19722 8421
rect 19664 8412 19676 8415
rect 18932 8384 19676 8412
rect 18932 8372 18938 8384
rect 19664 8381 19676 8384
rect 19710 8412 19722 8415
rect 20073 8415 20131 8421
rect 20073 8412 20085 8415
rect 19710 8384 20085 8412
rect 19710 8381 19722 8384
rect 19664 8375 19722 8381
rect 20073 8381 20085 8384
rect 20119 8381 20131 8415
rect 20073 8375 20131 8381
rect 5074 8344 5080 8356
rect 5035 8316 5080 8344
rect 5074 8304 5080 8316
rect 5132 8304 5138 8356
rect 7146 8347 7204 8353
rect 7146 8344 7158 8347
rect 6656 8316 7158 8344
rect 6656 8288 6684 8316
rect 7146 8313 7158 8316
rect 7192 8344 7204 8347
rect 7282 8344 7288 8356
rect 7192 8316 7288 8344
rect 7192 8313 7204 8316
rect 7146 8307 7204 8313
rect 7282 8304 7288 8316
rect 7340 8344 7346 8356
rect 8018 8344 8024 8356
rect 7340 8316 8024 8344
rect 7340 8304 7346 8316
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 9766 8344 9772 8356
rect 9727 8316 9772 8344
rect 9766 8304 9772 8316
rect 9824 8344 9830 8356
rect 10134 8344 10140 8356
rect 9824 8316 10140 8344
rect 9824 8304 9830 8316
rect 10134 8304 10140 8316
rect 10192 8344 10198 8356
rect 10597 8347 10655 8353
rect 10597 8344 10609 8347
rect 10192 8316 10609 8344
rect 10192 8304 10198 8316
rect 10597 8313 10609 8316
rect 10643 8313 10655 8347
rect 10597 8307 10655 8313
rect 12618 8304 12624 8356
rect 12676 8344 12682 8356
rect 14090 8344 14096 8356
rect 12676 8316 12721 8344
rect 14051 8316 14096 8344
rect 12676 8304 12682 8316
rect 14090 8304 14096 8316
rect 14148 8304 14154 8356
rect 14185 8347 14243 8353
rect 14185 8313 14197 8347
rect 14231 8313 14243 8347
rect 14185 8307 14243 8313
rect 16301 8347 16359 8353
rect 16301 8313 16313 8347
rect 16347 8344 16359 8347
rect 16577 8347 16635 8353
rect 16577 8344 16589 8347
rect 16347 8316 16589 8344
rect 16347 8313 16359 8316
rect 16301 8307 16359 8313
rect 16577 8313 16589 8316
rect 16623 8344 16635 8347
rect 16942 8344 16948 8356
rect 16623 8316 16948 8344
rect 16623 8313 16635 8316
rect 16577 8307 16635 8313
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 4065 8279 4123 8285
rect 4065 8276 4077 8279
rect 4028 8248 4077 8276
rect 4028 8236 4034 8248
rect 4065 8245 4077 8248
rect 4111 8245 4123 8279
rect 6638 8276 6644 8288
rect 6599 8248 6644 8276
rect 4065 8239 4123 8245
rect 6638 8236 6644 8248
rect 6696 8236 6702 8288
rect 8481 8279 8539 8285
rect 8481 8245 8493 8279
rect 8527 8276 8539 8279
rect 8662 8276 8668 8288
rect 8527 8248 8668 8276
rect 8527 8245 8539 8248
rect 8481 8239 8539 8245
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 11054 8276 11060 8288
rect 11015 8248 11060 8276
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 11606 8236 11612 8288
rect 11664 8276 11670 8288
rect 11977 8279 12035 8285
rect 11977 8276 11989 8279
rect 11664 8248 11989 8276
rect 11664 8236 11670 8248
rect 11977 8245 11989 8248
rect 12023 8245 12035 8279
rect 13906 8276 13912 8288
rect 13819 8248 13912 8276
rect 11977 8239 12035 8245
rect 13906 8236 13912 8248
rect 13964 8276 13970 8288
rect 14200 8276 14228 8307
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 17129 8347 17187 8353
rect 17129 8313 17141 8347
rect 17175 8344 17187 8347
rect 17402 8344 17408 8356
rect 17175 8316 17408 8344
rect 17175 8313 17187 8316
rect 17129 8307 17187 8313
rect 17402 8304 17408 8316
rect 17460 8304 17466 8356
rect 17862 8344 17868 8356
rect 17823 8316 17868 8344
rect 17862 8304 17868 8316
rect 17920 8304 17926 8356
rect 18230 8344 18236 8356
rect 18191 8316 18236 8344
rect 18230 8304 18236 8316
rect 18288 8304 18294 8356
rect 19751 8347 19809 8353
rect 19751 8313 19763 8347
rect 19797 8344 19809 8347
rect 21450 8344 21456 8356
rect 19797 8316 21456 8344
rect 19797 8313 19809 8316
rect 19751 8307 19809 8313
rect 21450 8304 21456 8316
rect 21508 8304 21514 8356
rect 15930 8276 15936 8288
rect 13964 8248 14228 8276
rect 15891 8248 15936 8276
rect 13964 8236 13970 8248
rect 15930 8236 15936 8248
rect 15988 8236 15994 8288
rect 19150 8276 19156 8288
rect 19111 8248 19156 8276
rect 19150 8236 19156 8248
rect 19208 8236 19214 8288
rect 1104 8186 20884 8208
rect 1104 8134 8315 8186
rect 8367 8134 8379 8186
rect 8431 8134 8443 8186
rect 8495 8134 8507 8186
rect 8559 8134 15648 8186
rect 15700 8134 15712 8186
rect 15764 8134 15776 8186
rect 15828 8134 15840 8186
rect 15892 8134 20884 8186
rect 1104 8112 20884 8134
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 9766 8072 9772 8084
rect 8803 8044 9772 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 10042 8072 10048 8084
rect 10003 8044 10048 8072
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 15930 8032 15936 8084
rect 15988 8072 15994 8084
rect 16209 8075 16267 8081
rect 16209 8072 16221 8075
rect 15988 8044 16221 8072
rect 15988 8032 15994 8044
rect 16209 8041 16221 8044
rect 16255 8041 16267 8075
rect 16209 8035 16267 8041
rect 5899 8007 5957 8013
rect 5899 7973 5911 8007
rect 5945 8004 5957 8007
rect 6638 8004 6644 8016
rect 5945 7976 6644 8004
rect 5945 7973 5957 7976
rect 5899 7967 5957 7973
rect 6638 7964 6644 7976
rect 6696 8004 6702 8016
rect 6696 7976 6960 8004
rect 6696 7964 6702 7976
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4571 7840 5181 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 5169 7837 5181 7840
rect 5215 7868 5227 7871
rect 5258 7868 5264 7880
rect 5215 7840 5264 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5534 7868 5540 7880
rect 5495 7840 5540 7868
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 4433 7735 4491 7741
rect 4433 7701 4445 7735
rect 4479 7732 4491 7735
rect 5166 7732 5172 7744
rect 4479 7704 5172 7732
rect 4479 7701 4491 7704
rect 4433 7695 4491 7701
rect 5166 7692 5172 7704
rect 5224 7692 5230 7744
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 6932 7741 6960 7976
rect 8018 7964 8024 8016
rect 8076 8004 8082 8016
rect 8158 8007 8216 8013
rect 8158 8004 8170 8007
rect 8076 7976 8170 8004
rect 8076 7964 8082 7976
rect 8158 7973 8170 7976
rect 8204 7973 8216 8007
rect 8158 7967 8216 7973
rect 11606 7964 11612 8016
rect 11664 8004 11670 8016
rect 11930 8007 11988 8013
rect 11930 8004 11942 8007
rect 11664 7976 11942 8004
rect 11664 7964 11670 7976
rect 11930 7973 11942 7976
rect 11976 7973 11988 8007
rect 13541 8007 13599 8013
rect 13541 8004 13553 8007
rect 11930 7967 11988 7973
rect 13188 7976 13553 8004
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 7926 7936 7932 7948
rect 7883 7908 7932 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 7926 7896 7932 7908
rect 7984 7896 7990 7948
rect 13188 7945 13216 7976
rect 13541 7973 13553 7976
rect 13587 8004 13599 8007
rect 13906 8004 13912 8016
rect 13587 7976 13912 8004
rect 13587 7973 13599 7976
rect 13541 7967 13599 7973
rect 13906 7964 13912 7976
rect 13964 7964 13970 8016
rect 15651 8007 15709 8013
rect 15651 7973 15663 8007
rect 15697 8004 15709 8007
rect 16022 8004 16028 8016
rect 15697 7976 16028 8004
rect 15697 7973 15709 7976
rect 15651 7967 15709 7973
rect 16022 7964 16028 7976
rect 16080 7964 16086 8016
rect 16224 8004 16252 8035
rect 16298 8032 16304 8084
rect 16356 8072 16362 8084
rect 16853 8075 16911 8081
rect 16853 8072 16865 8075
rect 16356 8044 16865 8072
rect 16356 8032 16362 8044
rect 16853 8041 16865 8044
rect 16899 8041 16911 8075
rect 16853 8035 16911 8041
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 18049 8075 18107 8081
rect 18049 8072 18061 8075
rect 17000 8044 18061 8072
rect 17000 8032 17006 8044
rect 18049 8041 18061 8044
rect 18095 8072 18107 8075
rect 18230 8072 18236 8084
rect 18095 8044 18236 8072
rect 18095 8041 18107 8044
rect 18049 8035 18107 8041
rect 18230 8032 18236 8044
rect 18288 8032 18294 8084
rect 16574 8004 16580 8016
rect 16224 7976 16580 8004
rect 16574 7964 16580 7976
rect 16632 8004 16638 8016
rect 17221 8007 17279 8013
rect 17221 8004 17233 8007
rect 16632 7976 17233 8004
rect 16632 7964 16638 7976
rect 17221 7973 17233 7976
rect 17267 8004 17279 8007
rect 17310 8004 17316 8016
rect 17267 7976 17316 8004
rect 17267 7973 17279 7976
rect 17221 7967 17279 7973
rect 17310 7964 17316 7976
rect 17368 7964 17374 8016
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7936 12587 7939
rect 13173 7939 13231 7945
rect 13173 7936 13185 7939
rect 12575 7908 13185 7936
rect 12575 7905 12587 7908
rect 12529 7899 12587 7905
rect 13173 7905 13185 7908
rect 13219 7905 13231 7939
rect 18598 7936 18604 7948
rect 18559 7908 18604 7936
rect 13173 7899 13231 7905
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 9766 7868 9772 7880
rect 9723 7840 9772 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 9766 7828 9772 7840
rect 9824 7868 9830 7880
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 9824 7840 10885 7868
rect 9824 7828 9830 7840
rect 10873 7837 10885 7840
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 11514 7828 11520 7880
rect 11572 7868 11578 7880
rect 11609 7871 11667 7877
rect 11609 7868 11621 7871
rect 11572 7840 11621 7868
rect 11572 7828 11578 7840
rect 11609 7837 11621 7840
rect 11655 7837 11667 7871
rect 13446 7868 13452 7880
rect 13407 7840 13452 7868
rect 11609 7831 11667 7837
rect 13446 7828 13452 7840
rect 13504 7828 13510 7880
rect 13538 7828 13544 7880
rect 13596 7868 13602 7880
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13596 7840 13737 7868
rect 13596 7828 13602 7840
rect 13725 7837 13737 7840
rect 13771 7837 13783 7871
rect 15286 7868 15292 7880
rect 15247 7840 15292 7868
rect 13725 7831 13783 7837
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7868 17187 7871
rect 17218 7868 17224 7880
rect 17175 7840 17224 7868
rect 17175 7837 17187 7840
rect 17129 7831 17187 7837
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 17402 7868 17408 7880
rect 17363 7840 17408 7868
rect 17402 7828 17408 7840
rect 17460 7868 17466 7880
rect 18782 7868 18788 7880
rect 17460 7840 18788 7868
rect 17460 7828 17466 7840
rect 18782 7828 18788 7840
rect 18840 7828 18846 7880
rect 19610 7868 19616 7880
rect 19571 7840 19616 7868
rect 19610 7828 19616 7840
rect 19668 7828 19674 7880
rect 10597 7803 10655 7809
rect 10597 7769 10609 7803
rect 10643 7800 10655 7803
rect 12618 7800 12624 7812
rect 10643 7772 12624 7800
rect 10643 7769 10655 7772
rect 10597 7763 10655 7769
rect 12618 7760 12624 7772
rect 12676 7800 12682 7812
rect 12805 7803 12863 7809
rect 12805 7800 12817 7803
rect 12676 7772 12817 7800
rect 12676 7760 12682 7772
rect 12805 7769 12817 7772
rect 12851 7769 12863 7803
rect 12805 7763 12863 7769
rect 6457 7735 6515 7741
rect 6457 7732 6469 7735
rect 5408 7704 6469 7732
rect 5408 7692 5414 7704
rect 6457 7701 6469 7704
rect 6503 7701 6515 7735
rect 6457 7695 6515 7701
rect 6917 7735 6975 7741
rect 6917 7701 6929 7735
rect 6963 7732 6975 7735
rect 7190 7732 7196 7744
rect 6963 7704 7196 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 7561 7735 7619 7741
rect 7561 7701 7573 7735
rect 7607 7732 7619 7735
rect 8202 7732 8208 7744
rect 7607 7704 8208 7732
rect 7607 7701 7619 7704
rect 7561 7695 7619 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 9033 7735 9091 7741
rect 9033 7732 9045 7735
rect 8720 7704 9045 7732
rect 8720 7692 8726 7704
rect 9033 7701 9045 7704
rect 9079 7701 9091 7735
rect 9398 7732 9404 7744
rect 9359 7704 9404 7732
rect 9033 7695 9091 7701
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 11514 7732 11520 7744
rect 11475 7704 11520 7732
rect 11514 7692 11520 7704
rect 11572 7692 11578 7744
rect 12342 7692 12348 7744
rect 12400 7732 12406 7744
rect 13630 7732 13636 7744
rect 12400 7704 13636 7732
rect 12400 7692 12406 7704
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 14461 7735 14519 7741
rect 14461 7701 14473 7735
rect 14507 7732 14519 7735
rect 15102 7732 15108 7744
rect 14507 7704 15108 7732
rect 14507 7701 14519 7704
rect 14461 7695 14519 7701
rect 15102 7692 15108 7704
rect 15160 7692 15166 7744
rect 16482 7732 16488 7744
rect 16443 7704 16488 7732
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 18138 7692 18144 7744
rect 18196 7732 18202 7744
rect 18739 7735 18797 7741
rect 18739 7732 18751 7735
rect 18196 7704 18751 7732
rect 18196 7692 18202 7704
rect 18739 7701 18751 7704
rect 18785 7701 18797 7735
rect 18739 7695 18797 7701
rect 1104 7642 20884 7664
rect 1104 7590 4648 7642
rect 4700 7590 4712 7642
rect 4764 7590 4776 7642
rect 4828 7590 4840 7642
rect 4892 7590 11982 7642
rect 12034 7590 12046 7642
rect 12098 7590 12110 7642
rect 12162 7590 12174 7642
rect 12226 7590 19315 7642
rect 19367 7590 19379 7642
rect 19431 7590 19443 7642
rect 19495 7590 19507 7642
rect 19559 7590 20884 7642
rect 1104 7568 20884 7590
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 4479 7500 6684 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 1670 7460 1676 7472
rect 1583 7432 1676 7460
rect 1670 7420 1676 7432
rect 1728 7460 1734 7472
rect 6656 7469 6684 7500
rect 9306 7488 9312 7540
rect 9364 7528 9370 7540
rect 10689 7531 10747 7537
rect 10689 7528 10701 7531
rect 9364 7500 10701 7528
rect 9364 7488 9370 7500
rect 10689 7497 10701 7500
rect 10735 7497 10747 7531
rect 10689 7491 10747 7497
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 12986 7528 12992 7540
rect 12299 7500 12992 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 13630 7528 13636 7540
rect 13591 7500 13636 7528
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 16942 7488 16948 7540
rect 17000 7528 17006 7540
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 17000 7500 17049 7528
rect 17000 7488 17006 7500
rect 17037 7497 17049 7500
rect 17083 7497 17095 7531
rect 17310 7528 17316 7540
rect 17271 7500 17316 7528
rect 17037 7491 17095 7497
rect 17310 7488 17316 7500
rect 17368 7488 17374 7540
rect 17494 7488 17500 7540
rect 17552 7528 17558 7540
rect 18233 7531 18291 7537
rect 18233 7528 18245 7531
rect 17552 7500 18245 7528
rect 17552 7488 17558 7500
rect 18233 7497 18245 7500
rect 18279 7497 18291 7531
rect 18233 7491 18291 7497
rect 6641 7463 6699 7469
rect 1728 7432 5948 7460
rect 1728 7420 1734 7432
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4387 7364 4445 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 5258 7392 5264 7404
rect 5219 7364 5264 7392
rect 4433 7355 4491 7361
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5920 7401 5948 7432
rect 6641 7429 6653 7463
rect 6687 7460 6699 7463
rect 8478 7460 8484 7472
rect 6687 7432 8484 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 8478 7420 8484 7432
rect 8536 7460 8542 7472
rect 9122 7460 9128 7472
rect 8536 7432 9128 7460
rect 8536 7420 8542 7432
rect 9122 7420 9128 7432
rect 9180 7420 9186 7472
rect 10870 7420 10876 7472
rect 10928 7460 10934 7472
rect 10928 7432 19196 7460
rect 10928 7420 10934 7432
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 9858 7392 9864 7404
rect 5951 7364 9864 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7392 15347 7395
rect 16117 7395 16175 7401
rect 16117 7392 16129 7395
rect 15335 7364 16129 7392
rect 15335 7361 15347 7364
rect 15289 7355 15347 7361
rect 16117 7361 16129 7364
rect 16163 7392 16175 7395
rect 16482 7392 16488 7404
rect 16163 7364 16488 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 17770 7392 17776 7404
rect 17731 7364 17776 7392
rect 17770 7352 17776 7364
rect 17828 7352 17834 7404
rect 3513 7327 3571 7333
rect 3513 7293 3525 7327
rect 3559 7324 3571 7327
rect 3694 7324 3700 7336
rect 3559 7296 3700 7324
rect 3559 7293 3571 7296
rect 3513 7287 3571 7293
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 7466 7324 7472 7336
rect 7427 7296 7472 7324
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 8202 7324 8208 7336
rect 8163 7296 8208 7324
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8478 7324 8484 7336
rect 8439 7296 8484 7324
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 8662 7324 8668 7336
rect 8623 7296 8668 7324
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 8754 7284 8760 7336
rect 8812 7324 8818 7336
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 8812 7296 9781 7324
rect 8812 7284 8818 7296
rect 9769 7293 9781 7296
rect 9815 7324 9827 7327
rect 9950 7324 9956 7336
rect 9815 7296 9956 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 11606 7324 11612 7336
rect 10888 7296 11612 7324
rect 4709 7259 4767 7265
rect 4709 7225 4721 7259
rect 4755 7256 4767 7259
rect 5350 7256 5356 7268
rect 4755 7228 5356 7256
rect 4755 7225 4767 7228
rect 4709 7219 4767 7225
rect 5350 7216 5356 7228
rect 5408 7216 5414 7268
rect 6273 7259 6331 7265
rect 6273 7225 6285 7259
rect 6319 7256 6331 7259
rect 7190 7256 7196 7268
rect 6319 7228 7196 7256
rect 6319 7225 6331 7228
rect 6273 7219 6331 7225
rect 7190 7216 7196 7228
rect 7248 7256 7254 7268
rect 9217 7259 9275 7265
rect 9217 7256 9229 7259
rect 7248 7228 9229 7256
rect 7248 7216 7254 7228
rect 9217 7225 9229 7228
rect 9263 7256 9275 7259
rect 9585 7259 9643 7265
rect 9585 7256 9597 7259
rect 9263 7228 9597 7256
rect 9263 7225 9275 7228
rect 9217 7219 9275 7225
rect 9585 7225 9597 7228
rect 9631 7256 9643 7259
rect 10042 7256 10048 7268
rect 9631 7228 10048 7256
rect 9631 7225 9643 7228
rect 9585 7219 9643 7225
rect 10042 7216 10048 7228
rect 10100 7265 10106 7268
rect 10100 7259 10148 7265
rect 10100 7225 10102 7259
rect 10136 7256 10148 7259
rect 10888 7256 10916 7296
rect 11606 7284 11612 7296
rect 11664 7284 11670 7336
rect 12575 7327 12633 7333
rect 12575 7293 12587 7327
rect 12621 7324 12633 7327
rect 13446 7324 13452 7336
rect 12621 7296 13452 7324
rect 12621 7293 12633 7296
rect 12575 7287 12633 7293
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 13630 7284 13636 7336
rect 13688 7324 13694 7336
rect 13817 7327 13875 7333
rect 13817 7324 13829 7327
rect 13688 7296 13829 7324
rect 13688 7284 13694 7296
rect 13817 7293 13829 7296
rect 13863 7324 13875 7327
rect 13998 7324 14004 7336
rect 13863 7296 14004 7324
rect 13863 7293 13875 7296
rect 13817 7287 13875 7293
rect 13998 7284 14004 7296
rect 14056 7284 14062 7336
rect 14277 7327 14335 7333
rect 14277 7293 14289 7327
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 11977 7259 12035 7265
rect 11977 7256 11989 7259
rect 10136 7228 10916 7256
rect 10980 7228 11989 7256
rect 10136 7225 10148 7228
rect 10100 7219 10148 7225
rect 10100 7216 10106 7219
rect 2038 7188 2044 7200
rect 1999 7160 2044 7188
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 2406 7188 2412 7200
rect 2367 7160 2412 7188
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 2682 7188 2688 7200
rect 2643 7160 2688 7188
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 3050 7188 3056 7200
rect 3011 7160 3056 7188
rect 3050 7148 3056 7160
rect 3108 7148 3114 7200
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7188 5135 7191
rect 6086 7188 6092 7200
rect 5123 7160 6092 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 6086 7148 6092 7160
rect 6144 7148 6150 7200
rect 7377 7191 7435 7197
rect 7377 7157 7389 7191
rect 7423 7188 7435 7191
rect 7466 7188 7472 7200
rect 7423 7160 7472 7188
rect 7423 7157 7435 7160
rect 7377 7151 7435 7157
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 7745 7191 7803 7197
rect 7745 7157 7757 7191
rect 7791 7188 7803 7191
rect 7926 7188 7932 7200
rect 7791 7160 7932 7188
rect 7791 7157 7803 7160
rect 7745 7151 7803 7157
rect 7926 7148 7932 7160
rect 7984 7148 7990 7200
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 10980 7197 11008 7228
rect 11977 7225 11989 7228
rect 12023 7225 12035 7259
rect 14292 7256 14320 7287
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 14700 7296 14745 7324
rect 14700 7284 14706 7296
rect 15102 7284 15108 7336
rect 15160 7324 15166 7336
rect 15197 7327 15255 7333
rect 15197 7324 15209 7327
rect 15160 7296 15209 7324
rect 15160 7284 15166 7296
rect 15197 7293 15209 7296
rect 15243 7324 15255 7327
rect 16206 7324 16212 7336
rect 15243 7296 16212 7324
rect 15243 7293 15255 7296
rect 15197 7287 15255 7293
rect 16206 7284 16212 7296
rect 16264 7284 16270 7336
rect 17788 7324 17816 7352
rect 19168 7333 19196 7432
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17788 7296 18061 7324
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 19153 7327 19211 7333
rect 19153 7293 19165 7327
rect 19199 7324 19211 7327
rect 19705 7327 19763 7333
rect 19705 7324 19717 7327
rect 19199 7296 19717 7324
rect 19199 7293 19211 7296
rect 19153 7287 19211 7293
rect 19705 7293 19717 7296
rect 19751 7293 19763 7327
rect 19705 7287 19763 7293
rect 16438 7259 16496 7265
rect 16438 7256 16450 7259
rect 11977 7219 12035 7225
rect 13280 7228 14320 7256
rect 16040 7228 16450 7256
rect 10965 7191 11023 7197
rect 10965 7188 10977 7191
rect 10928 7160 10977 7188
rect 10928 7148 10934 7160
rect 10965 7157 10977 7160
rect 11011 7157 11023 7191
rect 10965 7151 11023 7157
rect 12710 7148 12716 7200
rect 12768 7188 12774 7200
rect 13280 7197 13308 7228
rect 16040 7200 16068 7228
rect 16438 7225 16450 7228
rect 16484 7225 16496 7259
rect 16438 7219 16496 7225
rect 18598 7216 18604 7268
rect 18656 7256 18662 7268
rect 18693 7259 18751 7265
rect 18693 7256 18705 7259
rect 18656 7228 18705 7256
rect 18656 7216 18662 7228
rect 18693 7225 18705 7228
rect 18739 7256 18751 7259
rect 19794 7256 19800 7268
rect 18739 7228 19800 7256
rect 18739 7225 18751 7228
rect 18693 7219 18751 7225
rect 19794 7216 19800 7228
rect 19852 7216 19858 7268
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 12768 7160 13277 7188
rect 12768 7148 12774 7160
rect 13265 7157 13277 7160
rect 13311 7157 13323 7191
rect 13265 7151 13323 7157
rect 15657 7191 15715 7197
rect 15657 7157 15669 7191
rect 15703 7188 15715 7191
rect 16022 7188 16028 7200
rect 15703 7160 16028 7188
rect 15703 7157 15715 7160
rect 15657 7151 15715 7157
rect 16022 7148 16028 7160
rect 16080 7148 16086 7200
rect 18966 7148 18972 7200
rect 19024 7188 19030 7200
rect 19337 7191 19395 7197
rect 19337 7188 19349 7191
rect 19024 7160 19349 7188
rect 19024 7148 19030 7160
rect 19337 7157 19349 7160
rect 19383 7157 19395 7191
rect 19337 7151 19395 7157
rect 1104 7098 20884 7120
rect 1104 7046 8315 7098
rect 8367 7046 8379 7098
rect 8431 7046 8443 7098
rect 8495 7046 8507 7098
rect 8559 7046 15648 7098
rect 15700 7046 15712 7098
rect 15764 7046 15776 7098
rect 15828 7046 15840 7098
rect 15892 7046 20884 7098
rect 1104 7024 20884 7046
rect 4525 6987 4583 6993
rect 4525 6953 4537 6987
rect 4571 6984 4583 6987
rect 5077 6987 5135 6993
rect 5077 6984 5089 6987
rect 4571 6956 5089 6984
rect 4571 6953 4583 6956
rect 4525 6947 4583 6953
rect 5077 6953 5089 6956
rect 5123 6984 5135 6987
rect 5534 6984 5540 6996
rect 5123 6956 5540 6984
rect 5123 6953 5135 6956
rect 5077 6947 5135 6953
rect 5534 6944 5540 6956
rect 5592 6944 5598 6996
rect 9766 6984 9772 6996
rect 9727 6956 9772 6984
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 11514 6944 11520 6996
rect 11572 6984 11578 6996
rect 12069 6987 12127 6993
rect 12069 6984 12081 6987
rect 11572 6956 12081 6984
rect 11572 6944 11578 6956
rect 12069 6953 12081 6956
rect 12115 6953 12127 6987
rect 12069 6947 12127 6953
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 14645 6987 14703 6993
rect 14645 6984 14657 6987
rect 13504 6956 14657 6984
rect 13504 6944 13510 6956
rect 14645 6953 14657 6956
rect 14691 6953 14703 6987
rect 14645 6947 14703 6953
rect 15105 6987 15163 6993
rect 15105 6953 15117 6987
rect 15151 6984 15163 6987
rect 15286 6984 15292 6996
rect 15151 6956 15292 6984
rect 15151 6953 15163 6956
rect 15105 6947 15163 6953
rect 15286 6944 15292 6956
rect 15344 6984 15350 6996
rect 15381 6987 15439 6993
rect 15381 6984 15393 6987
rect 15344 6956 15393 6984
rect 15344 6944 15350 6956
rect 15381 6953 15393 6956
rect 15427 6953 15439 6987
rect 15381 6947 15439 6953
rect 17218 6944 17224 6996
rect 17276 6984 17282 6996
rect 17405 6987 17463 6993
rect 17405 6984 17417 6987
rect 17276 6956 17417 6984
rect 17276 6944 17282 6956
rect 17405 6953 17417 6956
rect 17451 6953 17463 6987
rect 17405 6947 17463 6953
rect 8754 6916 8760 6928
rect 6196 6888 8524 6916
rect 8715 6888 8760 6916
rect 6196 6860 6224 6888
rect 1464 6851 1522 6857
rect 1464 6817 1476 6851
rect 1510 6848 1522 6851
rect 1670 6848 1676 6860
rect 1510 6820 1676 6848
rect 1510 6817 1522 6820
rect 1464 6811 1522 6817
rect 1670 6808 1676 6820
rect 1728 6808 1734 6860
rect 5258 6848 5264 6860
rect 5219 6820 5264 6848
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 5718 6848 5724 6860
rect 5679 6820 5724 6848
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 5994 6848 6000 6860
rect 5955 6820 6000 6848
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 6178 6848 6184 6860
rect 6139 6820 6184 6848
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 7466 6848 7472 6860
rect 7427 6820 7472 6848
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7926 6848 7932 6860
rect 7887 6820 7932 6848
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 8496 6857 8524 6888
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 13909 6919 13967 6925
rect 13909 6916 13921 6919
rect 9968 6888 11928 6916
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6817 8171 6851
rect 8113 6811 8171 6817
rect 8481 6851 8539 6857
rect 8481 6817 8493 6851
rect 8527 6848 8539 6851
rect 8662 6848 8668 6860
rect 8527 6820 8668 6848
rect 8527 6817 8539 6820
rect 8481 6811 8539 6817
rect 8018 6780 8024 6792
rect 4126 6752 8024 6780
rect 2547 6715 2605 6721
rect 2547 6681 2559 6715
rect 2593 6712 2605 6715
rect 4126 6712 4154 6752
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 2593 6684 4154 6712
rect 2593 6681 2605 6684
rect 2547 6675 2605 6681
rect 4522 6672 4528 6724
rect 4580 6712 4586 6724
rect 6730 6712 6736 6724
rect 4580 6684 6736 6712
rect 4580 6672 4586 6684
rect 6730 6672 6736 6684
rect 6788 6712 6794 6724
rect 6825 6715 6883 6721
rect 6825 6712 6837 6715
rect 6788 6684 6837 6712
rect 6788 6672 6794 6684
rect 6825 6681 6837 6684
rect 6871 6681 6883 6715
rect 6825 6675 6883 6681
rect 7834 6672 7840 6724
rect 7892 6712 7898 6724
rect 8128 6712 8156 6811
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 9030 6808 9036 6860
rect 9088 6848 9094 6860
rect 9968 6857 9996 6888
rect 11900 6860 11928 6888
rect 12728 6888 13921 6916
rect 12728 6860 12756 6888
rect 13909 6885 13921 6888
rect 13955 6916 13967 6919
rect 17770 6916 17776 6928
rect 13955 6888 15792 6916
rect 17731 6888 17776 6916
rect 13955 6885 13967 6888
rect 13909 6879 13967 6885
rect 15764 6860 15792 6888
rect 17770 6876 17776 6888
rect 17828 6876 17834 6928
rect 18325 6919 18383 6925
rect 18325 6885 18337 6919
rect 18371 6916 18383 6919
rect 18414 6916 18420 6928
rect 18371 6888 18420 6916
rect 18371 6885 18383 6888
rect 18325 6879 18383 6885
rect 18414 6876 18420 6888
rect 18472 6876 18478 6928
rect 9493 6851 9551 6857
rect 9493 6848 9505 6851
rect 9088 6820 9505 6848
rect 9088 6808 9094 6820
rect 9493 6817 9505 6820
rect 9539 6848 9551 6851
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9539 6820 9965 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 9953 6817 9965 6820
rect 9999 6817 10011 6851
rect 10410 6848 10416 6860
rect 10371 6820 10416 6848
rect 9953 6811 10011 6817
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 10686 6848 10692 6860
rect 10647 6820 10692 6848
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 10870 6848 10876 6860
rect 10783 6820 10876 6848
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 11882 6848 11888 6860
rect 11795 6820 11888 6848
rect 11882 6808 11888 6820
rect 11940 6848 11946 6860
rect 12253 6851 12311 6857
rect 12253 6848 12265 6851
rect 11940 6820 12265 6848
rect 11940 6808 11946 6820
rect 12253 6817 12265 6820
rect 12299 6848 12311 6851
rect 12342 6848 12348 6860
rect 12299 6820 12348 6848
rect 12299 6817 12311 6820
rect 12253 6811 12311 6817
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 12710 6848 12716 6860
rect 12671 6820 12716 6848
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 12894 6848 12900 6860
rect 12855 6820 12900 6848
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13173 6851 13231 6857
rect 13173 6817 13185 6851
rect 13219 6817 13231 6851
rect 13173 6811 13231 6817
rect 14369 6851 14427 6857
rect 14369 6817 14381 6851
rect 14415 6848 14427 6851
rect 14642 6848 14648 6860
rect 14415 6820 14648 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 8680 6780 8708 6808
rect 10888 6780 10916 6808
rect 11238 6780 11244 6792
rect 8680 6752 11244 6780
rect 11238 6740 11244 6752
rect 11296 6780 11302 6792
rect 11425 6783 11483 6789
rect 11425 6780 11437 6783
rect 11296 6752 11437 6780
rect 11296 6740 11302 6752
rect 11425 6749 11437 6752
rect 11471 6780 11483 6783
rect 13188 6780 13216 6811
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 15470 6848 15476 6860
rect 15431 6820 15476 6848
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 15746 6848 15752 6860
rect 15659 6820 15752 6848
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 16117 6851 16175 6857
rect 16117 6848 16129 6851
rect 15988 6820 16129 6848
rect 15988 6808 15994 6820
rect 16117 6817 16129 6820
rect 16163 6817 16175 6851
rect 16117 6811 16175 6817
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 16485 6851 16543 6857
rect 16485 6848 16497 6851
rect 16264 6820 16497 6848
rect 16264 6808 16270 6820
rect 16485 6817 16497 6820
rect 16531 6817 16543 6851
rect 16485 6811 16543 6817
rect 19058 6808 19064 6860
rect 19116 6848 19122 6860
rect 19153 6851 19211 6857
rect 19153 6848 19165 6851
rect 19116 6820 19165 6848
rect 19116 6808 19122 6820
rect 19153 6817 19165 6820
rect 19199 6817 19211 6851
rect 19153 6811 19211 6817
rect 11471 6752 13216 6780
rect 17681 6783 17739 6789
rect 11471 6749 11483 6752
rect 11425 6743 11483 6749
rect 17681 6749 17693 6783
rect 17727 6780 17739 6783
rect 18138 6780 18144 6792
rect 17727 6752 18144 6780
rect 17727 6749 17739 6752
rect 17681 6743 17739 6749
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 7892 6684 8156 6712
rect 7892 6672 7898 6684
rect 18598 6672 18604 6724
rect 18656 6712 18662 6724
rect 19337 6715 19395 6721
rect 19337 6712 19349 6715
rect 18656 6684 19349 6712
rect 18656 6672 18662 6684
rect 19337 6681 19349 6684
rect 19383 6681 19395 6715
rect 19337 6675 19395 6681
rect 106 6604 112 6656
rect 164 6644 170 6656
rect 1535 6647 1593 6653
rect 1535 6644 1547 6647
rect 164 6616 1547 6644
rect 164 6604 170 6616
rect 1535 6613 1547 6616
rect 1581 6613 1593 6647
rect 2130 6644 2136 6656
rect 2091 6616 2136 6644
rect 1535 6607 1593 6613
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 2869 6647 2927 6653
rect 2869 6644 2881 6647
rect 2832 6616 2881 6644
rect 2832 6604 2838 6616
rect 2869 6613 2881 6616
rect 2915 6613 2927 6647
rect 2869 6607 2927 6613
rect 3329 6647 3387 6653
rect 3329 6613 3341 6647
rect 3375 6644 3387 6647
rect 3602 6644 3608 6656
rect 3375 6616 3608 6644
rect 3375 6613 3387 6616
rect 3329 6607 3387 6613
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 4893 6647 4951 6653
rect 4893 6613 4905 6647
rect 4939 6644 4951 6647
rect 4982 6644 4988 6656
rect 4939 6616 4988 6644
rect 4939 6613 4951 6616
rect 4893 6607 4951 6613
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 9033 6647 9091 6653
rect 9033 6644 9045 6647
rect 6972 6616 9045 6644
rect 6972 6604 6978 6616
rect 9033 6613 9045 6616
rect 9079 6613 9091 6647
rect 9033 6607 9091 6613
rect 16206 6604 16212 6656
rect 16264 6644 16270 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 16264 6616 17049 6644
rect 16264 6604 16270 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 18690 6644 18696 6656
rect 18651 6616 18696 6644
rect 17037 6607 17095 6613
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 1104 6554 20884 6576
rect 1104 6502 4648 6554
rect 4700 6502 4712 6554
rect 4764 6502 4776 6554
rect 4828 6502 4840 6554
rect 4892 6502 11982 6554
rect 12034 6502 12046 6554
rect 12098 6502 12110 6554
rect 12162 6502 12174 6554
rect 12226 6502 19315 6554
rect 19367 6502 19379 6554
rect 19431 6502 19443 6554
rect 19495 6502 19507 6554
rect 19559 6502 20884 6554
rect 1104 6480 20884 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1854 6440 1860 6452
rect 1627 6412 1860 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1854 6400 1860 6412
rect 1912 6400 1918 6452
rect 6730 6400 6736 6452
rect 6788 6440 6794 6452
rect 6963 6443 7021 6449
rect 6963 6440 6975 6443
rect 6788 6412 6975 6440
rect 6788 6400 6794 6412
rect 6963 6409 6975 6412
rect 7009 6409 7021 6443
rect 6963 6403 7021 6409
rect 10502 6400 10508 6452
rect 10560 6440 10566 6452
rect 12575 6443 12633 6449
rect 12575 6440 12587 6443
rect 10560 6412 12587 6440
rect 10560 6400 10566 6412
rect 12575 6409 12587 6412
rect 12621 6409 12633 6443
rect 12575 6403 12633 6409
rect 15746 6400 15752 6452
rect 15804 6440 15810 6452
rect 16025 6443 16083 6449
rect 16025 6440 16037 6443
rect 15804 6412 16037 6440
rect 15804 6400 15810 6412
rect 16025 6409 16037 6412
rect 16071 6409 16083 6443
rect 16025 6403 16083 6409
rect 17129 6443 17187 6449
rect 17129 6409 17141 6443
rect 17175 6440 17187 6443
rect 17497 6443 17555 6449
rect 17497 6440 17509 6443
rect 17175 6412 17509 6440
rect 17175 6409 17187 6412
rect 17129 6403 17187 6409
rect 17497 6409 17509 6412
rect 17543 6440 17555 6443
rect 17770 6440 17776 6452
rect 17543 6412 17776 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 18690 6400 18696 6452
rect 18748 6440 18754 6452
rect 19751 6443 19809 6449
rect 19751 6440 19763 6443
rect 18748 6412 19763 6440
rect 18748 6400 18754 6412
rect 19751 6409 19763 6412
rect 19797 6409 19809 6443
rect 19751 6403 19809 6409
rect 7098 6372 7104 6384
rect 7059 6344 7104 6372
rect 7098 6332 7104 6344
rect 7156 6332 7162 6384
rect 7466 6332 7472 6384
rect 7524 6372 7530 6384
rect 9493 6375 9551 6381
rect 9493 6372 9505 6375
rect 7524 6344 9505 6372
rect 7524 6332 7530 6344
rect 9493 6341 9505 6344
rect 9539 6372 9551 6375
rect 9539 6344 9674 6372
rect 9539 6341 9551 6344
rect 9493 6335 9551 6341
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 6604 6276 7205 6304
rect 6604 6264 6610 6276
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 9214 6304 9220 6316
rect 8619 6276 9220 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6236 1458 6248
rect 1949 6239 2007 6245
rect 1949 6236 1961 6239
rect 1452 6208 1961 6236
rect 1452 6196 1458 6208
rect 1949 6205 1961 6208
rect 1995 6236 2007 6239
rect 2314 6236 2320 6248
rect 1995 6208 2320 6236
rect 1995 6205 2007 6208
rect 1949 6199 2007 6205
rect 2314 6196 2320 6208
rect 2372 6236 2378 6248
rect 2536 6239 2594 6245
rect 2536 6236 2548 6239
rect 2372 6208 2548 6236
rect 2372 6196 2378 6208
rect 2536 6205 2548 6208
rect 2582 6236 2594 6239
rect 2961 6239 3019 6245
rect 2961 6236 2973 6239
rect 2582 6208 2973 6236
rect 2582 6205 2594 6208
rect 2536 6199 2594 6205
rect 2961 6205 2973 6208
rect 3007 6205 3019 6239
rect 2961 6199 3019 6205
rect 3513 6239 3571 6245
rect 3513 6205 3525 6239
rect 3559 6236 3571 6239
rect 4249 6239 4307 6245
rect 4249 6236 4261 6239
rect 3559 6208 4261 6236
rect 3559 6205 3571 6208
rect 3513 6199 3571 6205
rect 4249 6205 4261 6208
rect 4295 6236 4307 6239
rect 4430 6236 4436 6248
rect 4295 6208 4436 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 5350 6236 5356 6248
rect 5311 6208 5356 6236
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6236 6883 6239
rect 6914 6236 6920 6248
rect 6871 6208 6920 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 7926 6236 7932 6248
rect 7024 6208 7932 6236
rect 4338 6168 4344 6180
rect 4299 6140 4344 6168
rect 4338 6128 4344 6140
rect 4396 6128 4402 6180
rect 4709 6171 4767 6177
rect 4709 6137 4721 6171
rect 4755 6168 4767 6171
rect 5718 6168 5724 6180
rect 4755 6140 5724 6168
rect 4755 6137 4767 6140
rect 4709 6131 4767 6137
rect 5718 6128 5724 6140
rect 5776 6168 5782 6180
rect 5905 6171 5963 6177
rect 5905 6168 5917 6171
rect 5776 6140 5917 6168
rect 5776 6128 5782 6140
rect 5905 6137 5917 6140
rect 5951 6168 5963 6171
rect 7024 6168 7052 6208
rect 7926 6196 7932 6208
rect 7984 6196 7990 6248
rect 9646 6236 9674 6344
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 11425 6375 11483 6381
rect 11425 6372 11437 6375
rect 11112 6344 11437 6372
rect 11112 6332 11118 6344
rect 11425 6341 11437 6344
rect 11471 6341 11483 6375
rect 11425 6335 11483 6341
rect 11974 6264 11980 6316
rect 12032 6304 12038 6316
rect 12710 6304 12716 6316
rect 12032 6276 12716 6304
rect 12032 6264 12038 6276
rect 12710 6264 12716 6276
rect 12768 6304 12774 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12768 6276 12909 6304
rect 12768 6264 12774 6276
rect 12897 6273 12909 6276
rect 12943 6304 12955 6307
rect 15381 6307 15439 6313
rect 12943 6276 14412 6304
rect 12943 6273 12955 6276
rect 12897 6267 12955 6273
rect 10045 6239 10103 6245
rect 10045 6236 10057 6239
rect 9646 6208 10057 6236
rect 10045 6205 10057 6208
rect 10091 6205 10103 6239
rect 10045 6199 10103 6205
rect 10410 6196 10416 6248
rect 10468 6236 10474 6248
rect 10505 6239 10563 6245
rect 10505 6236 10517 6239
rect 10468 6208 10517 6236
rect 10468 6196 10474 6208
rect 10505 6205 10517 6208
rect 10551 6205 10563 6239
rect 10505 6199 10563 6205
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6205 11115 6239
rect 11238 6236 11244 6248
rect 11199 6208 11244 6236
rect 11057 6199 11115 6205
rect 7558 6168 7564 6180
rect 5951 6140 7052 6168
rect 7519 6140 7564 6168
rect 5951 6137 5963 6140
rect 5905 6131 5963 6137
rect 7558 6128 7564 6140
rect 7616 6128 7622 6180
rect 8665 6171 8723 6177
rect 8665 6137 8677 6171
rect 8711 6168 8723 6171
rect 8754 6168 8760 6180
rect 8711 6140 8760 6168
rect 8711 6137 8723 6140
rect 8665 6131 8723 6137
rect 8754 6128 8760 6140
rect 8812 6128 8818 6180
rect 9214 6168 9220 6180
rect 9175 6140 9220 6168
rect 9214 6128 9220 6140
rect 9272 6128 9278 6180
rect 11072 6168 11100 6199
rect 11238 6196 11244 6208
rect 11296 6196 11302 6248
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 12472 6239 12530 6245
rect 12472 6236 12484 6239
rect 11848 6208 12484 6236
rect 11848 6196 11854 6208
rect 12472 6205 12484 6208
rect 12518 6236 12530 6239
rect 13265 6239 13323 6245
rect 13265 6236 13277 6239
rect 12518 6208 13277 6236
rect 12518 6205 12530 6208
rect 12472 6199 12530 6205
rect 13265 6205 13277 6208
rect 13311 6205 13323 6239
rect 13998 6236 14004 6248
rect 13959 6208 14004 6236
rect 13265 6199 13323 6205
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14384 6245 14412 6276
rect 15381 6273 15393 6307
rect 15427 6304 15439 6307
rect 16206 6304 16212 6316
rect 15427 6276 16212 6304
rect 15427 6273 15439 6276
rect 15381 6267 15439 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 18141 6307 18199 6313
rect 18141 6273 18153 6307
rect 18187 6304 18199 6307
rect 18708 6304 18736 6400
rect 18187 6276 18736 6304
rect 18187 6273 18199 6276
rect 18141 6267 18199 6273
rect 18782 6264 18788 6316
rect 18840 6304 18846 6316
rect 18840 6276 18885 6304
rect 18840 6264 18846 6276
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6205 14427 6239
rect 14369 6199 14427 6205
rect 14737 6239 14795 6245
rect 14737 6205 14749 6239
rect 14783 6205 14795 6239
rect 15102 6236 15108 6248
rect 15063 6208 15108 6236
rect 14737 6199 14795 6205
rect 11072 6140 11652 6168
rect 11624 6112 11652 6140
rect 1762 6060 1768 6112
rect 1820 6100 1826 6112
rect 2406 6100 2412 6112
rect 1820 6072 2412 6100
rect 1820 6060 1826 6072
rect 2406 6060 2412 6072
rect 2464 6100 2470 6112
rect 2639 6103 2697 6109
rect 2639 6100 2651 6103
rect 2464 6072 2651 6100
rect 2464 6060 2470 6072
rect 2639 6069 2651 6072
rect 2685 6069 2697 6103
rect 2639 6063 2697 6069
rect 5077 6103 5135 6109
rect 5077 6069 5089 6103
rect 5123 6100 5135 6103
rect 5258 6100 5264 6112
rect 5123 6072 5264 6100
rect 5123 6069 5135 6072
rect 5077 6063 5135 6069
rect 5258 6060 5264 6072
rect 5316 6100 5322 6112
rect 5810 6100 5816 6112
rect 5316 6072 5816 6100
rect 5316 6060 5322 6072
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 5994 6060 6000 6112
rect 6052 6100 6058 6112
rect 6273 6103 6331 6109
rect 6273 6100 6285 6103
rect 6052 6072 6285 6100
rect 6052 6060 6058 6072
rect 6273 6069 6285 6072
rect 6319 6100 6331 6103
rect 6362 6100 6368 6112
rect 6319 6072 6368 6100
rect 6319 6069 6331 6072
rect 6273 6063 6331 6069
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6546 6100 6552 6112
rect 6507 6072 6552 6100
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 7834 6100 7840 6112
rect 7795 6072 7840 6100
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 7926 6060 7932 6112
rect 7984 6100 7990 6112
rect 8297 6103 8355 6109
rect 8297 6100 8309 6103
rect 7984 6072 8309 6100
rect 7984 6060 7990 6072
rect 8297 6069 8309 6072
rect 8343 6100 8355 6103
rect 9306 6100 9312 6112
rect 8343 6072 9312 6100
rect 8343 6069 8355 6072
rect 8297 6063 8355 6069
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 9861 6103 9919 6109
rect 9861 6100 9873 6103
rect 9824 6072 9873 6100
rect 9824 6060 9830 6072
rect 9861 6069 9873 6072
rect 9907 6069 9919 6103
rect 9861 6063 9919 6069
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 11238 6100 11244 6112
rect 10100 6072 11244 6100
rect 10100 6060 10106 6072
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 11606 6060 11612 6112
rect 11664 6100 11670 6112
rect 11977 6103 12035 6109
rect 11977 6100 11989 6103
rect 11664 6072 11989 6100
rect 11664 6060 11670 6072
rect 11977 6069 11989 6072
rect 12023 6100 12035 6103
rect 12894 6100 12900 6112
rect 12023 6072 12900 6100
rect 12023 6069 12035 6072
rect 11977 6063 12035 6069
rect 12894 6060 12900 6072
rect 12952 6100 12958 6112
rect 13725 6103 13783 6109
rect 13725 6100 13737 6103
rect 12952 6072 13737 6100
rect 12952 6060 12958 6072
rect 13725 6069 13737 6072
rect 13771 6100 13783 6103
rect 14752 6100 14780 6199
rect 15102 6196 15108 6208
rect 15160 6196 15166 6248
rect 19702 6245 19708 6248
rect 19680 6239 19708 6245
rect 19680 6236 19692 6239
rect 19615 6208 19692 6236
rect 19680 6205 19692 6208
rect 19760 6236 19766 6248
rect 20073 6239 20131 6245
rect 20073 6236 20085 6239
rect 19760 6208 20085 6236
rect 19680 6199 19708 6205
rect 19702 6196 19708 6199
rect 19760 6196 19766 6208
rect 20073 6205 20085 6208
rect 20119 6205 20131 6239
rect 20073 6199 20131 6205
rect 16114 6128 16120 6180
rect 16172 6168 16178 6180
rect 16530 6171 16588 6177
rect 16530 6168 16542 6171
rect 16172 6140 16542 6168
rect 16172 6128 16178 6140
rect 16530 6137 16542 6140
rect 16576 6137 16588 6171
rect 16530 6131 16588 6137
rect 17770 6128 17776 6180
rect 17828 6168 17834 6180
rect 18233 6171 18291 6177
rect 18233 6168 18245 6171
rect 17828 6140 18245 6168
rect 17828 6128 17834 6140
rect 18233 6137 18245 6140
rect 18279 6137 18291 6171
rect 18233 6131 18291 6137
rect 15657 6103 15715 6109
rect 15657 6100 15669 6103
rect 13771 6072 15669 6100
rect 13771 6069 13783 6072
rect 13725 6063 13783 6069
rect 15657 6069 15669 6072
rect 15703 6100 15715 6103
rect 15930 6100 15936 6112
rect 15703 6072 15936 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 19058 6100 19064 6112
rect 16264 6072 19064 6100
rect 16264 6060 16270 6072
rect 19058 6060 19064 6072
rect 19116 6100 19122 6112
rect 19153 6103 19211 6109
rect 19153 6100 19165 6103
rect 19116 6072 19165 6100
rect 19116 6060 19122 6072
rect 19153 6069 19165 6072
rect 19199 6069 19211 6103
rect 19153 6063 19211 6069
rect 1104 6010 20884 6032
rect 1104 5958 8315 6010
rect 8367 5958 8379 6010
rect 8431 5958 8443 6010
rect 8495 5958 8507 6010
rect 8559 5958 15648 6010
rect 15700 5958 15712 6010
rect 15764 5958 15776 6010
rect 15828 5958 15840 6010
rect 15892 5958 20884 6010
rect 1104 5936 20884 5958
rect 6822 5896 6828 5908
rect 6783 5868 6828 5896
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 8846 5896 8852 5908
rect 8220 5868 8852 5896
rect 2958 5788 2964 5840
rect 3016 5828 3022 5840
rect 7006 5828 7012 5840
rect 3016 5800 7012 5828
rect 3016 5788 3022 5800
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 2130 5760 2136 5772
rect 1912 5732 2136 5760
rect 1912 5720 1918 5732
rect 2130 5720 2136 5732
rect 2188 5760 2194 5772
rect 2225 5763 2283 5769
rect 2225 5760 2237 5763
rect 2188 5732 2237 5760
rect 2188 5720 2194 5732
rect 2225 5729 2237 5732
rect 2271 5729 2283 5763
rect 2225 5723 2283 5729
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 4982 5760 4988 5772
rect 4111 5732 4988 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 3326 5652 3332 5704
rect 3384 5692 3390 5704
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3384 5664 3801 5692
rect 3384 5652 3390 5664
rect 3789 5661 3801 5664
rect 3835 5692 3847 5695
rect 4080 5692 4108 5723
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 6472 5769 6500 5800
rect 7006 5788 7012 5800
rect 7064 5788 7070 5840
rect 8110 5828 8116 5840
rect 8071 5800 8116 5828
rect 8110 5788 8116 5800
rect 8168 5788 8174 5840
rect 8220 5837 8248 5868
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 9122 5896 9128 5908
rect 9035 5868 9128 5896
rect 9122 5856 9128 5868
rect 9180 5896 9186 5908
rect 10686 5896 10692 5908
rect 9180 5868 10692 5896
rect 9180 5856 9186 5868
rect 10686 5856 10692 5868
rect 10744 5896 10750 5908
rect 11698 5896 11704 5908
rect 10744 5868 11560 5896
rect 11659 5868 11704 5896
rect 10744 5856 10750 5868
rect 8205 5831 8263 5837
rect 8205 5797 8217 5831
rect 8251 5797 8263 5831
rect 8205 5791 8263 5797
rect 8754 5788 8760 5840
rect 8812 5828 8818 5840
rect 9398 5828 9404 5840
rect 8812 5800 9404 5828
rect 8812 5788 8818 5800
rect 9398 5788 9404 5800
rect 9456 5828 9462 5840
rect 10229 5831 10287 5837
rect 10229 5828 10241 5831
rect 9456 5800 10241 5828
rect 9456 5788 9462 5800
rect 10229 5797 10241 5800
rect 10275 5828 10287 5831
rect 10870 5828 10876 5840
rect 10275 5800 10876 5828
rect 10275 5797 10287 5800
rect 10229 5791 10287 5797
rect 10870 5788 10876 5800
rect 10928 5788 10934 5840
rect 11532 5837 11560 5868
rect 11698 5856 11704 5868
rect 11756 5856 11762 5908
rect 12526 5896 12532 5908
rect 11808 5868 12532 5896
rect 11808 5840 11836 5868
rect 12526 5856 12532 5868
rect 12584 5896 12590 5908
rect 14642 5896 14648 5908
rect 12584 5868 14648 5896
rect 12584 5856 12590 5868
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 14737 5899 14795 5905
rect 14737 5865 14749 5899
rect 14783 5896 14795 5899
rect 15102 5896 15108 5908
rect 14783 5868 15108 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15470 5896 15476 5908
rect 15431 5868 15476 5896
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 16577 5899 16635 5905
rect 16577 5865 16589 5899
rect 16623 5896 16635 5899
rect 17402 5896 17408 5908
rect 16623 5868 17408 5896
rect 16623 5865 16635 5868
rect 16577 5859 16635 5865
rect 17402 5856 17408 5868
rect 17460 5896 17466 5908
rect 17460 5868 17632 5896
rect 17460 5856 17466 5868
rect 11517 5831 11575 5837
rect 11517 5797 11529 5831
rect 11563 5828 11575 5831
rect 11790 5828 11796 5840
rect 11563 5800 11796 5828
rect 11563 5797 11575 5800
rect 11517 5791 11575 5797
rect 11790 5788 11796 5800
rect 11848 5788 11854 5840
rect 12342 5828 12348 5840
rect 11900 5800 12348 5828
rect 11900 5772 11928 5800
rect 12342 5788 12348 5800
rect 12400 5828 12406 5840
rect 13541 5831 13599 5837
rect 13541 5828 13553 5831
rect 12400 5800 13553 5828
rect 12400 5788 12406 5800
rect 13541 5797 13553 5800
rect 13587 5828 13599 5831
rect 13725 5831 13783 5837
rect 13725 5828 13737 5831
rect 13587 5800 13737 5828
rect 13587 5797 13599 5800
rect 13541 5791 13599 5797
rect 13725 5797 13737 5800
rect 13771 5797 13783 5831
rect 13998 5828 14004 5840
rect 13959 5800 14004 5828
rect 13725 5791 13783 5797
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 16019 5831 16077 5837
rect 16019 5797 16031 5831
rect 16065 5828 16077 5831
rect 16114 5828 16120 5840
rect 16065 5800 16120 5828
rect 16065 5797 16077 5800
rect 16019 5791 16077 5797
rect 16114 5788 16120 5800
rect 16172 5828 16178 5840
rect 17604 5837 17632 5868
rect 18138 5856 18144 5908
rect 18196 5896 18202 5908
rect 18417 5899 18475 5905
rect 18417 5896 18429 5899
rect 18196 5868 18429 5896
rect 18196 5856 18202 5868
rect 18417 5865 18429 5868
rect 18463 5865 18475 5899
rect 18782 5896 18788 5908
rect 18743 5868 18788 5896
rect 18417 5859 18475 5865
rect 18782 5856 18788 5868
rect 18840 5856 18846 5908
rect 16853 5831 16911 5837
rect 16853 5828 16865 5831
rect 16172 5800 16865 5828
rect 16172 5788 16178 5800
rect 16853 5797 16865 5800
rect 16899 5797 16911 5831
rect 16853 5791 16911 5797
rect 17589 5831 17647 5837
rect 17589 5797 17601 5831
rect 17635 5797 17647 5831
rect 17589 5791 17647 5797
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5729 5687 5763
rect 5629 5723 5687 5729
rect 6365 5763 6423 5769
rect 6365 5729 6377 5763
rect 6411 5729 6423 5763
rect 6365 5723 6423 5729
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5729 6515 5763
rect 6457 5723 6515 5729
rect 6917 5763 6975 5769
rect 6917 5729 6929 5763
rect 6963 5760 6975 5763
rect 7834 5760 7840 5772
rect 6963 5732 7840 5760
rect 6963 5729 6975 5732
rect 6917 5723 6975 5729
rect 3835 5664 4108 5692
rect 4433 5695 4491 5701
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 4433 5661 4445 5695
rect 4479 5692 4491 5695
rect 4522 5692 4528 5704
rect 4479 5664 4528 5692
rect 4479 5661 4491 5664
rect 4433 5655 4491 5661
rect 4522 5652 4528 5664
rect 4580 5692 4586 5704
rect 5644 5692 5672 5723
rect 4580 5664 5672 5692
rect 6380 5692 6408 5723
rect 6638 5692 6644 5704
rect 6380 5664 6644 5692
rect 4580 5652 4586 5664
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 4062 5584 4068 5636
rect 4120 5624 4126 5636
rect 5169 5627 5227 5633
rect 5169 5624 5181 5627
rect 4120 5596 5181 5624
rect 4120 5584 4126 5596
rect 5169 5593 5181 5596
rect 5215 5624 5227 5627
rect 5350 5624 5356 5636
rect 5215 5596 5356 5624
rect 5215 5593 5227 5596
rect 5169 5587 5227 5593
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 5994 5584 6000 5636
rect 6052 5624 6058 5636
rect 6932 5624 6960 5723
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 11882 5760 11888 5772
rect 11843 5732 11888 5760
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 12069 5763 12127 5769
rect 12069 5760 12081 5763
rect 12032 5732 12081 5760
rect 12032 5720 12038 5732
rect 12069 5729 12081 5732
rect 12115 5729 12127 5763
rect 12526 5760 12532 5772
rect 12487 5732 12532 5760
rect 12069 5723 12127 5729
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 12802 5760 12808 5772
rect 12763 5732 12808 5760
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 13170 5720 13176 5772
rect 13228 5760 13234 5772
rect 14093 5763 14151 5769
rect 14093 5760 14105 5763
rect 13228 5732 14105 5760
rect 13228 5720 13234 5732
rect 14093 5729 14105 5732
rect 14139 5729 14151 5763
rect 14093 5723 14151 5729
rect 18141 5763 18199 5769
rect 18141 5729 18153 5763
rect 18187 5760 18199 5763
rect 18874 5760 18880 5772
rect 18187 5732 18880 5760
rect 18187 5729 18199 5732
rect 18141 5723 18199 5729
rect 18874 5720 18880 5732
rect 18932 5720 18938 5772
rect 19058 5760 19064 5772
rect 19019 5732 19064 5760
rect 19058 5720 19064 5732
rect 19116 5720 19122 5772
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5692 10195 5695
rect 10502 5692 10508 5704
rect 10183 5664 10508 5692
rect 10183 5661 10195 5664
rect 10137 5655 10195 5661
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5692 10839 5695
rect 12618 5692 12624 5704
rect 10827 5664 12624 5692
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 6052 5596 6960 5624
rect 6052 5584 6058 5596
rect 7190 5584 7196 5636
rect 7248 5624 7254 5636
rect 7745 5627 7803 5633
rect 7745 5624 7757 5627
rect 7248 5596 7757 5624
rect 7248 5584 7254 5596
rect 7745 5593 7757 5596
rect 7791 5593 7803 5627
rect 7745 5587 7803 5593
rect 8665 5627 8723 5633
rect 8665 5593 8677 5627
rect 8711 5624 8723 5627
rect 10796 5624 10824 5655
rect 12618 5652 12624 5664
rect 12676 5652 12682 5704
rect 13722 5692 13728 5704
rect 13635 5664 13728 5692
rect 13722 5652 13728 5664
rect 13780 5692 13786 5704
rect 15470 5692 15476 5704
rect 13780 5664 15476 5692
rect 13780 5652 13786 5664
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 15654 5692 15660 5704
rect 15615 5664 15660 5692
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 17313 5695 17371 5701
rect 17313 5661 17325 5695
rect 17359 5692 17371 5695
rect 17497 5695 17555 5701
rect 17497 5692 17509 5695
rect 17359 5664 17509 5692
rect 17359 5661 17371 5664
rect 17313 5655 17371 5661
rect 17497 5661 17509 5664
rect 17543 5692 17555 5695
rect 18414 5692 18420 5704
rect 17543 5664 18420 5692
rect 17543 5661 17555 5664
rect 17497 5655 17555 5661
rect 18414 5652 18420 5664
rect 18472 5652 18478 5704
rect 18506 5652 18512 5704
rect 18564 5692 18570 5704
rect 18969 5695 19027 5701
rect 18969 5692 18981 5695
rect 18564 5664 18981 5692
rect 18564 5652 18570 5664
rect 18969 5661 18981 5664
rect 19015 5661 19027 5695
rect 18969 5655 19027 5661
rect 8711 5596 10824 5624
rect 14277 5627 14335 5633
rect 8711 5593 8723 5596
rect 8665 5587 8723 5593
rect 14277 5593 14289 5627
rect 14323 5624 14335 5627
rect 15930 5624 15936 5636
rect 14323 5596 15936 5624
rect 14323 5593 14335 5596
rect 14277 5587 14335 5593
rect 15930 5584 15936 5596
rect 15988 5584 15994 5636
rect 1765 5559 1823 5565
rect 1765 5525 1777 5559
rect 1811 5556 1823 5559
rect 1854 5556 1860 5568
rect 1811 5528 1860 5556
rect 1811 5525 1823 5528
rect 1765 5519 1823 5525
rect 1854 5516 1860 5528
rect 1912 5516 1918 5568
rect 2406 5556 2412 5568
rect 2367 5528 2412 5556
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 3510 5556 3516 5568
rect 3471 5528 3516 5556
rect 3510 5516 3516 5528
rect 3568 5516 3574 5568
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 4203 5559 4261 5565
rect 4203 5556 4215 5559
rect 3936 5528 4215 5556
rect 3936 5516 3942 5528
rect 4203 5525 4215 5528
rect 4249 5525 4261 5559
rect 4203 5519 4261 5525
rect 4341 5559 4399 5565
rect 4341 5525 4353 5559
rect 4387 5556 4399 5559
rect 4430 5556 4436 5568
rect 4387 5528 4436 5556
rect 4387 5525 4399 5528
rect 4341 5519 4399 5525
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 4709 5559 4767 5565
rect 4709 5525 4721 5559
rect 4755 5556 4767 5559
rect 7282 5556 7288 5568
rect 4755 5528 7288 5556
rect 4755 5525 4767 5528
rect 4709 5519 4767 5525
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 7466 5556 7472 5568
rect 7427 5528 7472 5556
rect 7466 5516 7472 5528
rect 7524 5516 7530 5568
rect 9398 5556 9404 5568
rect 9359 5528 9404 5556
rect 9398 5516 9404 5528
rect 9456 5556 9462 5568
rect 9861 5559 9919 5565
rect 9861 5556 9873 5559
rect 9456 5528 9873 5556
rect 9456 5516 9462 5528
rect 9861 5525 9873 5528
rect 9907 5556 9919 5559
rect 10410 5556 10416 5568
rect 9907 5528 10416 5556
rect 9907 5525 9919 5528
rect 9861 5519 9919 5525
rect 10410 5516 10416 5528
rect 10468 5556 10474 5568
rect 10962 5556 10968 5568
rect 10468 5528 10968 5556
rect 10468 5516 10474 5528
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 11054 5516 11060 5568
rect 11112 5556 11118 5568
rect 11149 5559 11207 5565
rect 11149 5556 11161 5559
rect 11112 5528 11161 5556
rect 11112 5516 11118 5528
rect 11149 5525 11161 5528
rect 11195 5556 11207 5559
rect 12802 5556 12808 5568
rect 11195 5528 12808 5556
rect 11195 5525 11207 5528
rect 11149 5519 11207 5525
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 1104 5466 20884 5488
rect 1104 5414 4648 5466
rect 4700 5414 4712 5466
rect 4764 5414 4776 5466
rect 4828 5414 4840 5466
rect 4892 5414 11982 5466
rect 12034 5414 12046 5466
rect 12098 5414 12110 5466
rect 12162 5414 12174 5466
rect 12226 5414 19315 5466
rect 19367 5414 19379 5466
rect 19431 5414 19443 5466
rect 19495 5414 19507 5466
rect 19559 5414 20884 5466
rect 1104 5392 20884 5414
rect 2222 5312 2228 5364
rect 2280 5352 2286 5364
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 2280 5324 2605 5352
rect 2280 5312 2286 5324
rect 2593 5321 2605 5324
rect 2639 5352 2651 5355
rect 4246 5352 4252 5364
rect 2639 5324 4252 5352
rect 2639 5321 2651 5324
rect 2593 5315 2651 5321
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 4338 5312 4344 5364
rect 4396 5352 4402 5364
rect 5261 5355 5319 5361
rect 5261 5352 5273 5355
rect 4396 5324 5273 5352
rect 4396 5312 4402 5324
rect 5261 5321 5273 5324
rect 5307 5352 5319 5355
rect 6914 5352 6920 5364
rect 5307 5324 6920 5352
rect 5307 5321 5319 5324
rect 5261 5315 5319 5321
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 7929 5355 7987 5361
rect 7929 5321 7941 5355
rect 7975 5352 7987 5355
rect 8754 5352 8760 5364
rect 7975 5324 8760 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 10778 5312 10784 5364
rect 10836 5352 10842 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 10836 5324 10885 5352
rect 10836 5312 10842 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 4522 5244 4528 5296
rect 4580 5284 4586 5296
rect 4801 5287 4859 5293
rect 4801 5284 4813 5287
rect 4580 5256 4813 5284
rect 4580 5244 4586 5256
rect 4801 5253 4813 5256
rect 4847 5253 4859 5287
rect 4801 5247 4859 5253
rect 5150 5287 5208 5293
rect 5150 5253 5162 5287
rect 5196 5284 5208 5287
rect 5534 5284 5540 5296
rect 5196 5256 5540 5284
rect 5196 5253 5208 5256
rect 5150 5247 5208 5253
rect 4816 5216 4844 5247
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 5810 5244 5816 5296
rect 5868 5284 5874 5296
rect 7466 5284 7472 5296
rect 5868 5256 7472 5284
rect 5868 5244 5874 5256
rect 7466 5244 7472 5256
rect 7524 5244 7530 5296
rect 7834 5244 7840 5296
rect 7892 5284 7898 5296
rect 8573 5287 8631 5293
rect 8573 5284 8585 5287
rect 7892 5256 8585 5284
rect 7892 5244 7898 5256
rect 8573 5253 8585 5256
rect 8619 5253 8631 5287
rect 8573 5247 8631 5253
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 4816 5188 5365 5216
rect 5353 5185 5365 5188
rect 5399 5216 5411 5219
rect 5626 5216 5632 5228
rect 5399 5188 5632 5216
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 5721 5219 5779 5225
rect 5721 5185 5733 5219
rect 5767 5216 5779 5219
rect 6178 5216 6184 5228
rect 5767 5188 6184 5216
rect 5767 5185 5779 5188
rect 5721 5179 5779 5185
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 8588 5216 8616 5247
rect 8662 5244 8668 5296
rect 8720 5284 8726 5296
rect 9122 5284 9128 5296
rect 8720 5256 9128 5284
rect 8720 5244 8726 5256
rect 9122 5244 9128 5256
rect 9180 5244 9186 5296
rect 8754 5216 8760 5228
rect 8588 5188 8760 5216
rect 8754 5176 8760 5188
rect 8812 5216 8818 5228
rect 8812 5188 9628 5216
rect 8812 5176 8818 5188
rect 1578 5148 1584 5160
rect 1539 5120 1584 5148
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 3421 5151 3479 5157
rect 3421 5117 3433 5151
rect 3467 5117 3479 5151
rect 3421 5111 3479 5117
rect 2133 5083 2191 5089
rect 2133 5049 2145 5083
rect 2179 5080 2191 5083
rect 3326 5080 3332 5092
rect 2179 5052 3332 5080
rect 2179 5049 2191 5052
rect 2133 5043 2191 5049
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 3436 5080 3464 5111
rect 3510 5108 3516 5160
rect 3568 5148 3574 5160
rect 7009 5151 7067 5157
rect 7009 5148 7021 5151
rect 3568 5120 7021 5148
rect 3568 5108 3574 5120
rect 7009 5117 7021 5120
rect 7055 5148 7067 5151
rect 7834 5148 7840 5160
rect 7055 5120 7840 5148
rect 7055 5117 7067 5120
rect 7009 5111 7067 5117
rect 7834 5108 7840 5120
rect 7892 5108 7898 5160
rect 8018 5108 8024 5160
rect 8076 5148 8082 5160
rect 8202 5148 8208 5160
rect 8076 5120 8208 5148
rect 8076 5108 8082 5120
rect 8202 5108 8208 5120
rect 8260 5148 8266 5160
rect 9030 5148 9036 5160
rect 8260 5120 8892 5148
rect 8991 5120 9036 5148
rect 8260 5108 8266 5120
rect 3602 5080 3608 5092
rect 3436 5052 3608 5080
rect 3602 5040 3608 5052
rect 3660 5040 3666 5092
rect 3694 5040 3700 5092
rect 3752 5080 3758 5092
rect 4982 5080 4988 5092
rect 3752 5052 4819 5080
rect 4895 5052 4988 5080
rect 3752 5040 3758 5052
rect 2958 5012 2964 5024
rect 2919 4984 2964 5012
rect 2958 4972 2964 4984
rect 3016 4972 3022 5024
rect 3510 5012 3516 5024
rect 3471 4984 3516 5012
rect 3510 4972 3516 4984
rect 3568 4972 3574 5024
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 4065 5015 4123 5021
rect 4065 5012 4077 5015
rect 3936 4984 4077 5012
rect 3936 4972 3942 4984
rect 4065 4981 4077 4984
rect 4111 4981 4123 5015
rect 4430 5012 4436 5024
rect 4391 4984 4436 5012
rect 4065 4975 4123 4981
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 4791 5012 4819 5052
rect 4982 5040 4988 5052
rect 5040 5080 5046 5092
rect 7098 5080 7104 5092
rect 5040 5052 7104 5080
rect 5040 5040 5046 5052
rect 7098 5040 7104 5052
rect 7156 5040 7162 5092
rect 7190 5040 7196 5092
rect 7248 5080 7254 5092
rect 7330 5083 7388 5089
rect 7330 5080 7342 5083
rect 7248 5052 7342 5080
rect 7248 5040 7254 5052
rect 7330 5049 7342 5052
rect 7376 5049 7388 5083
rect 8864 5080 8892 5120
rect 9030 5108 9036 5120
rect 9088 5108 9094 5160
rect 9217 5151 9275 5157
rect 9217 5117 9229 5151
rect 9263 5148 9275 5151
rect 9398 5148 9404 5160
rect 9263 5120 9404 5148
rect 9263 5117 9275 5120
rect 9217 5111 9275 5117
rect 9232 5080 9260 5111
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 9600 5157 9628 5188
rect 9585 5151 9643 5157
rect 9585 5117 9597 5151
rect 9631 5148 9643 5151
rect 9766 5148 9772 5160
rect 9631 5120 9772 5148
rect 9631 5117 9643 5120
rect 9585 5111 9643 5117
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 10134 5148 10140 5160
rect 10047 5120 10140 5148
rect 10134 5108 10140 5120
rect 10192 5148 10198 5160
rect 10689 5151 10747 5157
rect 10689 5148 10701 5151
rect 10192 5120 10701 5148
rect 10192 5108 10198 5120
rect 10689 5117 10701 5120
rect 10735 5117 10747 5151
rect 10888 5148 10916 5315
rect 10962 5312 10968 5364
rect 11020 5352 11026 5364
rect 11609 5355 11667 5361
rect 11609 5352 11621 5355
rect 11020 5324 11621 5352
rect 11020 5312 11026 5324
rect 11609 5321 11621 5324
rect 11655 5321 11667 5355
rect 11609 5315 11667 5321
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12986 5352 12992 5364
rect 12299 5324 12992 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 11624 5284 11652 5315
rect 11882 5284 11888 5296
rect 11624 5256 11888 5284
rect 11882 5244 11888 5256
rect 11940 5244 11946 5296
rect 12452 5157 12480 5324
rect 12986 5312 12992 5324
rect 13044 5312 13050 5364
rect 17402 5352 17408 5364
rect 17363 5324 17408 5352
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 18414 5312 18420 5364
rect 18472 5352 18478 5364
rect 19058 5352 19064 5364
rect 18472 5324 19064 5352
rect 18472 5312 18478 5324
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 12710 5244 12716 5296
rect 12768 5284 12774 5296
rect 13541 5287 13599 5293
rect 13541 5284 13553 5287
rect 12768 5256 13553 5284
rect 12768 5244 12774 5256
rect 13541 5253 13553 5256
rect 13587 5253 13599 5287
rect 13541 5247 13599 5253
rect 18693 5287 18751 5293
rect 18693 5253 18705 5287
rect 18739 5284 18751 5287
rect 18874 5284 18880 5296
rect 18739 5256 18880 5284
rect 18739 5253 18751 5256
rect 18693 5247 18751 5253
rect 13556 5216 13584 5247
rect 18874 5244 18880 5256
rect 18932 5244 18938 5296
rect 15197 5219 15255 5225
rect 13556 5188 14228 5216
rect 11057 5151 11115 5157
rect 11057 5148 11069 5151
rect 10888 5120 11069 5148
rect 10689 5111 10747 5117
rect 11057 5117 11069 5120
rect 11103 5117 11115 5151
rect 11057 5111 11115 5117
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5117 12495 5151
rect 13722 5148 13728 5160
rect 13683 5120 13728 5148
rect 12437 5111 12495 5117
rect 13722 5108 13728 5120
rect 13780 5108 13786 5160
rect 14200 5157 14228 5188
rect 15197 5185 15209 5219
rect 15243 5216 15255 5219
rect 15654 5216 15660 5228
rect 15243 5188 15660 5216
rect 15243 5185 15255 5188
rect 15197 5179 15255 5185
rect 15654 5176 15660 5188
rect 15712 5216 15718 5228
rect 16758 5216 16764 5228
rect 15712 5188 16764 5216
rect 15712 5176 15718 5188
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 18141 5219 18199 5225
rect 18141 5185 18153 5219
rect 18187 5216 18199 5219
rect 18782 5216 18788 5228
rect 18187 5188 18788 5216
rect 18187 5185 18199 5188
rect 18141 5179 18199 5185
rect 18782 5176 18788 5188
rect 18840 5176 18846 5228
rect 14185 5151 14243 5157
rect 14185 5117 14197 5151
rect 14231 5117 14243 5151
rect 14642 5148 14648 5160
rect 14603 5120 14648 5148
rect 14185 5111 14243 5117
rect 14642 5108 14648 5120
rect 14700 5108 14706 5160
rect 15102 5148 15108 5160
rect 15063 5120 15108 5148
rect 15102 5108 15108 5120
rect 15160 5108 15166 5160
rect 16022 5148 16028 5160
rect 15983 5120 16028 5148
rect 16022 5108 16028 5120
rect 16080 5108 16086 5160
rect 16945 5151 17003 5157
rect 16945 5117 16957 5151
rect 16991 5148 17003 5151
rect 17773 5151 17831 5157
rect 17773 5148 17785 5151
rect 16991 5120 17785 5148
rect 16991 5117 17003 5120
rect 16945 5111 17003 5117
rect 17773 5117 17785 5120
rect 17819 5117 17831 5151
rect 17773 5111 17831 5117
rect 13170 5080 13176 5092
rect 8864 5052 9260 5080
rect 10381 5052 13176 5080
rect 7330 5043 7388 5049
rect 5994 5012 6000 5024
rect 4791 4984 6000 5012
rect 5994 4972 6000 4984
rect 6052 4972 6058 5024
rect 6457 5015 6515 5021
rect 6457 4981 6469 5015
rect 6503 5012 6515 5015
rect 6638 5012 6644 5024
rect 6503 4984 6644 5012
rect 6503 4981 6515 4984
rect 6457 4975 6515 4981
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 9030 5012 9036 5024
rect 8991 4984 9036 5012
rect 9030 4972 9036 4984
rect 9088 4972 9094 5024
rect 9582 4972 9588 5024
rect 9640 5012 9646 5024
rect 10381 5012 10409 5052
rect 13170 5040 13176 5052
rect 13228 5040 13234 5092
rect 16346 5083 16404 5089
rect 16346 5049 16358 5083
rect 16392 5049 16404 5083
rect 16346 5043 16404 5049
rect 9640 4984 10409 5012
rect 10597 5015 10655 5021
rect 9640 4972 9646 4984
rect 10597 4981 10609 5015
rect 10643 5012 10655 5015
rect 10689 5015 10747 5021
rect 10689 5012 10701 5015
rect 10643 4984 10701 5012
rect 10643 4981 10655 4984
rect 10597 4975 10655 4981
rect 10689 4981 10701 4984
rect 10735 5012 10747 5015
rect 10962 5012 10968 5024
rect 10735 4984 10968 5012
rect 10735 4981 10747 4984
rect 10689 4975 10747 4981
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 11241 5015 11299 5021
rect 11241 5012 11253 5015
rect 11112 4984 11253 5012
rect 11112 4972 11118 4984
rect 11241 4981 11253 4984
rect 11287 4981 11299 5015
rect 11241 4975 11299 4981
rect 12621 5015 12679 5021
rect 12621 4981 12633 5015
rect 12667 5012 12679 5015
rect 12894 5012 12900 5024
rect 12667 4984 12900 5012
rect 12667 4981 12679 4984
rect 12621 4975 12679 4981
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 15473 5015 15531 5021
rect 15473 5012 15485 5015
rect 15436 4984 15485 5012
rect 15436 4972 15442 4984
rect 15473 4981 15485 4984
rect 15519 5012 15531 5015
rect 15841 5015 15899 5021
rect 15841 5012 15853 5015
rect 15519 4984 15853 5012
rect 15519 4981 15531 4984
rect 15473 4975 15531 4981
rect 15841 4981 15853 4984
rect 15887 5012 15899 5015
rect 16114 5012 16120 5024
rect 15887 4984 16120 5012
rect 15887 4981 15899 4984
rect 15841 4975 15899 4981
rect 16114 4972 16120 4984
rect 16172 5012 16178 5024
rect 16361 5012 16389 5043
rect 16172 4984 16389 5012
rect 17788 5012 17816 5111
rect 18233 5083 18291 5089
rect 18233 5049 18245 5083
rect 18279 5049 18291 5083
rect 18233 5043 18291 5049
rect 18248 5012 18276 5043
rect 17788 4984 18276 5012
rect 16172 4972 16178 4984
rect 19150 4972 19156 5024
rect 19208 5012 19214 5024
rect 19613 5015 19671 5021
rect 19613 5012 19625 5015
rect 19208 4984 19625 5012
rect 19208 4972 19214 4984
rect 19613 4981 19625 4984
rect 19659 4981 19671 5015
rect 19613 4975 19671 4981
rect 1104 4922 20884 4944
rect 1104 4870 8315 4922
rect 8367 4870 8379 4922
rect 8431 4870 8443 4922
rect 8495 4870 8507 4922
rect 8559 4870 15648 4922
rect 15700 4870 15712 4922
rect 15764 4870 15776 4922
rect 15828 4870 15840 4922
rect 15892 4870 20884 4922
rect 1104 4848 20884 4870
rect 842 4768 848 4820
rect 900 4808 906 4820
rect 1578 4808 1584 4820
rect 900 4780 1584 4808
rect 900 4768 906 4780
rect 1578 4768 1584 4780
rect 1636 4768 1642 4820
rect 2222 4808 2228 4820
rect 2183 4780 2228 4808
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 3326 4768 3332 4820
rect 3384 4808 3390 4820
rect 3421 4811 3479 4817
rect 3421 4808 3433 4811
rect 3384 4780 3433 4808
rect 3384 4768 3390 4780
rect 3421 4777 3433 4780
rect 3467 4777 3479 4811
rect 3421 4771 3479 4777
rect 4341 4811 4399 4817
rect 4341 4777 4353 4811
rect 4387 4808 4399 4811
rect 4522 4808 4528 4820
rect 4387 4780 4528 4808
rect 4387 4777 4399 4780
rect 4341 4771 4399 4777
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 5626 4808 5632 4820
rect 5587 4780 5632 4808
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 6454 4808 6460 4820
rect 6415 4780 6460 4808
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 7282 4768 7288 4820
rect 7340 4808 7346 4820
rect 8297 4811 8355 4817
rect 8297 4808 8309 4811
rect 7340 4780 8309 4808
rect 7340 4768 7346 4780
rect 8297 4777 8309 4780
rect 8343 4808 8355 4811
rect 9122 4808 9128 4820
rect 8343 4780 9128 4808
rect 8343 4777 8355 4780
rect 8297 4771 8355 4777
rect 9122 4768 9128 4780
rect 9180 4808 9186 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9180 4780 9413 4808
rect 9180 4768 9186 4780
rect 9401 4777 9413 4780
rect 9447 4808 9459 4811
rect 10134 4808 10140 4820
rect 9447 4780 10140 4808
rect 9447 4777 9459 4780
rect 9401 4771 9459 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 10870 4808 10876 4820
rect 10831 4780 10876 4808
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 12069 4811 12127 4817
rect 12069 4777 12081 4811
rect 12115 4808 12127 4811
rect 12115 4780 15148 4808
rect 12115 4777 12127 4780
rect 12069 4771 12127 4777
rect 2406 4700 2412 4752
rect 2464 4740 2470 4752
rect 2501 4743 2559 4749
rect 2501 4740 2513 4743
rect 2464 4712 2513 4740
rect 2464 4700 2470 4712
rect 2501 4709 2513 4712
rect 2547 4709 2559 4743
rect 3050 4740 3056 4752
rect 3011 4712 3056 4740
rect 2501 4703 2559 4709
rect 3050 4700 3056 4712
rect 3108 4700 3114 4752
rect 4246 4700 4252 4752
rect 4304 4740 4310 4752
rect 4801 4743 4859 4749
rect 4801 4740 4813 4743
rect 4304 4712 4813 4740
rect 4304 4700 4310 4712
rect 4801 4709 4813 4712
rect 4847 4740 4859 4743
rect 4847 4712 5580 4740
rect 4847 4709 4859 4712
rect 4801 4703 4859 4709
rect 5350 4632 5356 4684
rect 5408 4672 5414 4684
rect 5408 4644 5453 4672
rect 5408 4632 5414 4644
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2682 4604 2688 4616
rect 2455 4576 2688 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4212 4576 4721 4604
rect 4212 4564 4218 4576
rect 4709 4573 4721 4576
rect 4755 4573 4767 4607
rect 5552 4604 5580 4712
rect 5644 4672 5672 4768
rect 6089 4743 6147 4749
rect 6089 4709 6101 4743
rect 6135 4740 6147 4743
rect 6914 4740 6920 4752
rect 6135 4712 6920 4740
rect 6135 4709 6147 4712
rect 6089 4703 6147 4709
rect 6914 4700 6920 4712
rect 6972 4700 6978 4752
rect 7745 4743 7803 4749
rect 7745 4709 7757 4743
rect 7791 4740 7803 4743
rect 7791 4712 9904 4740
rect 7791 4709 7803 4712
rect 7745 4703 7803 4709
rect 5718 4672 5724 4684
rect 5631 4644 5724 4672
rect 5718 4632 5724 4644
rect 5776 4672 5782 4684
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 5776 4644 6193 4672
rect 5776 4632 5782 4644
rect 6181 4641 6193 4644
rect 6227 4641 6239 4675
rect 6638 4672 6644 4684
rect 6599 4644 6644 4672
rect 6181 4635 6239 4641
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 7006 4672 7012 4684
rect 6967 4644 7012 4672
rect 7006 4632 7012 4644
rect 7064 4632 7070 4684
rect 7561 4675 7619 4681
rect 7561 4641 7573 4675
rect 7607 4672 7619 4675
rect 7837 4675 7895 4681
rect 7837 4672 7849 4675
rect 7607 4644 7849 4672
rect 7607 4641 7619 4644
rect 7561 4635 7619 4641
rect 7837 4641 7849 4644
rect 7883 4641 7895 4675
rect 7837 4635 7895 4641
rect 5552 4576 5902 4604
rect 4709 4567 4767 4573
rect 3881 4539 3939 4545
rect 3881 4505 3893 4539
rect 3927 4536 3939 4539
rect 5874 4536 5902 4576
rect 5994 4564 6000 4616
rect 6052 4604 6058 4616
rect 6362 4604 6368 4616
rect 6052 4576 6368 4604
rect 6052 4564 6058 4576
rect 6362 4564 6368 4576
rect 6420 4604 6426 4616
rect 7576 4604 7604 4635
rect 7926 4632 7932 4684
rect 7984 4672 7990 4684
rect 8608 4675 8666 4681
rect 8608 4672 8620 4675
rect 7984 4644 8620 4672
rect 7984 4632 7990 4644
rect 8608 4641 8620 4644
rect 8654 4641 8666 4675
rect 8608 4635 8666 4641
rect 8938 4632 8944 4684
rect 8996 4672 9002 4684
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8996 4644 9045 4672
rect 8996 4632 9002 4644
rect 9033 4641 9045 4644
rect 9079 4641 9091 4675
rect 9033 4635 9091 4641
rect 9214 4632 9220 4684
rect 9272 4672 9278 4684
rect 9876 4681 9904 4712
rect 11238 4700 11244 4752
rect 11296 4740 11302 4752
rect 11470 4743 11528 4749
rect 11470 4740 11482 4743
rect 11296 4712 11482 4740
rect 11296 4700 11302 4712
rect 11470 4709 11482 4712
rect 11516 4709 11528 4743
rect 12342 4740 12348 4752
rect 12303 4712 12348 4740
rect 11470 4703 11528 4709
rect 12342 4700 12348 4712
rect 12400 4700 12406 4752
rect 13906 4740 13912 4752
rect 13188 4712 13912 4740
rect 9677 4675 9735 4681
rect 9677 4672 9689 4675
rect 9272 4644 9689 4672
rect 9272 4632 9278 4644
rect 9677 4641 9689 4644
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 9861 4675 9919 4681
rect 9861 4641 9873 4675
rect 9907 4672 9919 4675
rect 10505 4675 10563 4681
rect 10505 4672 10517 4675
rect 9907 4644 10517 4672
rect 9907 4641 9919 4644
rect 9861 4635 9919 4641
rect 10505 4641 10517 4644
rect 10551 4641 10563 4675
rect 10505 4635 10563 4641
rect 11149 4675 11207 4681
rect 11149 4641 11161 4675
rect 11195 4672 11207 4675
rect 11698 4672 11704 4684
rect 11195 4644 11704 4672
rect 11195 4641 11207 4644
rect 11149 4635 11207 4641
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 13078 4632 13084 4684
rect 13136 4672 13142 4684
rect 13188 4681 13216 4712
rect 13906 4700 13912 4712
rect 13964 4700 13970 4752
rect 14642 4740 14648 4752
rect 14016 4712 14648 4740
rect 13173 4675 13231 4681
rect 13173 4672 13185 4675
rect 13136 4644 13185 4672
rect 13136 4632 13142 4644
rect 13173 4641 13185 4644
rect 13219 4641 13231 4675
rect 13354 4672 13360 4684
rect 13315 4644 13360 4672
rect 13173 4635 13231 4641
rect 13354 4632 13360 4644
rect 13412 4632 13418 4684
rect 13722 4632 13728 4684
rect 13780 4672 13786 4684
rect 13817 4675 13875 4681
rect 13817 4672 13829 4675
rect 13780 4644 13829 4672
rect 13780 4632 13786 4644
rect 13817 4641 13829 4644
rect 13863 4672 13875 4675
rect 14016 4672 14044 4712
rect 14642 4700 14648 4712
rect 14700 4700 14706 4752
rect 15120 4740 15148 4780
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 16022 4808 16028 4820
rect 15344 4780 16028 4808
rect 15344 4768 15350 4780
rect 16022 4768 16028 4780
rect 16080 4808 16086 4820
rect 17129 4811 17187 4817
rect 17129 4808 17141 4811
rect 16080 4780 17141 4808
rect 16080 4768 16086 4780
rect 17129 4777 17141 4780
rect 17175 4777 17187 4811
rect 18693 4811 18751 4817
rect 18693 4808 18705 4811
rect 17129 4771 17187 4777
rect 17236 4780 18705 4808
rect 15927 4743 15985 4749
rect 15120 4712 15675 4740
rect 13863 4644 14044 4672
rect 13863 4641 13875 4644
rect 13817 4635 13875 4641
rect 14090 4632 14096 4684
rect 14148 4672 14154 4684
rect 14277 4675 14335 4681
rect 14277 4672 14289 4675
rect 14148 4644 14289 4672
rect 14148 4632 14154 4644
rect 14277 4641 14289 4644
rect 14323 4672 14335 4675
rect 14918 4672 14924 4684
rect 14323 4644 14924 4672
rect 14323 4641 14335 4644
rect 14277 4635 14335 4641
rect 14918 4632 14924 4644
rect 14976 4672 14982 4684
rect 15102 4672 15108 4684
rect 14976 4644 15108 4672
rect 14976 4632 14982 4644
rect 15102 4632 15108 4644
rect 15160 4632 15166 4684
rect 15647 4672 15675 4712
rect 15927 4709 15939 4743
rect 15973 4740 15985 4743
rect 16114 4740 16120 4752
rect 15973 4712 16120 4740
rect 15973 4709 15985 4712
rect 15927 4703 15985 4709
rect 16114 4700 16120 4712
rect 16172 4700 16178 4752
rect 16298 4700 16304 4752
rect 16356 4740 16362 4752
rect 17236 4740 17264 4780
rect 18693 4777 18705 4780
rect 18739 4777 18751 4811
rect 18693 4771 18751 4777
rect 16356 4712 17264 4740
rect 16356 4700 16362 4712
rect 17402 4700 17408 4752
rect 17460 4740 17466 4752
rect 17497 4743 17555 4749
rect 17497 4740 17509 4743
rect 17460 4712 17509 4740
rect 17460 4700 17466 4712
rect 17497 4709 17509 4712
rect 17543 4709 17555 4743
rect 17497 4703 17555 4709
rect 16390 4672 16396 4684
rect 15647 4644 16396 4672
rect 16390 4632 16396 4644
rect 16448 4632 16454 4684
rect 16758 4672 16764 4684
rect 16719 4644 16764 4672
rect 16758 4632 16764 4644
rect 16816 4632 16822 4684
rect 19058 4672 19064 4684
rect 19019 4644 19064 4672
rect 19058 4632 19064 4644
rect 19116 4632 19122 4684
rect 6420 4576 7604 4604
rect 6420 4564 6426 4576
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 8168 4576 10241 4604
rect 8168 4564 8174 4576
rect 10229 4573 10241 4576
rect 10275 4604 10287 4607
rect 10318 4604 10324 4616
rect 10275 4576 10324 4604
rect 10275 4573 10287 4576
rect 10229 4567 10287 4573
rect 10318 4564 10324 4576
rect 10376 4564 10382 4616
rect 11716 4604 11744 4632
rect 13630 4604 13636 4616
rect 11716 4576 13636 4604
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4604 14427 4607
rect 15565 4607 15623 4613
rect 15565 4604 15577 4607
rect 14415 4576 15577 4604
rect 14415 4573 14427 4576
rect 14369 4567 14427 4573
rect 15565 4573 15577 4576
rect 15611 4604 15623 4607
rect 16666 4604 16672 4616
rect 15611 4576 16672 4604
rect 15611 4573 15623 4576
rect 15565 4567 15623 4573
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 17402 4604 17408 4616
rect 17363 4576 17408 4604
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 17678 4604 17684 4616
rect 17639 4576 17684 4604
rect 17678 4564 17684 4576
rect 17736 4564 17742 4616
rect 17770 4564 17776 4616
rect 17828 4604 17834 4616
rect 18877 4607 18935 4613
rect 18877 4604 18889 4607
rect 17828 4576 18889 4604
rect 17828 4564 17834 4576
rect 18877 4573 18889 4576
rect 18923 4573 18935 4607
rect 18877 4567 18935 4573
rect 8846 4536 8852 4548
rect 3927 4508 4154 4536
rect 5874 4508 8852 4536
rect 3927 4505 3939 4508
rect 3881 4499 3939 4505
rect 4126 4468 4154 4508
rect 8846 4496 8852 4508
rect 8904 4496 8910 4548
rect 9306 4496 9312 4548
rect 9364 4536 9370 4548
rect 11330 4536 11336 4548
rect 9364 4508 11336 4536
rect 9364 4496 9370 4508
rect 11330 4496 11336 4508
rect 11388 4536 11394 4548
rect 12805 4539 12863 4545
rect 12805 4536 12817 4539
rect 11388 4508 12817 4536
rect 11388 4496 11394 4508
rect 12805 4505 12817 4508
rect 12851 4536 12863 4539
rect 13354 4536 13360 4548
rect 12851 4508 13360 4536
rect 12851 4505 12863 4508
rect 12805 4499 12863 4505
rect 13354 4496 13360 4508
rect 13412 4496 13418 4548
rect 16485 4539 16543 4545
rect 16485 4505 16497 4539
rect 16531 4536 16543 4539
rect 18230 4536 18236 4548
rect 16531 4508 18236 4536
rect 16531 4505 16543 4508
rect 16485 4499 16543 4505
rect 18230 4496 18236 4508
rect 18288 4536 18294 4548
rect 18325 4539 18383 4545
rect 18325 4536 18337 4539
rect 18288 4508 18337 4536
rect 18288 4496 18294 4508
rect 18325 4505 18337 4508
rect 18371 4505 18383 4539
rect 18325 4499 18383 4505
rect 5534 4468 5540 4480
rect 4126 4440 5540 4468
rect 5534 4428 5540 4440
rect 5592 4468 5598 4480
rect 7745 4471 7803 4477
rect 7745 4468 7757 4471
rect 5592 4440 7757 4468
rect 5592 4428 5598 4440
rect 7745 4437 7757 4440
rect 7791 4437 7803 4471
rect 7745 4431 7803 4437
rect 7837 4471 7895 4477
rect 7837 4437 7849 4471
rect 7883 4468 7895 4471
rect 8021 4471 8079 4477
rect 8021 4468 8033 4471
rect 7883 4440 8033 4468
rect 7883 4437 7895 4440
rect 7837 4431 7895 4437
rect 8021 4437 8033 4440
rect 8067 4468 8079 4471
rect 8570 4468 8576 4480
rect 8067 4440 8576 4468
rect 8067 4437 8079 4440
rect 8021 4431 8079 4437
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 8711 4471 8769 4477
rect 8711 4437 8723 4471
rect 8757 4468 8769 4471
rect 8938 4468 8944 4480
rect 8757 4440 8944 4468
rect 8757 4437 8769 4440
rect 8711 4431 8769 4437
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 10594 4428 10600 4480
rect 10652 4468 10658 4480
rect 15102 4468 15108 4480
rect 10652 4440 15108 4468
rect 10652 4428 10658 4440
rect 15102 4428 15108 4440
rect 15160 4428 15166 4480
rect 1104 4378 20884 4400
rect 1104 4326 4648 4378
rect 4700 4326 4712 4378
rect 4764 4326 4776 4378
rect 4828 4326 4840 4378
rect 4892 4326 11982 4378
rect 12034 4326 12046 4378
rect 12098 4326 12110 4378
rect 12162 4326 12174 4378
rect 12226 4326 19315 4378
rect 19367 4326 19379 4378
rect 19431 4326 19443 4378
rect 19495 4326 19507 4378
rect 19559 4326 20884 4378
rect 1104 4304 20884 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2685 4267 2743 4273
rect 2685 4264 2697 4267
rect 2464 4236 2697 4264
rect 2464 4224 2470 4236
rect 2685 4233 2697 4236
rect 2731 4233 2743 4267
rect 2685 4227 2743 4233
rect 2958 4224 2964 4276
rect 3016 4264 3022 4276
rect 3053 4267 3111 4273
rect 3053 4264 3065 4267
rect 3016 4236 3065 4264
rect 3016 4224 3022 4236
rect 3053 4233 3065 4236
rect 3099 4233 3111 4267
rect 3053 4227 3111 4233
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 5629 4267 5687 4273
rect 5629 4264 5641 4267
rect 4120 4236 5641 4264
rect 4120 4224 4126 4236
rect 5629 4233 5641 4236
rect 5675 4233 5687 4267
rect 5629 4227 5687 4233
rect 5718 4224 5724 4276
rect 5776 4264 5782 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 5776 4236 6561 4264
rect 5776 4224 5782 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 12621 4267 12679 4273
rect 12621 4233 12633 4267
rect 12667 4264 12679 4267
rect 12667 4236 13584 4264
rect 12667 4233 12679 4236
rect 12621 4227 12679 4233
rect 4890 4156 4896 4208
rect 4948 4196 4954 4208
rect 5810 4196 5816 4208
rect 4948 4168 5816 4196
rect 4948 4156 4954 4168
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 7466 4156 7472 4208
rect 7524 4196 7530 4208
rect 7653 4199 7711 4205
rect 7653 4196 7665 4199
rect 7524 4168 7665 4196
rect 7524 4156 7530 4168
rect 7653 4165 7665 4168
rect 7699 4196 7711 4199
rect 8202 4196 8208 4208
rect 7699 4168 8208 4196
rect 7699 4165 7711 4168
rect 7653 4159 7711 4165
rect 1762 4128 1768 4140
rect 1723 4100 1768 4128
rect 1762 4088 1768 4100
rect 1820 4088 1826 4140
rect 5534 4128 5540 4140
rect 5495 4100 5540 4128
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4128 5687 4131
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 5675 4100 7205 4128
rect 5675 4097 5687 4100
rect 5629 4091 5687 4097
rect 7193 4097 7205 4100
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 4709 4063 4767 4069
rect 4709 4060 4721 4063
rect 4126 4032 4721 4060
rect 1854 3992 1860 4004
rect 1815 3964 1860 3992
rect 1854 3952 1860 3964
rect 1912 3952 1918 4004
rect 2409 3995 2467 4001
rect 2409 3961 2421 3995
rect 2455 3992 2467 3995
rect 3050 3992 3056 4004
rect 2455 3964 3056 3992
rect 2455 3961 2467 3964
rect 2409 3955 2467 3961
rect 3050 3952 3056 3964
rect 3108 3992 3114 4004
rect 3329 3995 3387 4001
rect 3329 3992 3341 3995
rect 3108 3964 3341 3992
rect 3108 3952 3114 3964
rect 3329 3961 3341 3964
rect 3375 3961 3387 3995
rect 3329 3955 3387 3961
rect 3421 3995 3479 4001
rect 3421 3961 3433 3995
rect 3467 3992 3479 3995
rect 3602 3992 3608 4004
rect 3467 3964 3608 3992
rect 3467 3961 3479 3964
rect 3421 3955 3479 3961
rect 3602 3952 3608 3964
rect 3660 3952 3666 4004
rect 3970 3992 3976 4004
rect 3931 3964 3976 3992
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 3878 3884 3884 3936
rect 3936 3924 3942 3936
rect 4126 3924 4154 4032
rect 4709 4029 4721 4032
rect 4755 4060 4767 4063
rect 5445 4063 5503 4069
rect 5445 4060 5457 4063
rect 4755 4032 5457 4060
rect 4755 4029 4767 4032
rect 4709 4023 4767 4029
rect 5445 4029 5457 4032
rect 5491 4060 5503 4063
rect 6546 4060 6552 4072
rect 5491 4032 6552 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 4338 3992 4344 4004
rect 4251 3964 4344 3992
rect 4338 3952 4344 3964
rect 4396 3992 4402 4004
rect 5994 3992 6000 4004
rect 4396 3964 6000 3992
rect 4396 3952 4402 3964
rect 5994 3952 6000 3964
rect 6052 3952 6058 4004
rect 7208 3992 7236 4091
rect 7852 4069 7880 4168
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 9306 4156 9312 4208
rect 9364 4196 9370 4208
rect 11146 4196 11152 4208
rect 9364 4168 11152 4196
rect 9364 4156 9370 4168
rect 11146 4156 11152 4168
rect 11204 4156 11210 4208
rect 11790 4196 11796 4208
rect 11751 4168 11796 4196
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 13078 4196 13084 4208
rect 13039 4168 13084 4196
rect 13078 4156 13084 4168
rect 13136 4196 13142 4208
rect 13357 4199 13415 4205
rect 13357 4196 13369 4199
rect 13136 4168 13369 4196
rect 13136 4156 13142 4168
rect 13357 4165 13369 4168
rect 13403 4165 13415 4199
rect 13556 4196 13584 4236
rect 13630 4224 13636 4276
rect 13688 4264 13694 4276
rect 17221 4267 17279 4273
rect 17221 4264 17233 4267
rect 13688 4236 17233 4264
rect 13688 4224 13694 4236
rect 17221 4233 17233 4236
rect 17267 4233 17279 4267
rect 17221 4227 17279 4233
rect 17865 4267 17923 4273
rect 17865 4233 17877 4267
rect 17911 4264 17923 4267
rect 18138 4264 18144 4276
rect 17911 4236 18144 4264
rect 17911 4233 17923 4236
rect 17865 4227 17923 4233
rect 18138 4224 18144 4236
rect 18196 4264 18202 4276
rect 18196 4224 18230 4264
rect 18782 4224 18788 4276
rect 18840 4264 18846 4276
rect 19058 4264 19064 4276
rect 18840 4236 19064 4264
rect 18840 4224 18846 4236
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 14090 4196 14096 4208
rect 13556 4168 14096 4196
rect 13357 4159 13415 4165
rect 14090 4156 14096 4168
rect 14148 4156 14154 4208
rect 15286 4196 15292 4208
rect 15247 4168 15292 4196
rect 15286 4156 15292 4168
rect 15344 4156 15350 4208
rect 15470 4156 15476 4208
rect 15528 4196 15534 4208
rect 17402 4196 17408 4208
rect 15528 4168 17408 4196
rect 15528 4156 15534 4168
rect 17402 4156 17408 4168
rect 17460 4156 17466 4208
rect 18202 4196 18230 4224
rect 19610 4196 19616 4208
rect 18202 4168 19616 4196
rect 19610 4156 19616 4168
rect 19668 4156 19674 4208
rect 8846 4088 8852 4140
rect 8904 4128 8910 4140
rect 12158 4128 12164 4140
rect 8904 4100 11008 4128
rect 12119 4100 12164 4128
rect 8904 4088 8910 4100
rect 7837 4063 7895 4069
rect 7837 4029 7849 4063
rect 7883 4029 7895 4063
rect 7837 4023 7895 4029
rect 8205 4063 8263 4069
rect 8205 4029 8217 4063
rect 8251 4029 8263 4063
rect 8570 4060 8576 4072
rect 8531 4032 8576 4060
rect 8205 4023 8263 4029
rect 8018 3992 8024 4004
rect 7208 3964 8024 3992
rect 8018 3952 8024 3964
rect 8076 3992 8082 4004
rect 8220 3992 8248 4023
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 9122 4060 9128 4072
rect 9035 4032 9128 4060
rect 9122 4020 9128 4032
rect 9180 4060 9186 4072
rect 9490 4060 9496 4072
rect 9180 4032 9496 4060
rect 9180 4020 9186 4032
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 10980 4069 11008 4100
rect 12158 4088 12164 4100
rect 12216 4128 12222 4140
rect 16025 4131 16083 4137
rect 16025 4128 16037 4131
rect 12216 4100 12480 4128
rect 12216 4088 12222 4100
rect 12452 4069 12480 4100
rect 12544 4100 16037 4128
rect 10045 4063 10103 4069
rect 10045 4029 10057 4063
rect 10091 4060 10103 4063
rect 10965 4063 11023 4069
rect 10091 4032 10916 4060
rect 10091 4029 10103 4032
rect 10045 4023 10103 4029
rect 8076 3964 8248 3992
rect 8076 3952 8082 3964
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 10060 3992 10088 4023
rect 9088 3964 10088 3992
rect 10366 3995 10424 4001
rect 9088 3952 9094 3964
rect 10366 3961 10378 3995
rect 10412 3961 10424 3995
rect 10888 3992 10916 4032
rect 10965 4029 10977 4063
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 12544 3992 12572 4100
rect 16025 4097 16037 4100
rect 16071 4097 16083 4131
rect 16025 4091 16083 4097
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4128 17003 4131
rect 17678 4128 17684 4140
rect 16991 4100 17684 4128
rect 16991 4097 17003 4100
rect 16945 4091 17003 4097
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 18138 4128 18144 4140
rect 18099 4100 18144 4128
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 18785 4131 18843 4137
rect 18785 4097 18797 4131
rect 18831 4128 18843 4131
rect 18874 4128 18880 4140
rect 18831 4100 18880 4128
rect 18831 4097 18843 4100
rect 18785 4091 18843 4097
rect 18874 4088 18880 4100
rect 18932 4088 18938 4140
rect 13906 4060 13912 4072
rect 13867 4032 13912 4060
rect 13906 4020 13912 4032
rect 13964 4020 13970 4072
rect 14366 4060 14372 4072
rect 14327 4032 14372 4060
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 14826 4060 14832 4072
rect 14787 4032 14832 4060
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 14918 4020 14924 4072
rect 14976 4060 14982 4072
rect 15105 4063 15163 4069
rect 15105 4060 15117 4063
rect 14976 4032 15117 4060
rect 14976 4020 14982 4032
rect 15105 4029 15117 4032
rect 15151 4029 15163 4063
rect 19610 4060 19616 4072
rect 19574 4032 19616 4060
rect 15105 4023 15163 4029
rect 19610 4020 19616 4032
rect 19668 4069 19674 4072
rect 19668 4063 19722 4069
rect 19668 4029 19676 4063
rect 19710 4060 19722 4063
rect 20073 4063 20131 4069
rect 20073 4060 20085 4063
rect 19710 4032 20085 4060
rect 19710 4029 19722 4032
rect 19668 4023 19722 4029
rect 20073 4029 20085 4032
rect 20119 4029 20131 4063
rect 20073 4023 20131 4029
rect 19668 4020 19674 4023
rect 10888 3964 12572 3992
rect 10366 3955 10424 3961
rect 6178 3924 6184 3936
rect 3936 3896 4154 3924
rect 6139 3896 6184 3924
rect 3936 3884 3942 3896
rect 6178 3884 6184 3896
rect 6236 3924 6242 3936
rect 6638 3924 6644 3936
rect 6236 3896 6644 3924
rect 6236 3884 6242 3896
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 7834 3924 7840 3936
rect 7795 3896 7840 3924
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 7984 3896 9505 3924
rect 7984 3884 7990 3896
rect 9493 3893 9505 3896
rect 9539 3924 9551 3927
rect 9582 3924 9588 3936
rect 9539 3896 9588 3924
rect 9539 3893 9551 3896
rect 9493 3887 9551 3893
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 9858 3924 9864 3936
rect 9819 3896 9864 3924
rect 9858 3884 9864 3896
rect 9916 3924 9922 3936
rect 10381 3924 10409 3955
rect 12618 3952 12624 4004
rect 12676 3992 12682 4004
rect 13538 3992 13544 4004
rect 12676 3964 13544 3992
rect 12676 3952 12682 3964
rect 13538 3952 13544 3964
rect 13596 3992 13602 4004
rect 16298 3992 16304 4004
rect 13596 3964 16304 3992
rect 13596 3952 13602 3964
rect 16298 3952 16304 3964
rect 16356 3952 16362 4004
rect 16390 3952 16396 4004
rect 16448 3992 16454 4004
rect 18230 3992 18236 4004
rect 16448 3964 16493 3992
rect 18191 3964 18236 3992
rect 16448 3952 16454 3964
rect 18230 3952 18236 3964
rect 18288 3952 18294 4004
rect 19751 3995 19809 4001
rect 19751 3961 19763 3995
rect 19797 3992 19809 3995
rect 20162 3992 20168 4004
rect 19797 3964 20168 3992
rect 19797 3961 19809 3964
rect 19751 3955 19809 3961
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 11238 3924 11244 3936
rect 9916 3896 11244 3924
rect 9916 3884 9922 3896
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 13817 3927 13875 3933
rect 13817 3924 13829 3927
rect 11756 3896 13829 3924
rect 11756 3884 11762 3896
rect 13817 3893 13829 3896
rect 13863 3924 13875 3927
rect 14826 3924 14832 3936
rect 13863 3896 14832 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 15378 3884 15384 3936
rect 15436 3924 15442 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 15436 3896 15669 3924
rect 15436 3884 15442 3896
rect 15657 3893 15669 3896
rect 15703 3893 15715 3927
rect 15657 3887 15715 3893
rect 17402 3884 17408 3936
rect 17460 3924 17466 3936
rect 19429 3927 19487 3933
rect 19429 3924 19441 3927
rect 17460 3896 19441 3924
rect 17460 3884 17466 3896
rect 19429 3893 19441 3896
rect 19475 3893 19487 3927
rect 19429 3887 19487 3893
rect 1104 3834 20884 3856
rect 1104 3782 8315 3834
rect 8367 3782 8379 3834
rect 8431 3782 8443 3834
rect 8495 3782 8507 3834
rect 8559 3782 15648 3834
rect 15700 3782 15712 3834
rect 15764 3782 15776 3834
rect 15828 3782 15840 3834
rect 15892 3782 20884 3834
rect 1104 3760 20884 3782
rect 1854 3680 1860 3732
rect 1912 3720 1918 3732
rect 2869 3723 2927 3729
rect 2869 3720 2881 3723
rect 1912 3692 2881 3720
rect 1912 3680 1918 3692
rect 2869 3689 2881 3692
rect 2915 3689 2927 3723
rect 2869 3683 2927 3689
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 3016 3692 3433 3720
rect 3016 3680 3022 3692
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 3421 3683 3479 3689
rect 3881 3723 3939 3729
rect 3881 3689 3893 3723
rect 3927 3720 3939 3723
rect 4338 3720 4344 3732
rect 3927 3692 4344 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 4890 3720 4896 3732
rect 4851 3692 4896 3720
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 5077 3723 5135 3729
rect 5077 3689 5089 3723
rect 5123 3689 5135 3723
rect 5077 3683 5135 3689
rect 2314 3661 2320 3664
rect 2311 3652 2320 3661
rect 2275 3624 2320 3652
rect 2311 3615 2320 3624
rect 2314 3612 2320 3615
rect 2372 3612 2378 3664
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 5092 3652 5120 3683
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 7377 3723 7435 3729
rect 7377 3720 7389 3723
rect 5224 3692 7389 3720
rect 5224 3680 5230 3692
rect 7377 3689 7389 3692
rect 7423 3689 7435 3723
rect 7377 3683 7435 3689
rect 8938 3680 8944 3732
rect 8996 3720 9002 3732
rect 13262 3720 13268 3732
rect 8996 3692 13268 3720
rect 8996 3680 9002 3692
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 13998 3680 14004 3732
rect 14056 3720 14062 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 14056 3692 14289 3720
rect 14056 3680 14062 3692
rect 14277 3689 14289 3692
rect 14323 3720 14335 3723
rect 14366 3720 14372 3732
rect 14323 3692 14372 3720
rect 14323 3689 14335 3692
rect 14277 3683 14335 3689
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 14645 3723 14703 3729
rect 14645 3689 14657 3723
rect 14691 3720 14703 3723
rect 14918 3720 14924 3732
rect 14691 3692 14924 3720
rect 14691 3689 14703 3692
rect 14645 3683 14703 3689
rect 14918 3680 14924 3692
rect 14976 3680 14982 3732
rect 16390 3720 16396 3732
rect 16351 3692 16396 3720
rect 16390 3680 16396 3692
rect 16448 3680 16454 3732
rect 16666 3720 16672 3732
rect 16627 3692 16672 3720
rect 16666 3680 16672 3692
rect 16724 3680 16730 3732
rect 17678 3680 17684 3732
rect 17736 3720 17742 3732
rect 19429 3723 19487 3729
rect 19429 3720 19441 3723
rect 17736 3692 19441 3720
rect 17736 3680 17742 3692
rect 19429 3689 19441 3692
rect 19475 3720 19487 3723
rect 19610 3720 19616 3732
rect 19475 3692 19616 3720
rect 19475 3689 19487 3692
rect 19429 3683 19487 3689
rect 19610 3680 19616 3692
rect 19668 3680 19674 3732
rect 2832 3624 5120 3652
rect 5276 3624 6868 3652
rect 2832 3612 2838 3624
rect 5276 3596 5304 3624
rect 5074 3544 5080 3596
rect 5132 3584 5138 3596
rect 5258 3584 5264 3596
rect 5132 3556 5264 3584
rect 5132 3544 5138 3556
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3553 5503 3587
rect 5994 3584 6000 3596
rect 5955 3556 6000 3584
rect 5445 3547 5503 3553
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3516 2007 3519
rect 2038 3516 2044 3528
rect 1995 3488 2044 3516
rect 1995 3485 2007 3488
rect 1949 3479 2007 3485
rect 2038 3476 2044 3488
rect 2096 3516 2102 3528
rect 4522 3516 4528 3528
rect 2096 3488 4528 3516
rect 2096 3476 2102 3488
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 5460 3516 5488 3547
rect 5994 3544 6000 3556
rect 6052 3544 6058 3596
rect 6362 3584 6368 3596
rect 6323 3556 6368 3584
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 6840 3593 6868 3624
rect 7098 3612 7104 3664
rect 7156 3652 7162 3664
rect 9033 3655 9091 3661
rect 9033 3652 9045 3655
rect 7156 3624 9045 3652
rect 7156 3612 7162 3624
rect 9033 3621 9045 3624
rect 9079 3652 9091 3655
rect 9214 3652 9220 3664
rect 9079 3624 9220 3652
rect 9079 3621 9091 3624
rect 9033 3615 9091 3621
rect 9214 3612 9220 3624
rect 9272 3652 9278 3664
rect 9493 3655 9551 3661
rect 9493 3652 9505 3655
rect 9272 3624 9505 3652
rect 9272 3612 9278 3624
rect 9493 3621 9505 3624
rect 9539 3621 9551 3655
rect 9493 3615 9551 3621
rect 10686 3612 10692 3664
rect 10744 3652 10750 3664
rect 13357 3655 13415 3661
rect 13357 3652 13369 3655
rect 10744 3624 13369 3652
rect 10744 3612 10750 3624
rect 13357 3621 13369 3624
rect 13403 3652 13415 3655
rect 15010 3652 15016 3664
rect 13403 3624 15016 3652
rect 13403 3621 13415 3624
rect 13357 3615 13415 3621
rect 15010 3612 15016 3624
rect 15068 3652 15074 3664
rect 15473 3655 15531 3661
rect 15473 3652 15485 3655
rect 15068 3624 15485 3652
rect 15068 3612 15074 3624
rect 15473 3621 15485 3624
rect 15519 3621 15531 3655
rect 15473 3615 15531 3621
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 17221 3655 17279 3661
rect 17221 3652 17233 3655
rect 17184 3624 17233 3652
rect 17184 3612 17190 3624
rect 17221 3621 17233 3624
rect 17267 3652 17279 3655
rect 17770 3652 17776 3664
rect 17267 3624 17776 3652
rect 17267 3621 17279 3624
rect 17221 3615 17279 3621
rect 17770 3612 17776 3624
rect 17828 3612 17834 3664
rect 18690 3612 18696 3664
rect 18748 3652 18754 3664
rect 18785 3655 18843 3661
rect 18785 3652 18797 3655
rect 18748 3624 18797 3652
rect 18748 3612 18754 3624
rect 18785 3621 18797 3624
rect 18831 3621 18843 3655
rect 18785 3615 18843 3621
rect 6825 3587 6883 3593
rect 6825 3553 6837 3587
rect 6871 3584 6883 3587
rect 6914 3584 6920 3596
rect 6871 3556 6920 3584
rect 6871 3553 6883 3556
rect 6825 3547 6883 3553
rect 6914 3544 6920 3556
rect 6972 3584 6978 3596
rect 7285 3587 7343 3593
rect 7285 3584 7297 3587
rect 6972 3556 7297 3584
rect 6972 3544 6978 3556
rect 7285 3553 7297 3556
rect 7331 3553 7343 3587
rect 7285 3547 7343 3553
rect 7745 3587 7803 3593
rect 7745 3553 7757 3587
rect 7791 3553 7803 3587
rect 8110 3584 8116 3596
rect 8023 3556 8116 3584
rect 7745 3547 7803 3553
rect 5000 3488 5488 3516
rect 5000 3392 5028 3488
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 7101 3519 7159 3525
rect 7101 3516 7113 3519
rect 6696 3488 7113 3516
rect 6696 3476 6702 3488
rect 7101 3485 7113 3488
rect 7147 3516 7159 3519
rect 7760 3516 7788 3547
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3584 8723 3587
rect 8754 3584 8760 3596
rect 8711 3556 8760 3584
rect 8711 3553 8723 3556
rect 8665 3547 8723 3553
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 9398 3544 9404 3596
rect 9456 3584 9462 3596
rect 9769 3587 9827 3593
rect 9769 3584 9781 3587
rect 9456 3556 9781 3584
rect 9456 3544 9462 3556
rect 9769 3553 9781 3556
rect 9815 3584 9827 3587
rect 10042 3584 10048 3596
rect 9815 3556 10048 3584
rect 9815 3553 9827 3556
rect 9769 3547 9827 3553
rect 10042 3544 10048 3556
rect 10100 3544 10106 3596
rect 11146 3584 11152 3596
rect 11107 3556 11152 3584
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 11330 3584 11336 3596
rect 11291 3556 11336 3584
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 11698 3584 11704 3596
rect 11485 3556 11704 3584
rect 7147 3488 7788 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 7006 3408 7012 3460
rect 7064 3448 7070 3460
rect 7742 3448 7748 3460
rect 7064 3420 7748 3448
rect 7064 3408 7070 3420
rect 7742 3408 7748 3420
rect 7800 3448 7806 3460
rect 8128 3448 8156 3544
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 10781 3519 10839 3525
rect 10781 3516 10793 3519
rect 8260 3488 10793 3516
rect 8260 3476 8266 3488
rect 10781 3485 10793 3488
rect 10827 3485 10839 3519
rect 10781 3479 10839 3485
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 11485 3516 11513 3556
rect 11698 3544 11704 3556
rect 11756 3544 11762 3596
rect 11790 3544 11796 3596
rect 11848 3584 11854 3596
rect 12253 3587 12311 3593
rect 12253 3584 12265 3587
rect 11848 3556 12265 3584
rect 11848 3544 11854 3556
rect 12253 3553 12265 3556
rect 12299 3584 12311 3587
rect 12805 3587 12863 3593
rect 12299 3556 12531 3584
rect 12299 3553 12311 3556
rect 12253 3547 12311 3553
rect 12342 3516 12348 3528
rect 11020 3488 11513 3516
rect 12303 3488 12348 3516
rect 11020 3476 11026 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 7800 3420 8156 3448
rect 9953 3451 10011 3457
rect 7800 3408 7806 3420
rect 9953 3417 9965 3451
rect 9999 3448 10011 3451
rect 12503 3448 12531 3556
rect 12805 3553 12817 3587
rect 12851 3584 12863 3587
rect 13078 3584 13084 3596
rect 12851 3556 13084 3584
rect 12851 3553 12863 3556
rect 12805 3547 12863 3553
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 13262 3516 13268 3528
rect 13223 3488 13268 3516
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 13538 3516 13544 3528
rect 13499 3488 13544 3516
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 15102 3476 15108 3528
rect 15160 3516 15166 3528
rect 15381 3519 15439 3525
rect 15381 3516 15393 3519
rect 15160 3488 15393 3516
rect 15160 3476 15166 3488
rect 15381 3485 15393 3488
rect 15427 3485 15439 3519
rect 15381 3479 15439 3485
rect 12802 3448 12808 3460
rect 9999 3420 11513 3448
rect 12503 3420 12808 3448
rect 9999 3417 10011 3420
rect 9953 3411 10011 3417
rect 1762 3380 1768 3392
rect 1723 3352 1768 3380
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 4430 3340 4436 3392
rect 4488 3380 4494 3392
rect 4525 3383 4583 3389
rect 4525 3380 4537 3383
rect 4488 3352 4537 3380
rect 4488 3340 4494 3352
rect 4525 3349 4537 3352
rect 4571 3380 4583 3383
rect 4982 3380 4988 3392
rect 4571 3352 4988 3380
rect 4571 3349 4583 3352
rect 4525 3343 4583 3349
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 9858 3340 9864 3392
rect 9916 3380 9922 3392
rect 10597 3383 10655 3389
rect 10597 3380 10609 3383
rect 9916 3352 10609 3380
rect 9916 3340 9922 3352
rect 10597 3349 10609 3352
rect 10643 3349 10655 3383
rect 10597 3343 10655 3349
rect 10781 3383 10839 3389
rect 10781 3349 10793 3383
rect 10827 3380 10839 3383
rect 11146 3380 11152 3392
rect 10827 3352 11152 3380
rect 10827 3349 10839 3352
rect 10781 3343 10839 3349
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 11485 3380 11513 3420
rect 12802 3408 12808 3420
rect 12860 3448 12866 3460
rect 13814 3448 13820 3460
rect 12860 3420 13820 3448
rect 12860 3408 12866 3420
rect 13814 3408 13820 3420
rect 13872 3408 13878 3460
rect 15396 3448 15424 3479
rect 15470 3476 15476 3528
rect 15528 3516 15534 3528
rect 15657 3519 15715 3525
rect 15657 3516 15669 3519
rect 15528 3488 15669 3516
rect 15528 3476 15534 3488
rect 15657 3485 15669 3488
rect 15703 3485 15715 3519
rect 15657 3479 15715 3485
rect 16945 3519 17003 3525
rect 16945 3485 16957 3519
rect 16991 3516 17003 3519
rect 17129 3519 17187 3525
rect 17129 3516 17141 3519
rect 16991 3488 17141 3516
rect 16991 3485 17003 3488
rect 16945 3479 17003 3485
rect 17129 3485 17141 3488
rect 17175 3485 17187 3519
rect 18693 3519 18751 3525
rect 17129 3479 17187 3485
rect 17512 3488 18552 3516
rect 17512 3448 17540 3488
rect 17678 3448 17684 3460
rect 15396 3420 17540 3448
rect 17639 3420 17684 3448
rect 17678 3408 17684 3420
rect 17736 3408 17742 3460
rect 17770 3408 17776 3460
rect 17828 3448 17834 3460
rect 18417 3451 18475 3457
rect 18417 3448 18429 3451
rect 17828 3420 18429 3448
rect 17828 3408 17834 3420
rect 18417 3417 18429 3420
rect 18463 3417 18475 3451
rect 18417 3411 18475 3417
rect 11698 3380 11704 3392
rect 11485 3352 11704 3380
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 16945 3383 17003 3389
rect 16945 3349 16957 3383
rect 16991 3380 17003 3383
rect 17218 3380 17224 3392
rect 16991 3352 17224 3380
rect 16991 3349 17003 3352
rect 16945 3343 17003 3349
rect 17218 3340 17224 3352
rect 17276 3340 17282 3392
rect 17310 3340 17316 3392
rect 17368 3380 17374 3392
rect 17586 3380 17592 3392
rect 17368 3352 17592 3380
rect 17368 3340 17374 3352
rect 17586 3340 17592 3352
rect 17644 3380 17650 3392
rect 18049 3383 18107 3389
rect 18049 3380 18061 3383
rect 17644 3352 18061 3380
rect 17644 3340 17650 3352
rect 18049 3349 18061 3352
rect 18095 3349 18107 3383
rect 18524 3380 18552 3488
rect 18693 3485 18705 3519
rect 18739 3516 18751 3519
rect 18874 3516 18880 3528
rect 18739 3488 18880 3516
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 18874 3476 18880 3488
rect 18932 3476 18938 3528
rect 19613 3383 19671 3389
rect 19613 3380 19625 3383
rect 18524 3352 19625 3380
rect 18049 3343 18107 3349
rect 19613 3349 19625 3352
rect 19659 3349 19671 3383
rect 19613 3343 19671 3349
rect 1104 3290 20884 3312
rect 1104 3238 4648 3290
rect 4700 3238 4712 3290
rect 4764 3238 4776 3290
rect 4828 3238 4840 3290
rect 4892 3238 11982 3290
rect 12034 3238 12046 3290
rect 12098 3238 12110 3290
rect 12162 3238 12174 3290
rect 12226 3238 19315 3290
rect 19367 3238 19379 3290
rect 19431 3238 19443 3290
rect 19495 3238 19507 3290
rect 19559 3238 20884 3290
rect 1104 3216 20884 3238
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 2004 3148 2145 3176
rect 2004 3136 2010 3148
rect 2133 3145 2145 3148
rect 2179 3145 2191 3179
rect 3602 3176 3608 3188
rect 3563 3148 3608 3176
rect 2133 3139 2191 3145
rect 3602 3136 3608 3148
rect 3660 3136 3666 3188
rect 3694 3136 3700 3188
rect 3752 3176 3758 3188
rect 4249 3179 4307 3185
rect 4249 3176 4261 3179
rect 3752 3148 4261 3176
rect 3752 3136 3758 3148
rect 4249 3145 4261 3148
rect 4295 3145 4307 3179
rect 4249 3139 4307 3145
rect 1811 3111 1869 3117
rect 1811 3077 1823 3111
rect 1857 3108 1869 3111
rect 2682 3108 2688 3120
rect 1857 3080 2688 3108
rect 1857 3077 1869 3080
rect 1811 3071 1869 3077
rect 2682 3068 2688 3080
rect 2740 3068 2746 3120
rect 4264 3040 4292 3139
rect 5994 3136 6000 3188
rect 6052 3176 6058 3188
rect 7101 3179 7159 3185
rect 7101 3176 7113 3179
rect 6052 3148 7113 3176
rect 6052 3136 6058 3148
rect 7101 3145 7113 3148
rect 7147 3145 7159 3179
rect 7101 3139 7159 3145
rect 7745 3179 7803 3185
rect 7745 3145 7757 3179
rect 7791 3176 7803 3179
rect 8113 3179 8171 3185
rect 8113 3176 8125 3179
rect 7791 3148 8125 3176
rect 7791 3145 7803 3148
rect 7745 3139 7803 3145
rect 8113 3145 8125 3148
rect 8159 3176 8171 3179
rect 8754 3176 8760 3188
rect 8159 3148 8760 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 8754 3136 8760 3148
rect 8812 3176 8818 3188
rect 10042 3176 10048 3188
rect 8812 3148 9674 3176
rect 10003 3148 10048 3176
rect 8812 3136 8818 3148
rect 4982 3068 4988 3120
rect 5040 3108 5046 3120
rect 6178 3108 6184 3120
rect 5040 3080 6184 3108
rect 5040 3068 5046 3080
rect 6178 3068 6184 3080
rect 6236 3068 6242 3120
rect 4264 3012 5672 3040
rect 1740 2975 1798 2981
rect 1740 2941 1752 2975
rect 1786 2972 1798 2975
rect 1946 2972 1952 2984
rect 1786 2944 1952 2972
rect 1786 2941 1798 2944
rect 1740 2935 1798 2941
rect 1946 2932 1952 2944
rect 2004 2932 2010 2984
rect 2685 2975 2743 2981
rect 2685 2941 2697 2975
rect 2731 2972 2743 2975
rect 2774 2972 2780 2984
rect 2731 2944 2780 2972
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 3973 2975 4031 2981
rect 3973 2941 3985 2975
rect 4019 2972 4031 2975
rect 4709 2975 4767 2981
rect 4709 2972 4721 2975
rect 4019 2944 4721 2972
rect 4019 2941 4031 2944
rect 3973 2935 4031 2941
rect 4709 2941 4721 2944
rect 4755 2941 4767 2975
rect 4982 2972 4988 2984
rect 4943 2944 4988 2972
rect 4709 2935 4767 2941
rect 3006 2907 3064 2913
rect 3006 2873 3018 2907
rect 3052 2873 3064 2907
rect 3006 2867 3064 2873
rect 2314 2796 2320 2848
rect 2372 2836 2378 2848
rect 2501 2839 2559 2845
rect 2501 2836 2513 2839
rect 2372 2808 2513 2836
rect 2372 2796 2378 2808
rect 2501 2805 2513 2808
rect 2547 2836 2559 2839
rect 3021 2836 3049 2867
rect 4614 2864 4620 2916
rect 4672 2904 4678 2916
rect 4724 2904 4752 2935
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5644 2981 5672 3012
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 9646 3040 9674 3148
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 10505 3179 10563 3185
rect 10505 3145 10517 3179
rect 10551 3176 10563 3179
rect 10962 3176 10968 3188
rect 10551 3148 10968 3176
rect 10551 3145 10563 3148
rect 10505 3139 10563 3145
rect 10520 3040 10548 3139
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 11330 3136 11336 3188
rect 11388 3176 11394 3188
rect 11793 3179 11851 3185
rect 11793 3176 11805 3179
rect 11388 3148 11805 3176
rect 11388 3136 11394 3148
rect 11793 3145 11805 3148
rect 11839 3176 11851 3179
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 11839 3148 12173 3176
rect 11839 3145 11851 3148
rect 11793 3139 11851 3145
rect 12161 3145 12173 3148
rect 12207 3176 12219 3179
rect 12207 3148 13216 3176
rect 12207 3145 12219 3148
rect 12161 3139 12219 3145
rect 11146 3068 11152 3120
rect 11204 3108 11210 3120
rect 11204 3080 13032 3108
rect 11204 3068 11210 3080
rect 8076 3012 8800 3040
rect 8076 3000 8082 3012
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2941 5503 2975
rect 5445 2935 5503 2941
rect 5629 2975 5687 2981
rect 5629 2941 5641 2975
rect 5675 2941 5687 2975
rect 5629 2935 5687 2941
rect 5258 2904 5264 2916
rect 4672 2876 5264 2904
rect 4672 2864 4678 2876
rect 5258 2864 5264 2876
rect 5316 2864 5322 2916
rect 5460 2904 5488 2935
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 6641 2975 6699 2981
rect 6641 2972 6653 2975
rect 6604 2944 6653 2972
rect 6604 2932 6610 2944
rect 6641 2941 6653 2944
rect 6687 2972 6699 2975
rect 7009 2975 7067 2981
rect 7009 2972 7021 2975
rect 6687 2944 7021 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 7009 2941 7021 2944
rect 7055 2941 7067 2975
rect 7009 2935 7067 2941
rect 8202 2932 8208 2984
rect 8260 2972 8266 2984
rect 8772 2981 8800 3012
rect 9324 3012 10548 3040
rect 10597 3043 10655 3049
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 8260 2944 8309 2972
rect 8260 2932 8266 2944
rect 8297 2941 8309 2944
rect 8343 2941 8355 2975
rect 8297 2935 8355 2941
rect 8757 2975 8815 2981
rect 8757 2941 8769 2975
rect 8803 2972 8815 2975
rect 9030 2972 9036 2984
rect 8803 2944 9036 2972
rect 8803 2941 8815 2944
rect 8757 2935 8815 2941
rect 9030 2932 9036 2944
rect 9088 2932 9094 2984
rect 9324 2981 9352 3012
rect 10597 3009 10609 3043
rect 10643 3040 10655 3043
rect 12342 3040 12348 3052
rect 10643 3012 12348 3040
rect 10643 3009 10655 3012
rect 10597 3003 10655 3009
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2941 9367 2975
rect 9490 2972 9496 2984
rect 9451 2944 9496 2972
rect 9309 2935 9367 2941
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 13004 2981 13032 3080
rect 13188 3040 13216 3148
rect 13262 3136 13268 3188
rect 13320 3176 13326 3188
rect 15010 3176 15016 3188
rect 13320 3148 14228 3176
rect 14971 3148 15016 3176
rect 13320 3136 13326 3148
rect 14200 3108 14228 3148
rect 15010 3136 15016 3148
rect 15068 3136 15074 3188
rect 17126 3176 17132 3188
rect 17087 3148 17132 3176
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 17497 3179 17555 3185
rect 17497 3176 17509 3179
rect 17276 3148 17509 3176
rect 17276 3136 17282 3148
rect 17497 3145 17509 3148
rect 17543 3176 17555 3179
rect 19150 3176 19156 3188
rect 17543 3148 19156 3176
rect 17543 3145 17555 3148
rect 17497 3139 17555 3145
rect 19150 3136 19156 3148
rect 19208 3136 19214 3188
rect 20073 3111 20131 3117
rect 20073 3108 20085 3111
rect 14200 3080 20085 3108
rect 20073 3077 20085 3080
rect 20119 3077 20131 3111
rect 20073 3071 20131 3077
rect 13998 3040 14004 3052
rect 13188 3012 14004 3040
rect 11517 2975 11575 2981
rect 11517 2941 11529 2975
rect 11563 2972 11575 2975
rect 12989 2975 13047 2981
rect 11563 2944 12480 2972
rect 11563 2941 11575 2944
rect 11517 2935 11575 2941
rect 5994 2904 6000 2916
rect 5460 2876 6000 2904
rect 5994 2864 6000 2876
rect 6052 2864 6058 2916
rect 6825 2907 6883 2913
rect 6825 2873 6837 2907
rect 6871 2904 6883 2907
rect 7098 2904 7104 2916
rect 6871 2876 7104 2904
rect 6871 2873 6883 2876
rect 6825 2867 6883 2873
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 9766 2904 9772 2916
rect 9727 2876 9772 2904
rect 9766 2864 9772 2876
rect 9824 2864 9830 2916
rect 9858 2864 9864 2916
rect 9916 2904 9922 2916
rect 10918 2907 10976 2913
rect 10918 2904 10930 2907
rect 9916 2876 10930 2904
rect 9916 2864 9922 2876
rect 10918 2873 10930 2876
rect 10964 2904 10976 2907
rect 12250 2904 12256 2916
rect 10964 2876 12256 2904
rect 10964 2873 10976 2876
rect 10918 2867 10976 2873
rect 12250 2864 12256 2876
rect 12308 2864 12314 2916
rect 4522 2836 4528 2848
rect 2547 2808 3049 2836
rect 4483 2808 4528 2836
rect 2547 2805 2559 2808
rect 2501 2799 2559 2805
rect 4522 2796 4528 2808
rect 4580 2796 4586 2848
rect 12452 2836 12480 2944
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 13078 2972 13084 2984
rect 13035 2944 13084 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 13188 2981 13216 3012
rect 13998 3000 14004 3012
rect 14056 3000 14062 3052
rect 14182 3000 14188 3052
rect 14240 3040 14246 3052
rect 17310 3040 17316 3052
rect 14240 3012 17316 3040
rect 14240 3000 14246 3012
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 17678 3000 17684 3052
rect 17736 3040 17742 3052
rect 17736 3012 19707 3040
rect 17736 3000 17742 3012
rect 13173 2975 13231 2981
rect 13173 2941 13185 2975
rect 13219 2941 13231 2975
rect 13722 2972 13728 2984
rect 13683 2944 13728 2972
rect 13173 2935 13231 2941
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 13814 2932 13820 2984
rect 13872 2972 13878 2984
rect 14093 2975 14151 2981
rect 14093 2972 14105 2975
rect 13872 2944 14105 2972
rect 13872 2932 13878 2944
rect 14093 2941 14105 2944
rect 14139 2972 14151 2975
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 14139 2944 14473 2972
rect 14139 2941 14151 2944
rect 14093 2935 14151 2941
rect 14461 2941 14473 2944
rect 14507 2941 14519 2975
rect 14461 2935 14519 2941
rect 14918 2932 14924 2984
rect 14976 2972 14982 2984
rect 15565 2975 15623 2981
rect 15565 2972 15577 2975
rect 14976 2944 15577 2972
rect 14976 2932 14982 2944
rect 15565 2941 15577 2944
rect 15611 2972 15623 2975
rect 17770 2972 17776 2984
rect 15611 2944 17776 2972
rect 15611 2941 15623 2944
rect 15565 2935 15623 2941
rect 17770 2932 17776 2944
rect 17828 2932 17834 2984
rect 18966 2932 18972 2984
rect 19024 2972 19030 2984
rect 19679 2981 19707 3012
rect 19061 2975 19119 2981
rect 19061 2972 19073 2975
rect 19024 2944 19073 2972
rect 19024 2932 19030 2944
rect 19061 2941 19073 2944
rect 19107 2941 19119 2975
rect 19061 2935 19119 2941
rect 19664 2975 19722 2981
rect 19664 2941 19676 2975
rect 19710 2972 19722 2975
rect 20441 2975 20499 2981
rect 20441 2972 20453 2975
rect 19710 2944 20453 2972
rect 19710 2941 19722 2944
rect 19664 2935 19722 2941
rect 20441 2941 20453 2944
rect 20487 2941 20499 2975
rect 20441 2935 20499 2941
rect 13354 2864 13360 2916
rect 13412 2904 13418 2916
rect 13998 2904 14004 2916
rect 13412 2876 14004 2904
rect 13412 2864 13418 2876
rect 13998 2864 14004 2876
rect 14056 2904 14062 2916
rect 15378 2904 15384 2916
rect 14056 2876 15384 2904
rect 14056 2864 14062 2876
rect 15378 2864 15384 2876
rect 15436 2904 15442 2916
rect 15886 2907 15944 2913
rect 15886 2904 15898 2907
rect 15436 2876 15898 2904
rect 15436 2864 15442 2876
rect 15886 2873 15898 2876
rect 15932 2873 15944 2907
rect 17586 2904 17592 2916
rect 15886 2867 15944 2873
rect 16408 2876 17592 2904
rect 16408 2836 16436 2876
rect 17586 2864 17592 2876
rect 17644 2864 17650 2916
rect 17862 2864 17868 2916
rect 17920 2904 17926 2916
rect 18141 2907 18199 2913
rect 18141 2904 18153 2907
rect 17920 2876 18153 2904
rect 17920 2864 17926 2876
rect 18141 2873 18153 2876
rect 18187 2873 18199 2907
rect 18141 2867 18199 2873
rect 18233 2907 18291 2913
rect 18233 2873 18245 2907
rect 18279 2904 18291 2907
rect 18414 2904 18420 2916
rect 18279 2876 18420 2904
rect 18279 2873 18291 2876
rect 18233 2867 18291 2873
rect 12452 2808 16436 2836
rect 16485 2839 16543 2845
rect 16485 2805 16497 2839
rect 16531 2836 16543 2839
rect 16666 2836 16672 2848
rect 16531 2808 16672 2836
rect 16531 2805 16543 2808
rect 16485 2799 16543 2805
rect 16666 2796 16672 2808
rect 16724 2796 16730 2848
rect 17770 2836 17776 2848
rect 17731 2808 17776 2836
rect 17770 2796 17776 2808
rect 17828 2836 17834 2848
rect 18248 2836 18276 2867
rect 18414 2864 18420 2876
rect 18472 2864 18478 2916
rect 18782 2904 18788 2916
rect 18743 2876 18788 2904
rect 18782 2864 18788 2876
rect 18840 2864 18846 2916
rect 19751 2907 19809 2913
rect 19751 2873 19763 2907
rect 19797 2904 19809 2907
rect 21542 2904 21548 2916
rect 19797 2876 21548 2904
rect 19797 2873 19809 2876
rect 19751 2867 19809 2873
rect 21542 2864 21548 2876
rect 21600 2864 21606 2916
rect 19426 2836 19432 2848
rect 17828 2808 18276 2836
rect 19387 2808 19432 2836
rect 17828 2796 17834 2808
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 1104 2746 20884 2768
rect 1104 2694 8315 2746
rect 8367 2694 8379 2746
rect 8431 2694 8443 2746
rect 8495 2694 8507 2746
rect 8559 2694 15648 2746
rect 15700 2694 15712 2746
rect 15764 2694 15776 2746
rect 15828 2694 15840 2746
rect 15892 2694 20884 2746
rect 1104 2672 20884 2694
rect 1397 2635 1455 2641
rect 1397 2601 1409 2635
rect 1443 2632 1455 2635
rect 1762 2632 1768 2644
rect 1443 2604 1768 2632
rect 1443 2601 1455 2604
rect 1397 2595 1455 2601
rect 1762 2592 1768 2604
rect 1820 2632 1826 2644
rect 3510 2632 3516 2644
rect 1820 2604 2544 2632
rect 1820 2592 1826 2604
rect 2516 2573 2544 2604
rect 2608 2604 3516 2632
rect 2608 2573 2636 2604
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 3881 2635 3939 2641
rect 3881 2601 3893 2635
rect 3927 2632 3939 2635
rect 4614 2632 4620 2644
rect 3927 2604 4620 2632
rect 3927 2601 3939 2604
rect 3881 2595 3939 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 6362 2632 6368 2644
rect 6275 2604 6368 2632
rect 6362 2592 6368 2604
rect 6420 2632 6426 2644
rect 8297 2635 8355 2641
rect 6420 2604 8156 2632
rect 6420 2592 6426 2604
rect 2501 2567 2559 2573
rect 2501 2533 2513 2567
rect 2547 2533 2559 2567
rect 2501 2527 2559 2533
rect 2593 2567 2651 2573
rect 2593 2533 2605 2567
rect 2639 2533 2651 2567
rect 5398 2567 5456 2573
rect 5398 2564 5410 2567
rect 2593 2527 2651 2533
rect 4908 2536 5410 2564
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2496 3203 2499
rect 3970 2496 3976 2508
rect 3191 2468 3976 2496
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 3970 2456 3976 2468
rect 4028 2496 4034 2508
rect 4908 2505 4936 2536
rect 5398 2533 5410 2536
rect 5444 2564 5456 2567
rect 6089 2567 6147 2573
rect 6089 2564 6101 2567
rect 5444 2536 6101 2564
rect 5444 2533 5456 2536
rect 5398 2527 5456 2533
rect 6089 2533 6101 2536
rect 6135 2533 6147 2567
rect 6089 2527 6147 2533
rect 6178 2524 6184 2576
rect 6236 2564 6242 2576
rect 6641 2567 6699 2573
rect 6641 2564 6653 2567
rect 6236 2536 6653 2564
rect 6236 2524 6242 2536
rect 6641 2533 6653 2536
rect 6687 2564 6699 2567
rect 6687 2536 7420 2564
rect 6687 2533 6699 2536
rect 6641 2527 6699 2533
rect 4100 2499 4158 2505
rect 4100 2496 4112 2499
rect 4028 2468 4112 2496
rect 4028 2456 4034 2468
rect 4100 2465 4112 2468
rect 4146 2465 4158 2499
rect 4893 2499 4951 2505
rect 4893 2496 4905 2499
rect 4100 2459 4158 2465
rect 4724 2468 4905 2496
rect 2314 2388 2320 2440
rect 2372 2428 2378 2440
rect 4724 2428 4752 2468
rect 4893 2465 4905 2468
rect 4939 2465 4951 2499
rect 4893 2459 4951 2465
rect 5077 2499 5135 2505
rect 5077 2465 5089 2499
rect 5123 2496 5135 2499
rect 5166 2496 5172 2508
rect 5123 2468 5172 2496
rect 5123 2465 5135 2468
rect 5077 2459 5135 2465
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 6914 2496 6920 2508
rect 6875 2468 6920 2496
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7392 2505 7420 2536
rect 7377 2499 7435 2505
rect 7377 2465 7389 2499
rect 7423 2465 7435 2499
rect 7742 2496 7748 2508
rect 7703 2468 7748 2496
rect 7377 2459 7435 2465
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 8128 2505 8156 2604
rect 8297 2601 8309 2635
rect 8343 2632 8355 2635
rect 11514 2632 11520 2644
rect 8343 2604 11520 2632
rect 8343 2601 8355 2604
rect 8297 2595 8355 2601
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 11655 2635 11713 2641
rect 11655 2601 11667 2635
rect 11701 2632 11713 2635
rect 15611 2635 15669 2641
rect 11701 2604 15567 2632
rect 11701 2601 11713 2604
rect 11655 2595 11713 2601
rect 9030 2564 9036 2576
rect 8991 2536 9036 2564
rect 9030 2524 9036 2536
rect 9088 2524 9094 2576
rect 9858 2524 9864 2576
rect 9916 2564 9922 2576
rect 10090 2567 10148 2573
rect 10090 2564 10102 2567
rect 9916 2536 10102 2564
rect 9916 2524 9922 2536
rect 10090 2533 10102 2536
rect 10136 2533 10148 2567
rect 10090 2527 10148 2533
rect 10318 2524 10324 2576
rect 10376 2564 10382 2576
rect 12345 2567 12403 2573
rect 12345 2564 12357 2567
rect 10376 2536 12357 2564
rect 10376 2524 10382 2536
rect 12345 2533 12357 2536
rect 12391 2533 12403 2567
rect 12345 2527 12403 2533
rect 12897 2567 12955 2573
rect 12897 2533 12909 2567
rect 12943 2564 12955 2567
rect 13630 2564 13636 2576
rect 12943 2536 13636 2564
rect 12943 2533 12955 2536
rect 12897 2527 12955 2533
rect 13630 2524 13636 2536
rect 13688 2524 13694 2576
rect 13903 2567 13961 2573
rect 13903 2533 13915 2567
rect 13949 2564 13961 2567
rect 13998 2564 14004 2576
rect 13949 2536 14004 2564
rect 13949 2533 13961 2536
rect 13903 2527 13961 2533
rect 13998 2524 14004 2536
rect 14056 2524 14062 2576
rect 14829 2567 14887 2573
rect 14829 2533 14841 2567
rect 14875 2564 14887 2567
rect 15010 2564 15016 2576
rect 14875 2536 15016 2564
rect 14875 2533 14887 2536
rect 14829 2527 14887 2533
rect 15010 2524 15016 2536
rect 15068 2524 15074 2576
rect 15539 2564 15567 2604
rect 15611 2601 15623 2635
rect 15657 2632 15669 2635
rect 17862 2632 17868 2644
rect 15657 2604 17868 2632
rect 15657 2601 15669 2604
rect 15611 2595 15669 2601
rect 17862 2592 17868 2604
rect 17920 2632 17926 2644
rect 19705 2635 19763 2641
rect 19705 2632 19717 2635
rect 17920 2604 19717 2632
rect 17920 2592 17926 2604
rect 19705 2601 19717 2604
rect 19751 2601 19763 2635
rect 19705 2595 19763 2601
rect 16666 2564 16672 2576
rect 15539 2536 16436 2564
rect 16627 2536 16672 2564
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2465 8171 2499
rect 10686 2496 10692 2508
rect 10647 2468 10692 2496
rect 8113 2459 8171 2465
rect 10686 2456 10692 2468
rect 10744 2456 10750 2508
rect 11584 2499 11642 2505
rect 11584 2496 11596 2499
rect 10796 2468 11596 2496
rect 2372 2400 4752 2428
rect 4801 2431 4859 2437
rect 2372 2388 2378 2400
rect 4801 2397 4813 2431
rect 4847 2428 4859 2431
rect 8202 2428 8208 2440
rect 4847 2400 8208 2428
rect 4847 2397 4859 2400
rect 4801 2391 4859 2397
rect 8202 2388 8208 2400
rect 8260 2428 8266 2440
rect 8665 2431 8723 2437
rect 8665 2428 8677 2431
rect 8260 2400 8677 2428
rect 8260 2388 8266 2400
rect 8665 2397 8677 2400
rect 8711 2397 8723 2431
rect 9766 2428 9772 2440
rect 9679 2400 9772 2428
rect 8665 2391 8723 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 10134 2388 10140 2440
rect 10192 2428 10198 2440
rect 10796 2428 10824 2468
rect 11584 2465 11596 2468
rect 11630 2496 11642 2499
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 11630 2468 11897 2496
rect 11630 2465 11642 2468
rect 11584 2459 11642 2465
rect 11885 2465 11897 2468
rect 11931 2465 11943 2499
rect 11885 2459 11943 2465
rect 12250 2456 12256 2508
rect 12308 2496 12314 2508
rect 13354 2496 13360 2508
rect 12308 2468 13360 2496
rect 12308 2456 12314 2468
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 13541 2499 13599 2505
rect 13541 2465 13553 2499
rect 13587 2496 13599 2499
rect 14182 2496 14188 2508
rect 13587 2468 14188 2496
rect 13587 2465 13599 2468
rect 13541 2459 13599 2465
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14461 2499 14519 2505
rect 14461 2465 14473 2499
rect 14507 2496 14519 2499
rect 15378 2496 15384 2508
rect 14507 2468 15384 2496
rect 14507 2465 14519 2468
rect 14461 2459 14519 2465
rect 15378 2456 15384 2468
rect 15436 2456 15442 2508
rect 15562 2505 15568 2508
rect 15540 2499 15568 2505
rect 15540 2465 15552 2499
rect 15620 2496 15626 2508
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 15620 2468 16037 2496
rect 15540 2459 15568 2465
rect 15562 2456 15568 2459
rect 15620 2456 15626 2468
rect 16025 2465 16037 2468
rect 16071 2496 16083 2499
rect 16206 2496 16212 2508
rect 16071 2468 16212 2496
rect 16071 2465 16083 2468
rect 16025 2459 16083 2465
rect 16206 2456 16212 2468
rect 16264 2456 16270 2508
rect 10192 2400 10824 2428
rect 11057 2431 11115 2437
rect 10192 2388 10198 2400
rect 11057 2397 11069 2431
rect 11103 2428 11115 2431
rect 11146 2428 11152 2440
rect 11103 2400 11152 2428
rect 11103 2397 11115 2400
rect 11057 2391 11115 2397
rect 11146 2388 11152 2400
rect 11204 2388 11210 2440
rect 11425 2431 11483 2437
rect 11425 2397 11437 2431
rect 11471 2428 11483 2431
rect 11790 2428 11796 2440
rect 11471 2400 11796 2428
rect 11471 2397 11483 2400
rect 11425 2391 11483 2397
rect 11790 2388 11796 2400
rect 11848 2388 11854 2440
rect 12342 2388 12348 2440
rect 12400 2428 12406 2440
rect 16301 2431 16359 2437
rect 16301 2428 16313 2431
rect 12400 2400 16313 2428
rect 12400 2388 12406 2400
rect 16301 2397 16313 2400
rect 16347 2397 16359 2431
rect 16301 2391 16359 2397
rect 4203 2363 4261 2369
rect 4203 2329 4215 2363
rect 4249 2360 4261 2363
rect 6454 2360 6460 2372
rect 4249 2332 6460 2360
rect 4249 2329 4261 2332
rect 4203 2323 4261 2329
rect 6454 2320 6460 2332
rect 6512 2320 6518 2372
rect 9784 2360 9812 2388
rect 15105 2363 15163 2369
rect 15105 2360 15117 2363
rect 9784 2332 15117 2360
rect 15105 2329 15117 2332
rect 15151 2329 15163 2363
rect 16408 2360 16436 2536
rect 16666 2524 16672 2536
rect 16724 2524 16730 2576
rect 17221 2567 17279 2573
rect 17221 2533 17233 2567
rect 17267 2564 17279 2567
rect 17678 2564 17684 2576
rect 17267 2536 17684 2564
rect 17267 2533 17279 2536
rect 17221 2527 17279 2533
rect 17678 2524 17684 2536
rect 17736 2524 17742 2576
rect 18141 2567 18199 2573
rect 18141 2533 18153 2567
rect 18187 2564 18199 2567
rect 18506 2564 18512 2576
rect 18187 2536 18512 2564
rect 18187 2533 18199 2536
rect 18141 2527 18199 2533
rect 18506 2524 18512 2536
rect 18564 2524 18570 2576
rect 18874 2524 18880 2576
rect 18932 2564 18938 2576
rect 19337 2567 19395 2573
rect 19337 2564 19349 2567
rect 18932 2536 19349 2564
rect 18932 2524 18938 2536
rect 19337 2533 19349 2536
rect 19383 2533 19395 2567
rect 19337 2527 19395 2533
rect 17310 2456 17316 2508
rect 17368 2496 17374 2508
rect 17497 2499 17555 2505
rect 17497 2496 17509 2499
rect 17368 2468 17509 2496
rect 17368 2456 17374 2468
rect 17497 2465 17509 2468
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 16577 2431 16635 2437
rect 16577 2397 16589 2431
rect 16623 2428 16635 2431
rect 18414 2428 18420 2440
rect 16623 2400 18276 2428
rect 18375 2400 18420 2428
rect 16623 2397 16635 2400
rect 16577 2391 16635 2397
rect 18248 2360 18276 2400
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 18693 2431 18751 2437
rect 18693 2397 18705 2431
rect 18739 2428 18751 2431
rect 18782 2428 18788 2440
rect 18739 2400 18788 2428
rect 18739 2397 18751 2400
rect 18693 2391 18751 2397
rect 18708 2360 18736 2391
rect 18782 2388 18788 2400
rect 18840 2428 18846 2440
rect 20441 2431 20499 2437
rect 20441 2428 20453 2431
rect 18840 2400 20453 2428
rect 18840 2388 18846 2400
rect 20441 2397 20453 2400
rect 20487 2397 20499 2431
rect 20441 2391 20499 2397
rect 20073 2363 20131 2369
rect 20073 2360 20085 2363
rect 16408 2332 18184 2360
rect 18248 2332 18736 2360
rect 18800 2332 20085 2360
rect 15105 2323 15163 2329
rect 1762 2252 1768 2304
rect 1820 2292 1826 2304
rect 1949 2295 2007 2301
rect 1949 2292 1961 2295
rect 1820 2264 1961 2292
rect 1820 2252 1826 2264
rect 1949 2261 1961 2264
rect 1995 2292 2007 2295
rect 2314 2292 2320 2304
rect 1995 2264 2320 2292
rect 1995 2261 2007 2264
rect 1949 2255 2007 2261
rect 2314 2252 2320 2264
rect 2372 2252 2378 2304
rect 2774 2252 2780 2304
rect 2832 2292 2838 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 2832 2264 4813 2292
rect 2832 2252 2838 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 5994 2292 6000 2304
rect 5955 2264 6000 2292
rect 4801 2255 4859 2261
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 6089 2295 6147 2301
rect 6089 2261 6101 2295
rect 6135 2292 6147 2295
rect 9493 2295 9551 2301
rect 9493 2292 9505 2295
rect 6135 2264 9505 2292
rect 6135 2261 6147 2264
rect 6089 2255 6147 2261
rect 9493 2261 9505 2264
rect 9539 2292 9551 2295
rect 9858 2292 9864 2304
rect 9539 2264 9864 2292
rect 9539 2261 9551 2264
rect 9493 2255 9551 2261
rect 9858 2252 9864 2264
rect 9916 2252 9922 2304
rect 11885 2295 11943 2301
rect 11885 2261 11897 2295
rect 11931 2292 11943 2295
rect 12069 2295 12127 2301
rect 12069 2292 12081 2295
rect 11931 2264 12081 2292
rect 11931 2261 11943 2264
rect 11885 2255 11943 2261
rect 12069 2261 12081 2264
rect 12115 2292 12127 2295
rect 12342 2292 12348 2304
rect 12115 2264 12348 2292
rect 12115 2261 12127 2264
rect 12069 2255 12127 2261
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 18156 2292 18184 2332
rect 18414 2292 18420 2304
rect 18156 2264 18420 2292
rect 18414 2252 18420 2264
rect 18472 2292 18478 2304
rect 18800 2292 18828 2332
rect 20073 2329 20085 2332
rect 20119 2329 20131 2363
rect 20073 2323 20131 2329
rect 18472 2264 18828 2292
rect 18472 2252 18478 2264
rect 1104 2202 20884 2224
rect 1104 2150 4648 2202
rect 4700 2150 4712 2202
rect 4764 2150 4776 2202
rect 4828 2150 4840 2202
rect 4892 2150 11982 2202
rect 12034 2150 12046 2202
rect 12098 2150 12110 2202
rect 12162 2150 12174 2202
rect 12226 2150 19315 2202
rect 19367 2150 19379 2202
rect 19431 2150 19443 2202
rect 19495 2150 19507 2202
rect 19559 2150 20884 2202
rect 1104 2128 20884 2150
rect 9766 2048 9772 2100
rect 9824 2088 9830 2100
rect 15562 2088 15568 2100
rect 9824 2060 15568 2088
rect 9824 2048 9830 2060
rect 15562 2048 15568 2060
rect 15620 2048 15626 2100
rect 12342 76 12348 128
rect 12400 116 12406 128
rect 15102 116 15108 128
rect 12400 88 15108 116
rect 12400 76 12406 88
rect 15102 76 15108 88
rect 15160 76 15166 128
<< via1 >>
rect 16580 21496 16632 21548
rect 17224 21496 17276 21548
rect 4648 19558 4700 19610
rect 4712 19558 4764 19610
rect 4776 19558 4828 19610
rect 4840 19558 4892 19610
rect 11982 19558 12034 19610
rect 12046 19558 12098 19610
rect 12110 19558 12162 19610
rect 12174 19558 12226 19610
rect 19315 19558 19367 19610
rect 19379 19558 19431 19610
rect 19443 19558 19495 19610
rect 19507 19558 19559 19610
rect 8315 19014 8367 19066
rect 8379 19014 8431 19066
rect 8443 19014 8495 19066
rect 8507 19014 8559 19066
rect 15648 19014 15700 19066
rect 15712 19014 15764 19066
rect 15776 19014 15828 19066
rect 15840 19014 15892 19066
rect 4648 18470 4700 18522
rect 4712 18470 4764 18522
rect 4776 18470 4828 18522
rect 4840 18470 4892 18522
rect 11982 18470 12034 18522
rect 12046 18470 12098 18522
rect 12110 18470 12162 18522
rect 12174 18470 12226 18522
rect 19315 18470 19367 18522
rect 19379 18470 19431 18522
rect 19443 18470 19495 18522
rect 19507 18470 19559 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 4528 18368 4580 18420
rect 7656 18411 7708 18420
rect 7656 18377 7665 18411
rect 7665 18377 7699 18411
rect 7699 18377 7708 18411
rect 7656 18368 7708 18377
rect 1308 18164 1360 18216
rect 5264 18028 5316 18080
rect 10232 18028 10284 18080
rect 8315 17926 8367 17978
rect 8379 17926 8431 17978
rect 8443 17926 8495 17978
rect 8507 17926 8559 17978
rect 15648 17926 15700 17978
rect 15712 17926 15764 17978
rect 15776 17926 15828 17978
rect 15840 17926 15892 17978
rect 4648 17382 4700 17434
rect 4712 17382 4764 17434
rect 4776 17382 4828 17434
rect 4840 17382 4892 17434
rect 11982 17382 12034 17434
rect 12046 17382 12098 17434
rect 12110 17382 12162 17434
rect 12174 17382 12226 17434
rect 19315 17382 19367 17434
rect 19379 17382 19431 17434
rect 19443 17382 19495 17434
rect 19507 17382 19559 17434
rect 8315 16838 8367 16890
rect 8379 16838 8431 16890
rect 8443 16838 8495 16890
rect 8507 16838 8559 16890
rect 15648 16838 15700 16890
rect 15712 16838 15764 16890
rect 15776 16838 15828 16890
rect 15840 16838 15892 16890
rect 4648 16294 4700 16346
rect 4712 16294 4764 16346
rect 4776 16294 4828 16346
rect 4840 16294 4892 16346
rect 11982 16294 12034 16346
rect 12046 16294 12098 16346
rect 12110 16294 12162 16346
rect 12174 16294 12226 16346
rect 19315 16294 19367 16346
rect 19379 16294 19431 16346
rect 19443 16294 19495 16346
rect 19507 16294 19559 16346
rect 8315 15750 8367 15802
rect 8379 15750 8431 15802
rect 8443 15750 8495 15802
rect 8507 15750 8559 15802
rect 15648 15750 15700 15802
rect 15712 15750 15764 15802
rect 15776 15750 15828 15802
rect 15840 15750 15892 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 4648 15206 4700 15258
rect 4712 15206 4764 15258
rect 4776 15206 4828 15258
rect 4840 15206 4892 15258
rect 11982 15206 12034 15258
rect 12046 15206 12098 15258
rect 12110 15206 12162 15258
rect 12174 15206 12226 15258
rect 19315 15206 19367 15258
rect 19379 15206 19431 15258
rect 19443 15206 19495 15258
rect 19507 15206 19559 15258
rect 1400 14764 1452 14816
rect 5356 14764 5408 14816
rect 8315 14662 8367 14714
rect 8379 14662 8431 14714
rect 8443 14662 8495 14714
rect 8507 14662 8559 14714
rect 15648 14662 15700 14714
rect 15712 14662 15764 14714
rect 15776 14662 15828 14714
rect 15840 14662 15892 14714
rect 4648 14118 4700 14170
rect 4712 14118 4764 14170
rect 4776 14118 4828 14170
rect 4840 14118 4892 14170
rect 11982 14118 12034 14170
rect 12046 14118 12098 14170
rect 12110 14118 12162 14170
rect 12174 14118 12226 14170
rect 19315 14118 19367 14170
rect 19379 14118 19431 14170
rect 19443 14118 19495 14170
rect 19507 14118 19559 14170
rect 8315 13574 8367 13626
rect 8379 13574 8431 13626
rect 8443 13574 8495 13626
rect 8507 13574 8559 13626
rect 15648 13574 15700 13626
rect 15712 13574 15764 13626
rect 15776 13574 15828 13626
rect 15840 13574 15892 13626
rect 12992 13336 13044 13388
rect 13820 13336 13872 13388
rect 19064 13379 19116 13388
rect 19064 13345 19073 13379
rect 19073 13345 19107 13379
rect 19107 13345 19116 13379
rect 19064 13336 19116 13345
rect 19248 13243 19300 13252
rect 19248 13209 19257 13243
rect 19257 13209 19291 13243
rect 19291 13209 19300 13243
rect 19248 13200 19300 13209
rect 4648 13030 4700 13082
rect 4712 13030 4764 13082
rect 4776 13030 4828 13082
rect 4840 13030 4892 13082
rect 11982 13030 12034 13082
rect 12046 13030 12098 13082
rect 12110 13030 12162 13082
rect 12174 13030 12226 13082
rect 19315 13030 19367 13082
rect 19379 13030 19431 13082
rect 19443 13030 19495 13082
rect 19507 13030 19559 13082
rect 18512 12588 18564 12640
rect 19064 12631 19116 12640
rect 19064 12597 19073 12631
rect 19073 12597 19107 12631
rect 19107 12597 19116 12631
rect 19064 12588 19116 12597
rect 8315 12486 8367 12538
rect 8379 12486 8431 12538
rect 8443 12486 8495 12538
rect 8507 12486 8559 12538
rect 15648 12486 15700 12538
rect 15712 12486 15764 12538
rect 15776 12486 15828 12538
rect 15840 12486 15892 12538
rect 4648 11942 4700 11994
rect 4712 11942 4764 11994
rect 4776 11942 4828 11994
rect 4840 11942 4892 11994
rect 11982 11942 12034 11994
rect 12046 11942 12098 11994
rect 12110 11942 12162 11994
rect 12174 11942 12226 11994
rect 19315 11942 19367 11994
rect 19379 11942 19431 11994
rect 19443 11942 19495 11994
rect 19507 11942 19559 11994
rect 8315 11398 8367 11450
rect 8379 11398 8431 11450
rect 8443 11398 8495 11450
rect 8507 11398 8559 11450
rect 15648 11398 15700 11450
rect 15712 11398 15764 11450
rect 15776 11398 15828 11450
rect 15840 11398 15892 11450
rect 19340 11296 19392 11348
rect 9772 11160 9824 11212
rect 19064 11203 19116 11212
rect 19064 11169 19073 11203
rect 19073 11169 19107 11203
rect 19107 11169 19116 11203
rect 19064 11160 19116 11169
rect 8116 11092 8168 11144
rect 6920 10999 6972 11008
rect 6920 10965 6929 10999
rect 6929 10965 6963 10999
rect 6963 10965 6972 10999
rect 6920 10956 6972 10965
rect 9680 10956 9732 11008
rect 4648 10854 4700 10906
rect 4712 10854 4764 10906
rect 4776 10854 4828 10906
rect 4840 10854 4892 10906
rect 11982 10854 12034 10906
rect 12046 10854 12098 10906
rect 12110 10854 12162 10906
rect 12174 10854 12226 10906
rect 19315 10854 19367 10906
rect 19379 10854 19431 10906
rect 19443 10854 19495 10906
rect 19507 10854 19559 10906
rect 10324 10752 10376 10804
rect 8208 10548 8260 10600
rect 6920 10523 6972 10532
rect 6920 10489 6929 10523
rect 6929 10489 6963 10523
rect 6963 10489 6972 10523
rect 6920 10480 6972 10489
rect 7564 10523 7616 10532
rect 6000 10412 6052 10464
rect 7564 10489 7573 10523
rect 7573 10489 7607 10523
rect 7607 10489 7616 10523
rect 7564 10480 7616 10489
rect 7748 10480 7800 10532
rect 9588 10548 9640 10600
rect 10876 10548 10928 10600
rect 9772 10455 9824 10464
rect 9772 10421 9781 10455
rect 9781 10421 9815 10455
rect 9815 10421 9824 10455
rect 9772 10412 9824 10421
rect 10784 10412 10836 10464
rect 11336 10412 11388 10464
rect 12716 10412 12768 10464
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 15384 10412 15436 10464
rect 19064 10455 19116 10464
rect 19064 10421 19073 10455
rect 19073 10421 19107 10455
rect 19107 10421 19116 10455
rect 19064 10412 19116 10421
rect 8315 10310 8367 10362
rect 8379 10310 8431 10362
rect 8443 10310 8495 10362
rect 8507 10310 8559 10362
rect 15648 10310 15700 10362
rect 15712 10310 15764 10362
rect 15776 10310 15828 10362
rect 15840 10310 15892 10362
rect 7564 10251 7616 10260
rect 6552 10140 6604 10192
rect 7564 10217 7573 10251
rect 7573 10217 7607 10251
rect 7607 10217 7616 10251
rect 7564 10208 7616 10217
rect 8116 10183 8168 10192
rect 8116 10149 8125 10183
rect 8125 10149 8159 10183
rect 8159 10149 8168 10183
rect 8116 10140 8168 10149
rect 8208 10183 8260 10192
rect 8208 10149 8217 10183
rect 8217 10149 8251 10183
rect 8251 10149 8260 10183
rect 9772 10183 9824 10192
rect 8208 10140 8260 10149
rect 9772 10149 9781 10183
rect 9781 10149 9815 10183
rect 9815 10149 9824 10183
rect 9772 10140 9824 10149
rect 10140 10140 10192 10192
rect 12348 10115 12400 10124
rect 12348 10081 12357 10115
rect 12357 10081 12391 10115
rect 12391 10081 12400 10115
rect 12348 10072 12400 10081
rect 6368 10004 6420 10056
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 9588 10004 9640 10056
rect 6276 9936 6328 9988
rect 9772 10004 9824 10056
rect 9220 9911 9272 9920
rect 9220 9877 9229 9911
rect 9229 9877 9263 9911
rect 9263 9877 9272 9911
rect 13544 10004 13596 10056
rect 10784 9936 10836 9988
rect 13728 9936 13780 9988
rect 12440 9911 12492 9920
rect 9220 9868 9272 9877
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 4648 9766 4700 9818
rect 4712 9766 4764 9818
rect 4776 9766 4828 9818
rect 4840 9766 4892 9818
rect 11982 9766 12034 9818
rect 12046 9766 12098 9818
rect 12110 9766 12162 9818
rect 12174 9766 12226 9818
rect 19315 9766 19367 9818
rect 19379 9766 19431 9818
rect 19443 9766 19495 9818
rect 19507 9766 19559 9818
rect 6368 9664 6420 9716
rect 8208 9664 8260 9716
rect 9772 9664 9824 9716
rect 12348 9664 12400 9716
rect 16580 9664 16632 9716
rect 5264 9639 5316 9648
rect 5264 9605 5273 9639
rect 5273 9605 5307 9639
rect 5307 9605 5316 9639
rect 5264 9596 5316 9605
rect 6920 9596 6972 9648
rect 7564 9596 7616 9648
rect 21548 9596 21600 9648
rect 8392 9528 8444 9580
rect 9220 9571 9272 9580
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 12716 9528 12768 9580
rect 13728 9528 13780 9580
rect 17776 9528 17828 9580
rect 19708 9528 19760 9580
rect 5356 9460 5408 9512
rect 10968 9503 11020 9512
rect 10968 9469 10977 9503
rect 10977 9469 11011 9503
rect 11011 9469 11020 9503
rect 10968 9460 11020 9469
rect 11796 9460 11848 9512
rect 7748 9435 7800 9444
rect 7748 9401 7757 9435
rect 7757 9401 7791 9435
rect 7791 9401 7800 9435
rect 7748 9392 7800 9401
rect 9312 9435 9364 9444
rect 9312 9401 9321 9435
rect 9321 9401 9355 9435
rect 9355 9401 9364 9435
rect 9864 9435 9916 9444
rect 9312 9392 9364 9401
rect 9864 9401 9873 9435
rect 9873 9401 9907 9435
rect 9907 9401 9916 9435
rect 9864 9392 9916 9401
rect 11428 9392 11480 9444
rect 12624 9435 12676 9444
rect 12624 9401 12633 9435
rect 12633 9401 12667 9435
rect 12667 9401 12676 9435
rect 12624 9392 12676 9401
rect 13176 9435 13228 9444
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 13176 9392 13228 9401
rect 6368 9324 6420 9376
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 11152 9324 11204 9376
rect 12900 9324 12952 9376
rect 17868 9460 17920 9512
rect 18512 9503 18564 9512
rect 18512 9469 18521 9503
rect 18521 9469 18555 9503
rect 18555 9469 18564 9503
rect 18512 9460 18564 9469
rect 19248 9460 19300 9512
rect 17776 9392 17828 9444
rect 15200 9324 15252 9376
rect 15936 9324 15988 9376
rect 17224 9324 17276 9376
rect 18328 9324 18380 9376
rect 8315 9222 8367 9274
rect 8379 9222 8431 9274
rect 8443 9222 8495 9274
rect 8507 9222 8559 9274
rect 15648 9222 15700 9274
rect 15712 9222 15764 9274
rect 15776 9222 15828 9274
rect 15840 9222 15892 9274
rect 7288 9163 7340 9172
rect 7288 9129 7297 9163
rect 7297 9129 7331 9163
rect 7331 9129 7340 9163
rect 7288 9120 7340 9129
rect 7748 9120 7800 9172
rect 8116 9163 8168 9172
rect 8116 9129 8125 9163
rect 8125 9129 8159 9163
rect 8159 9129 8168 9163
rect 8116 9120 8168 9129
rect 9680 9120 9732 9172
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 18328 9120 18380 9172
rect 19156 9120 19208 9172
rect 6552 9052 6604 9104
rect 10048 9052 10100 9104
rect 1308 8984 1360 9036
rect 6000 9027 6052 9036
rect 6000 8993 6009 9027
rect 6009 8993 6043 9027
rect 6043 8993 6052 9027
rect 6000 8984 6052 8993
rect 9496 8984 9548 9036
rect 12624 9052 12676 9104
rect 13452 9052 13504 9104
rect 15936 9052 15988 9104
rect 16304 9052 16356 9104
rect 16580 9095 16632 9104
rect 16580 9061 16589 9095
rect 16589 9061 16623 9095
rect 16623 9061 16632 9095
rect 16580 9052 16632 9061
rect 6276 8848 6328 8900
rect 11060 8916 11112 8968
rect 8116 8848 8168 8900
rect 10600 8848 10652 8900
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 6460 8780 6512 8789
rect 6828 8823 6880 8832
rect 6828 8789 6837 8823
rect 6837 8789 6871 8823
rect 6871 8789 6880 8823
rect 6828 8780 6880 8789
rect 7932 8780 7984 8832
rect 9220 8823 9272 8832
rect 9220 8789 9229 8823
rect 9229 8789 9263 8823
rect 9263 8789 9272 8823
rect 9220 8780 9272 8789
rect 9956 8780 10008 8832
rect 10508 8823 10560 8832
rect 10508 8789 10517 8823
rect 10517 8789 10551 8823
rect 10551 8789 10560 8823
rect 10508 8780 10560 8789
rect 15108 8984 15160 9036
rect 17868 8984 17920 9036
rect 19156 8984 19208 9036
rect 11336 8916 11388 8968
rect 18420 8916 18472 8968
rect 13544 8891 13596 8900
rect 13544 8857 13553 8891
rect 13553 8857 13587 8891
rect 13587 8857 13596 8891
rect 13544 8848 13596 8857
rect 15384 8780 15436 8832
rect 16212 8780 16264 8832
rect 16488 8780 16540 8832
rect 4648 8678 4700 8730
rect 4712 8678 4764 8730
rect 4776 8678 4828 8730
rect 4840 8678 4892 8730
rect 11982 8678 12034 8730
rect 12046 8678 12098 8730
rect 12110 8678 12162 8730
rect 12174 8678 12226 8730
rect 19315 8678 19367 8730
rect 19379 8678 19431 8730
rect 19443 8678 19495 8730
rect 19507 8678 19559 8730
rect 1308 8576 1360 8628
rect 6000 8576 6052 8628
rect 13452 8619 13504 8628
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 15108 8576 15160 8628
rect 16212 8576 16264 8628
rect 3884 8508 3936 8560
rect 4160 8508 4212 8560
rect 9220 8508 9272 8560
rect 11428 8508 11480 8560
rect 2044 8440 2096 8492
rect 9496 8440 9548 8492
rect 9680 8483 9732 8492
rect 9680 8449 9689 8483
rect 9689 8449 9723 8483
rect 9723 8449 9732 8483
rect 9680 8440 9732 8449
rect 13176 8440 13228 8492
rect 16488 8483 16540 8492
rect 16488 8449 16497 8483
rect 16497 8449 16531 8483
rect 16531 8449 16540 8483
rect 16488 8440 16540 8449
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 18420 8440 18472 8449
rect 4528 8372 4580 8424
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 9036 8415 9088 8424
rect 9036 8381 9045 8415
rect 9045 8381 9079 8415
rect 9079 8381 9088 8415
rect 9036 8372 9088 8381
rect 10876 8372 10928 8424
rect 18880 8372 18932 8424
rect 5080 8347 5132 8356
rect 5080 8313 5089 8347
rect 5089 8313 5123 8347
rect 5123 8313 5132 8347
rect 5080 8304 5132 8313
rect 7288 8304 7340 8356
rect 8024 8347 8076 8356
rect 8024 8313 8033 8347
rect 8033 8313 8067 8347
rect 8067 8313 8076 8347
rect 8024 8304 8076 8313
rect 9772 8347 9824 8356
rect 9772 8313 9781 8347
rect 9781 8313 9815 8347
rect 9815 8313 9824 8347
rect 9772 8304 9824 8313
rect 10140 8304 10192 8356
rect 12624 8347 12676 8356
rect 12624 8313 12633 8347
rect 12633 8313 12667 8347
rect 12667 8313 12676 8347
rect 14096 8347 14148 8356
rect 12624 8304 12676 8313
rect 14096 8313 14105 8347
rect 14105 8313 14139 8347
rect 14139 8313 14148 8347
rect 14096 8304 14148 8313
rect 3976 8236 4028 8288
rect 6644 8279 6696 8288
rect 6644 8245 6653 8279
rect 6653 8245 6687 8279
rect 6687 8245 6696 8279
rect 6644 8236 6696 8245
rect 8668 8236 8720 8288
rect 11060 8279 11112 8288
rect 11060 8245 11069 8279
rect 11069 8245 11103 8279
rect 11103 8245 11112 8279
rect 11060 8236 11112 8245
rect 11612 8236 11664 8288
rect 13912 8279 13964 8288
rect 13912 8245 13921 8279
rect 13921 8245 13955 8279
rect 13955 8245 13964 8279
rect 16948 8304 17000 8356
rect 17408 8304 17460 8356
rect 17868 8347 17920 8356
rect 17868 8313 17877 8347
rect 17877 8313 17911 8347
rect 17911 8313 17920 8347
rect 17868 8304 17920 8313
rect 18236 8347 18288 8356
rect 18236 8313 18245 8347
rect 18245 8313 18279 8347
rect 18279 8313 18288 8347
rect 18236 8304 18288 8313
rect 21456 8304 21508 8356
rect 15936 8279 15988 8288
rect 13912 8236 13964 8245
rect 15936 8245 15945 8279
rect 15945 8245 15979 8279
rect 15979 8245 15988 8279
rect 15936 8236 15988 8245
rect 19156 8279 19208 8288
rect 19156 8245 19165 8279
rect 19165 8245 19199 8279
rect 19199 8245 19208 8279
rect 19156 8236 19208 8245
rect 8315 8134 8367 8186
rect 8379 8134 8431 8186
rect 8443 8134 8495 8186
rect 8507 8134 8559 8186
rect 15648 8134 15700 8186
rect 15712 8134 15764 8186
rect 15776 8134 15828 8186
rect 15840 8134 15892 8186
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 9772 8032 9824 8084
rect 10048 8075 10100 8084
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 15936 8032 15988 8084
rect 6644 7964 6696 8016
rect 5264 7828 5316 7880
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 5540 7828 5592 7837
rect 5172 7692 5224 7744
rect 5356 7692 5408 7744
rect 8024 7964 8076 8016
rect 11612 7964 11664 8016
rect 7932 7896 7984 7948
rect 13912 7964 13964 8016
rect 16028 7964 16080 8016
rect 16304 8032 16356 8084
rect 16948 8032 17000 8084
rect 18236 8032 18288 8084
rect 16580 7964 16632 8016
rect 17316 7964 17368 8016
rect 18604 7939 18656 7948
rect 18604 7905 18613 7939
rect 18613 7905 18647 7939
rect 18647 7905 18656 7939
rect 18604 7896 18656 7905
rect 9772 7828 9824 7880
rect 11520 7828 11572 7880
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 13544 7828 13596 7880
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 17224 7828 17276 7880
rect 17408 7871 17460 7880
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 17408 7828 17460 7837
rect 18788 7828 18840 7880
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 12624 7760 12676 7812
rect 7196 7692 7248 7744
rect 8208 7692 8260 7744
rect 8668 7692 8720 7744
rect 9404 7735 9456 7744
rect 9404 7701 9413 7735
rect 9413 7701 9447 7735
rect 9447 7701 9456 7735
rect 9404 7692 9456 7701
rect 11520 7735 11572 7744
rect 11520 7701 11529 7735
rect 11529 7701 11563 7735
rect 11563 7701 11572 7735
rect 11520 7692 11572 7701
rect 12348 7692 12400 7744
rect 13636 7692 13688 7744
rect 15108 7692 15160 7744
rect 16488 7735 16540 7744
rect 16488 7701 16497 7735
rect 16497 7701 16531 7735
rect 16531 7701 16540 7735
rect 16488 7692 16540 7701
rect 18144 7692 18196 7744
rect 4648 7590 4700 7642
rect 4712 7590 4764 7642
rect 4776 7590 4828 7642
rect 4840 7590 4892 7642
rect 11982 7590 12034 7642
rect 12046 7590 12098 7642
rect 12110 7590 12162 7642
rect 12174 7590 12226 7642
rect 19315 7590 19367 7642
rect 19379 7590 19431 7642
rect 19443 7590 19495 7642
rect 19507 7590 19559 7642
rect 1676 7463 1728 7472
rect 1676 7429 1685 7463
rect 1685 7429 1719 7463
rect 1719 7429 1728 7463
rect 9312 7488 9364 7540
rect 12992 7531 13044 7540
rect 12992 7497 13001 7531
rect 13001 7497 13035 7531
rect 13035 7497 13044 7531
rect 12992 7488 13044 7497
rect 13636 7531 13688 7540
rect 13636 7497 13645 7531
rect 13645 7497 13679 7531
rect 13679 7497 13688 7531
rect 13636 7488 13688 7497
rect 16948 7488 17000 7540
rect 17316 7531 17368 7540
rect 17316 7497 17325 7531
rect 17325 7497 17359 7531
rect 17359 7497 17368 7531
rect 17316 7488 17368 7497
rect 17500 7488 17552 7540
rect 1676 7420 1728 7429
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 8484 7420 8536 7472
rect 9128 7420 9180 7472
rect 10876 7420 10928 7472
rect 9864 7352 9916 7404
rect 16488 7352 16540 7404
rect 17776 7395 17828 7404
rect 17776 7361 17785 7395
rect 17785 7361 17819 7395
rect 17819 7361 17828 7395
rect 17776 7352 17828 7361
rect 3700 7327 3752 7336
rect 3700 7293 3709 7327
rect 3709 7293 3743 7327
rect 3743 7293 3752 7327
rect 3700 7284 3752 7293
rect 7472 7327 7524 7336
rect 7472 7293 7481 7327
rect 7481 7293 7515 7327
rect 7515 7293 7524 7327
rect 7472 7284 7524 7293
rect 8208 7327 8260 7336
rect 8208 7293 8217 7327
rect 8217 7293 8251 7327
rect 8251 7293 8260 7327
rect 8208 7284 8260 7293
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 8760 7284 8812 7336
rect 9956 7284 10008 7336
rect 11612 7327 11664 7336
rect 5356 7259 5408 7268
rect 5356 7225 5365 7259
rect 5365 7225 5399 7259
rect 5399 7225 5408 7259
rect 5356 7216 5408 7225
rect 7196 7216 7248 7268
rect 10048 7216 10100 7268
rect 11612 7293 11621 7327
rect 11621 7293 11655 7327
rect 11655 7293 11664 7327
rect 11612 7284 11664 7293
rect 13452 7284 13504 7336
rect 13636 7284 13688 7336
rect 14004 7284 14056 7336
rect 2044 7191 2096 7200
rect 2044 7157 2053 7191
rect 2053 7157 2087 7191
rect 2087 7157 2096 7191
rect 2044 7148 2096 7157
rect 2412 7191 2464 7200
rect 2412 7157 2421 7191
rect 2421 7157 2455 7191
rect 2455 7157 2464 7191
rect 2412 7148 2464 7157
rect 2688 7191 2740 7200
rect 2688 7157 2697 7191
rect 2697 7157 2731 7191
rect 2731 7157 2740 7191
rect 2688 7148 2740 7157
rect 3056 7191 3108 7200
rect 3056 7157 3065 7191
rect 3065 7157 3099 7191
rect 3099 7157 3108 7191
rect 3056 7148 3108 7157
rect 6092 7148 6144 7200
rect 7472 7148 7524 7200
rect 7932 7148 7984 7200
rect 10876 7148 10928 7200
rect 14648 7327 14700 7336
rect 14648 7293 14657 7327
rect 14657 7293 14691 7327
rect 14691 7293 14700 7327
rect 14648 7284 14700 7293
rect 15108 7284 15160 7336
rect 16212 7284 16264 7336
rect 12716 7148 12768 7200
rect 18604 7216 18656 7268
rect 19800 7216 19852 7268
rect 16028 7191 16080 7200
rect 16028 7157 16037 7191
rect 16037 7157 16071 7191
rect 16071 7157 16080 7191
rect 16028 7148 16080 7157
rect 18972 7148 19024 7200
rect 8315 7046 8367 7098
rect 8379 7046 8431 7098
rect 8443 7046 8495 7098
rect 8507 7046 8559 7098
rect 15648 7046 15700 7098
rect 15712 7046 15764 7098
rect 15776 7046 15828 7098
rect 15840 7046 15892 7098
rect 5540 6944 5592 6996
rect 9772 6987 9824 6996
rect 9772 6953 9781 6987
rect 9781 6953 9815 6987
rect 9815 6953 9824 6987
rect 9772 6944 9824 6953
rect 11520 6944 11572 6996
rect 13452 6944 13504 6996
rect 15292 6944 15344 6996
rect 17224 6944 17276 6996
rect 8760 6919 8812 6928
rect 1676 6808 1728 6860
rect 5264 6851 5316 6860
rect 5264 6817 5273 6851
rect 5273 6817 5307 6851
rect 5307 6817 5316 6851
rect 5264 6808 5316 6817
rect 5724 6851 5776 6860
rect 5724 6817 5733 6851
rect 5733 6817 5767 6851
rect 5767 6817 5776 6851
rect 5724 6808 5776 6817
rect 6000 6851 6052 6860
rect 6000 6817 6009 6851
rect 6009 6817 6043 6851
rect 6043 6817 6052 6851
rect 6000 6808 6052 6817
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 7932 6851 7984 6860
rect 7932 6817 7941 6851
rect 7941 6817 7975 6851
rect 7975 6817 7984 6851
rect 7932 6808 7984 6817
rect 8760 6885 8769 6919
rect 8769 6885 8803 6919
rect 8803 6885 8812 6919
rect 8760 6876 8812 6885
rect 8024 6740 8076 6792
rect 4528 6672 4580 6724
rect 6736 6672 6788 6724
rect 7840 6672 7892 6724
rect 8668 6808 8720 6860
rect 9036 6808 9088 6860
rect 17776 6919 17828 6928
rect 17776 6885 17785 6919
rect 17785 6885 17819 6919
rect 17819 6885 17828 6919
rect 17776 6876 17828 6885
rect 18420 6876 18472 6928
rect 10416 6851 10468 6860
rect 10416 6817 10425 6851
rect 10425 6817 10459 6851
rect 10459 6817 10468 6851
rect 10416 6808 10468 6817
rect 10692 6851 10744 6860
rect 10692 6817 10701 6851
rect 10701 6817 10735 6851
rect 10735 6817 10744 6851
rect 10692 6808 10744 6817
rect 10876 6851 10928 6860
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 11888 6851 11940 6860
rect 11888 6817 11897 6851
rect 11897 6817 11931 6851
rect 11931 6817 11940 6851
rect 11888 6808 11940 6817
rect 12348 6808 12400 6860
rect 12716 6851 12768 6860
rect 12716 6817 12725 6851
rect 12725 6817 12759 6851
rect 12759 6817 12768 6851
rect 12716 6808 12768 6817
rect 12900 6851 12952 6860
rect 12900 6817 12909 6851
rect 12909 6817 12943 6851
rect 12943 6817 12952 6851
rect 12900 6808 12952 6817
rect 11244 6740 11296 6792
rect 14648 6808 14700 6860
rect 15476 6851 15528 6860
rect 15476 6817 15485 6851
rect 15485 6817 15519 6851
rect 15519 6817 15528 6851
rect 15476 6808 15528 6817
rect 15752 6851 15804 6860
rect 15752 6817 15761 6851
rect 15761 6817 15795 6851
rect 15795 6817 15804 6851
rect 15752 6808 15804 6817
rect 15936 6808 15988 6860
rect 16212 6808 16264 6860
rect 19064 6808 19116 6860
rect 18144 6740 18196 6792
rect 18604 6672 18656 6724
rect 112 6604 164 6656
rect 2136 6647 2188 6656
rect 2136 6613 2145 6647
rect 2145 6613 2179 6647
rect 2179 6613 2188 6647
rect 2136 6604 2188 6613
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 2780 6604 2832 6656
rect 3608 6647 3660 6656
rect 3608 6613 3617 6647
rect 3617 6613 3651 6647
rect 3651 6613 3660 6647
rect 3608 6604 3660 6613
rect 4988 6604 5040 6656
rect 6920 6604 6972 6656
rect 16212 6604 16264 6656
rect 18696 6647 18748 6656
rect 18696 6613 18705 6647
rect 18705 6613 18739 6647
rect 18739 6613 18748 6647
rect 18696 6604 18748 6613
rect 4648 6502 4700 6554
rect 4712 6502 4764 6554
rect 4776 6502 4828 6554
rect 4840 6502 4892 6554
rect 11982 6502 12034 6554
rect 12046 6502 12098 6554
rect 12110 6502 12162 6554
rect 12174 6502 12226 6554
rect 19315 6502 19367 6554
rect 19379 6502 19431 6554
rect 19443 6502 19495 6554
rect 19507 6502 19559 6554
rect 1860 6400 1912 6452
rect 6736 6400 6788 6452
rect 10508 6400 10560 6452
rect 15752 6400 15804 6452
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 18696 6400 18748 6452
rect 7104 6375 7156 6384
rect 7104 6341 7113 6375
rect 7113 6341 7147 6375
rect 7147 6341 7156 6375
rect 7104 6332 7156 6341
rect 7472 6332 7524 6384
rect 6552 6264 6604 6316
rect 9220 6264 9272 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 2320 6239 2372 6248
rect 2320 6205 2329 6239
rect 2329 6205 2363 6239
rect 2363 6205 2372 6239
rect 2320 6196 2372 6205
rect 4436 6196 4488 6248
rect 5356 6239 5408 6248
rect 5356 6205 5365 6239
rect 5365 6205 5399 6239
rect 5399 6205 5408 6239
rect 5356 6196 5408 6205
rect 6920 6196 6972 6248
rect 4344 6171 4396 6180
rect 4344 6137 4353 6171
rect 4353 6137 4387 6171
rect 4387 6137 4396 6171
rect 4344 6128 4396 6137
rect 5724 6128 5776 6180
rect 7932 6196 7984 6248
rect 11060 6332 11112 6384
rect 11980 6264 12032 6316
rect 12716 6264 12768 6316
rect 10416 6196 10468 6248
rect 11244 6239 11296 6248
rect 7564 6171 7616 6180
rect 7564 6137 7573 6171
rect 7573 6137 7607 6171
rect 7607 6137 7616 6171
rect 7564 6128 7616 6137
rect 8760 6128 8812 6180
rect 9220 6171 9272 6180
rect 9220 6137 9229 6171
rect 9229 6137 9263 6171
rect 9263 6137 9272 6171
rect 9220 6128 9272 6137
rect 11244 6205 11253 6239
rect 11253 6205 11287 6239
rect 11287 6205 11296 6239
rect 11244 6196 11296 6205
rect 11796 6196 11848 6248
rect 14004 6239 14056 6248
rect 14004 6205 14013 6239
rect 14013 6205 14047 6239
rect 14047 6205 14056 6239
rect 14004 6196 14056 6205
rect 16212 6307 16264 6316
rect 16212 6273 16221 6307
rect 16221 6273 16255 6307
rect 16255 6273 16264 6307
rect 16212 6264 16264 6273
rect 18788 6307 18840 6316
rect 18788 6273 18797 6307
rect 18797 6273 18831 6307
rect 18831 6273 18840 6307
rect 18788 6264 18840 6273
rect 15108 6239 15160 6248
rect 1768 6060 1820 6112
rect 2412 6060 2464 6112
rect 5264 6060 5316 6112
rect 5816 6060 5868 6112
rect 6000 6060 6052 6112
rect 6368 6060 6420 6112
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 6552 6060 6604 6069
rect 7840 6103 7892 6112
rect 7840 6069 7849 6103
rect 7849 6069 7883 6103
rect 7883 6069 7892 6103
rect 7840 6060 7892 6069
rect 7932 6060 7984 6112
rect 9312 6060 9364 6112
rect 9772 6060 9824 6112
rect 10048 6060 10100 6112
rect 11244 6060 11296 6112
rect 11612 6060 11664 6112
rect 12900 6060 12952 6112
rect 15108 6205 15117 6239
rect 15117 6205 15151 6239
rect 15151 6205 15160 6239
rect 15108 6196 15160 6205
rect 19708 6239 19760 6248
rect 19708 6205 19726 6239
rect 19726 6205 19760 6239
rect 19708 6196 19760 6205
rect 16120 6128 16172 6180
rect 17776 6128 17828 6180
rect 15936 6060 15988 6112
rect 16212 6060 16264 6112
rect 19064 6060 19116 6112
rect 8315 5958 8367 6010
rect 8379 5958 8431 6010
rect 8443 5958 8495 6010
rect 8507 5958 8559 6010
rect 15648 5958 15700 6010
rect 15712 5958 15764 6010
rect 15776 5958 15828 6010
rect 15840 5958 15892 6010
rect 6828 5899 6880 5908
rect 6828 5865 6837 5899
rect 6837 5865 6871 5899
rect 6871 5865 6880 5899
rect 6828 5856 6880 5865
rect 2964 5788 3016 5840
rect 1860 5720 1912 5772
rect 2136 5720 2188 5772
rect 3332 5652 3384 5704
rect 4988 5720 5040 5772
rect 7012 5788 7064 5840
rect 8116 5831 8168 5840
rect 8116 5797 8125 5831
rect 8125 5797 8159 5831
rect 8159 5797 8168 5831
rect 8116 5788 8168 5797
rect 8852 5856 8904 5908
rect 9128 5899 9180 5908
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 10692 5856 10744 5908
rect 11704 5899 11756 5908
rect 8760 5788 8812 5840
rect 9404 5788 9456 5840
rect 10876 5788 10928 5840
rect 11704 5865 11713 5899
rect 11713 5865 11747 5899
rect 11747 5865 11756 5899
rect 11704 5856 11756 5865
rect 12532 5856 12584 5908
rect 14648 5856 14700 5908
rect 15108 5899 15160 5908
rect 15108 5865 15117 5899
rect 15117 5865 15151 5899
rect 15151 5865 15160 5899
rect 15108 5856 15160 5865
rect 15476 5899 15528 5908
rect 15476 5865 15485 5899
rect 15485 5865 15519 5899
rect 15519 5865 15528 5899
rect 15476 5856 15528 5865
rect 17408 5856 17460 5908
rect 11796 5788 11848 5840
rect 12348 5788 12400 5840
rect 14004 5831 14056 5840
rect 14004 5797 14013 5831
rect 14013 5797 14047 5831
rect 14047 5797 14056 5831
rect 14004 5788 14056 5797
rect 16120 5788 16172 5840
rect 18144 5856 18196 5908
rect 18788 5899 18840 5908
rect 18788 5865 18797 5899
rect 18797 5865 18831 5899
rect 18831 5865 18840 5899
rect 18788 5856 18840 5865
rect 4528 5652 4580 5704
rect 6644 5652 6696 5704
rect 4068 5584 4120 5636
rect 5356 5584 5408 5636
rect 6000 5584 6052 5636
rect 7840 5720 7892 5772
rect 11888 5763 11940 5772
rect 11888 5729 11897 5763
rect 11897 5729 11931 5763
rect 11931 5729 11940 5763
rect 11888 5720 11940 5729
rect 11980 5720 12032 5772
rect 12532 5763 12584 5772
rect 12532 5729 12541 5763
rect 12541 5729 12575 5763
rect 12575 5729 12584 5763
rect 12532 5720 12584 5729
rect 12808 5763 12860 5772
rect 12808 5729 12817 5763
rect 12817 5729 12851 5763
rect 12851 5729 12860 5763
rect 12808 5720 12860 5729
rect 13176 5720 13228 5772
rect 18880 5720 18932 5772
rect 19064 5763 19116 5772
rect 19064 5729 19073 5763
rect 19073 5729 19107 5763
rect 19107 5729 19116 5763
rect 19064 5720 19116 5729
rect 10508 5652 10560 5704
rect 7196 5584 7248 5636
rect 12624 5652 12676 5704
rect 13728 5695 13780 5704
rect 13728 5661 13737 5695
rect 13737 5661 13771 5695
rect 13771 5661 13780 5695
rect 13728 5652 13780 5661
rect 15476 5652 15528 5704
rect 15660 5695 15712 5704
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 18420 5652 18472 5704
rect 18512 5652 18564 5704
rect 15936 5584 15988 5636
rect 1860 5516 1912 5568
rect 2412 5559 2464 5568
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 3516 5559 3568 5568
rect 3516 5525 3525 5559
rect 3525 5525 3559 5559
rect 3559 5525 3568 5559
rect 3516 5516 3568 5525
rect 3884 5516 3936 5568
rect 4436 5516 4488 5568
rect 7288 5516 7340 5568
rect 7472 5559 7524 5568
rect 7472 5525 7481 5559
rect 7481 5525 7515 5559
rect 7515 5525 7524 5559
rect 7472 5516 7524 5525
rect 9404 5559 9456 5568
rect 9404 5525 9413 5559
rect 9413 5525 9447 5559
rect 9447 5525 9456 5559
rect 9404 5516 9456 5525
rect 10416 5516 10468 5568
rect 10968 5516 11020 5568
rect 11060 5516 11112 5568
rect 12808 5516 12860 5568
rect 4648 5414 4700 5466
rect 4712 5414 4764 5466
rect 4776 5414 4828 5466
rect 4840 5414 4892 5466
rect 11982 5414 12034 5466
rect 12046 5414 12098 5466
rect 12110 5414 12162 5466
rect 12174 5414 12226 5466
rect 19315 5414 19367 5466
rect 19379 5414 19431 5466
rect 19443 5414 19495 5466
rect 19507 5414 19559 5466
rect 2228 5312 2280 5364
rect 4252 5312 4304 5364
rect 4344 5312 4396 5364
rect 6920 5312 6972 5364
rect 8760 5312 8812 5364
rect 10784 5312 10836 5364
rect 4528 5244 4580 5296
rect 5540 5244 5592 5296
rect 5816 5244 5868 5296
rect 7472 5244 7524 5296
rect 7840 5244 7892 5296
rect 5632 5176 5684 5228
rect 6184 5176 6236 5228
rect 8668 5244 8720 5296
rect 9128 5244 9180 5296
rect 8760 5176 8812 5228
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 3332 5040 3384 5092
rect 3516 5108 3568 5160
rect 7840 5108 7892 5160
rect 8024 5108 8076 5160
rect 8208 5151 8260 5160
rect 8208 5117 8217 5151
rect 8217 5117 8251 5151
rect 8251 5117 8260 5151
rect 9036 5151 9088 5160
rect 8208 5108 8260 5117
rect 3608 5040 3660 5092
rect 3700 5040 3752 5092
rect 4988 5083 5040 5092
rect 2964 5015 3016 5024
rect 2964 4981 2973 5015
rect 2973 4981 3007 5015
rect 3007 4981 3016 5015
rect 2964 4972 3016 4981
rect 3516 5015 3568 5024
rect 3516 4981 3525 5015
rect 3525 4981 3559 5015
rect 3559 4981 3568 5015
rect 3516 4972 3568 4981
rect 3884 4972 3936 5024
rect 4436 5015 4488 5024
rect 4436 4981 4445 5015
rect 4445 4981 4479 5015
rect 4479 4981 4488 5015
rect 4436 4972 4488 4981
rect 4988 5049 4997 5083
rect 4997 5049 5031 5083
rect 5031 5049 5040 5083
rect 4988 5040 5040 5049
rect 7104 5040 7156 5092
rect 7196 5040 7248 5092
rect 9036 5117 9045 5151
rect 9045 5117 9079 5151
rect 9079 5117 9088 5151
rect 9036 5108 9088 5117
rect 9404 5108 9456 5160
rect 9772 5108 9824 5160
rect 10140 5151 10192 5160
rect 10140 5117 10149 5151
rect 10149 5117 10183 5151
rect 10183 5117 10192 5151
rect 10140 5108 10192 5117
rect 10968 5312 11020 5364
rect 11888 5244 11940 5296
rect 12992 5312 13044 5364
rect 17408 5355 17460 5364
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 18420 5312 18472 5364
rect 19064 5355 19116 5364
rect 19064 5321 19073 5355
rect 19073 5321 19107 5355
rect 19107 5321 19116 5355
rect 19064 5312 19116 5321
rect 12716 5244 12768 5296
rect 18880 5244 18932 5296
rect 13728 5151 13780 5160
rect 13728 5117 13737 5151
rect 13737 5117 13771 5151
rect 13771 5117 13780 5151
rect 13728 5108 13780 5117
rect 15660 5176 15712 5228
rect 16764 5176 16816 5228
rect 18788 5176 18840 5228
rect 14648 5151 14700 5160
rect 14648 5117 14657 5151
rect 14657 5117 14691 5151
rect 14691 5117 14700 5151
rect 14648 5108 14700 5117
rect 15108 5151 15160 5160
rect 15108 5117 15117 5151
rect 15117 5117 15151 5151
rect 15151 5117 15160 5151
rect 15108 5108 15160 5117
rect 16028 5151 16080 5160
rect 16028 5117 16037 5151
rect 16037 5117 16071 5151
rect 16071 5117 16080 5151
rect 16028 5108 16080 5117
rect 13176 5083 13228 5092
rect 6000 5015 6052 5024
rect 6000 4981 6009 5015
rect 6009 4981 6043 5015
rect 6043 4981 6052 5015
rect 6000 4972 6052 4981
rect 6644 4972 6696 5024
rect 9036 5015 9088 5024
rect 9036 4981 9045 5015
rect 9045 4981 9079 5015
rect 9079 4981 9088 5015
rect 9036 4972 9088 4981
rect 9588 4972 9640 5024
rect 13176 5049 13185 5083
rect 13185 5049 13219 5083
rect 13219 5049 13228 5083
rect 13176 5040 13228 5049
rect 10968 4972 11020 5024
rect 11060 4972 11112 5024
rect 12900 4972 12952 5024
rect 15384 4972 15436 5024
rect 16120 4972 16172 5024
rect 19156 4972 19208 5024
rect 8315 4870 8367 4922
rect 8379 4870 8431 4922
rect 8443 4870 8495 4922
rect 8507 4870 8559 4922
rect 15648 4870 15700 4922
rect 15712 4870 15764 4922
rect 15776 4870 15828 4922
rect 15840 4870 15892 4922
rect 848 4768 900 4820
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 2228 4811 2280 4820
rect 2228 4777 2237 4811
rect 2237 4777 2271 4811
rect 2271 4777 2280 4811
rect 2228 4768 2280 4777
rect 3332 4768 3384 4820
rect 4528 4768 4580 4820
rect 5632 4811 5684 4820
rect 5632 4777 5641 4811
rect 5641 4777 5675 4811
rect 5675 4777 5684 4811
rect 5632 4768 5684 4777
rect 6460 4811 6512 4820
rect 6460 4777 6469 4811
rect 6469 4777 6503 4811
rect 6503 4777 6512 4811
rect 6460 4768 6512 4777
rect 7288 4768 7340 4820
rect 9128 4768 9180 4820
rect 10140 4768 10192 4820
rect 10876 4811 10928 4820
rect 10876 4777 10885 4811
rect 10885 4777 10919 4811
rect 10919 4777 10928 4811
rect 10876 4768 10928 4777
rect 2412 4700 2464 4752
rect 3056 4743 3108 4752
rect 3056 4709 3065 4743
rect 3065 4709 3099 4743
rect 3099 4709 3108 4743
rect 3056 4700 3108 4709
rect 4252 4700 4304 4752
rect 5356 4675 5408 4684
rect 5356 4641 5365 4675
rect 5365 4641 5399 4675
rect 5399 4641 5408 4675
rect 5356 4632 5408 4641
rect 2688 4564 2740 4616
rect 4160 4564 4212 4616
rect 6920 4700 6972 4752
rect 5724 4632 5776 4684
rect 6644 4675 6696 4684
rect 6644 4641 6653 4675
rect 6653 4641 6687 4675
rect 6687 4641 6696 4675
rect 6644 4632 6696 4641
rect 7012 4675 7064 4684
rect 7012 4641 7021 4675
rect 7021 4641 7055 4675
rect 7055 4641 7064 4675
rect 7012 4632 7064 4641
rect 6000 4564 6052 4616
rect 6368 4564 6420 4616
rect 7932 4632 7984 4684
rect 8944 4632 8996 4684
rect 9220 4632 9272 4684
rect 11244 4700 11296 4752
rect 12348 4743 12400 4752
rect 12348 4709 12357 4743
rect 12357 4709 12391 4743
rect 12391 4709 12400 4743
rect 12348 4700 12400 4709
rect 11704 4632 11756 4684
rect 13084 4632 13136 4684
rect 13912 4700 13964 4752
rect 14648 4743 14700 4752
rect 13360 4675 13412 4684
rect 13360 4641 13369 4675
rect 13369 4641 13403 4675
rect 13403 4641 13412 4675
rect 13360 4632 13412 4641
rect 13728 4632 13780 4684
rect 14648 4709 14657 4743
rect 14657 4709 14691 4743
rect 14691 4709 14700 4743
rect 14648 4700 14700 4709
rect 15292 4768 15344 4820
rect 16028 4768 16080 4820
rect 14096 4632 14148 4684
rect 14924 4632 14976 4684
rect 15108 4675 15160 4684
rect 15108 4641 15117 4675
rect 15117 4641 15151 4675
rect 15151 4641 15160 4675
rect 15108 4632 15160 4641
rect 16120 4700 16172 4752
rect 16304 4700 16356 4752
rect 17408 4700 17460 4752
rect 16396 4632 16448 4684
rect 16764 4675 16816 4684
rect 16764 4641 16773 4675
rect 16773 4641 16807 4675
rect 16807 4641 16816 4675
rect 16764 4632 16816 4641
rect 19064 4675 19116 4684
rect 19064 4641 19073 4675
rect 19073 4641 19107 4675
rect 19107 4641 19116 4675
rect 19064 4632 19116 4641
rect 8116 4564 8168 4616
rect 10324 4564 10376 4616
rect 13636 4564 13688 4616
rect 16672 4564 16724 4616
rect 17408 4607 17460 4616
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 17408 4564 17460 4573
rect 17684 4607 17736 4616
rect 17684 4573 17693 4607
rect 17693 4573 17727 4607
rect 17727 4573 17736 4607
rect 17684 4564 17736 4573
rect 17776 4564 17828 4616
rect 8852 4496 8904 4548
rect 9312 4496 9364 4548
rect 11336 4496 11388 4548
rect 13360 4496 13412 4548
rect 18236 4496 18288 4548
rect 5540 4428 5592 4480
rect 8576 4428 8628 4480
rect 8944 4428 8996 4480
rect 10600 4428 10652 4480
rect 15108 4428 15160 4480
rect 4648 4326 4700 4378
rect 4712 4326 4764 4378
rect 4776 4326 4828 4378
rect 4840 4326 4892 4378
rect 11982 4326 12034 4378
rect 12046 4326 12098 4378
rect 12110 4326 12162 4378
rect 12174 4326 12226 4378
rect 19315 4326 19367 4378
rect 19379 4326 19431 4378
rect 19443 4326 19495 4378
rect 19507 4326 19559 4378
rect 2412 4224 2464 4276
rect 2964 4224 3016 4276
rect 4068 4224 4120 4276
rect 5724 4224 5776 4276
rect 4896 4156 4948 4208
rect 5816 4199 5868 4208
rect 5816 4165 5825 4199
rect 5825 4165 5859 4199
rect 5859 4165 5868 4199
rect 5816 4156 5868 4165
rect 7472 4156 7524 4208
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 5540 4131 5592 4140
rect 5540 4097 5549 4131
rect 5549 4097 5583 4131
rect 5583 4097 5592 4131
rect 5540 4088 5592 4097
rect 1860 3995 1912 4004
rect 1860 3961 1869 3995
rect 1869 3961 1903 3995
rect 1903 3961 1912 3995
rect 1860 3952 1912 3961
rect 3056 3952 3108 4004
rect 3608 3952 3660 4004
rect 3976 3995 4028 4004
rect 3976 3961 3985 3995
rect 3985 3961 4019 3995
rect 4019 3961 4028 3995
rect 3976 3952 4028 3961
rect 3884 3884 3936 3936
rect 6552 4020 6604 4072
rect 4344 3995 4396 4004
rect 4344 3961 4353 3995
rect 4353 3961 4387 3995
rect 4387 3961 4396 3995
rect 4344 3952 4396 3961
rect 6000 3952 6052 4004
rect 8208 4156 8260 4208
rect 9312 4156 9364 4208
rect 11152 4156 11204 4208
rect 11796 4199 11848 4208
rect 11796 4165 11805 4199
rect 11805 4165 11839 4199
rect 11839 4165 11848 4199
rect 11796 4156 11848 4165
rect 13084 4199 13136 4208
rect 13084 4165 13093 4199
rect 13093 4165 13127 4199
rect 13127 4165 13136 4199
rect 13084 4156 13136 4165
rect 13636 4224 13688 4276
rect 18144 4224 18196 4276
rect 18788 4224 18840 4276
rect 19064 4267 19116 4276
rect 19064 4233 19073 4267
rect 19073 4233 19107 4267
rect 19107 4233 19116 4267
rect 19064 4224 19116 4233
rect 14096 4156 14148 4208
rect 15292 4199 15344 4208
rect 15292 4165 15301 4199
rect 15301 4165 15335 4199
rect 15335 4165 15344 4199
rect 15292 4156 15344 4165
rect 15476 4156 15528 4208
rect 17408 4156 17460 4208
rect 19616 4156 19668 4208
rect 8852 4088 8904 4140
rect 12164 4131 12216 4140
rect 8576 4063 8628 4072
rect 8024 3952 8076 4004
rect 8576 4029 8585 4063
rect 8585 4029 8619 4063
rect 8619 4029 8628 4063
rect 8576 4020 8628 4029
rect 9128 4063 9180 4072
rect 9128 4029 9137 4063
rect 9137 4029 9171 4063
rect 9171 4029 9180 4063
rect 9128 4020 9180 4029
rect 9496 4020 9548 4072
rect 12164 4097 12173 4131
rect 12173 4097 12207 4131
rect 12207 4097 12216 4131
rect 12164 4088 12216 4097
rect 9036 3952 9088 4004
rect 17684 4088 17736 4140
rect 18144 4131 18196 4140
rect 18144 4097 18153 4131
rect 18153 4097 18187 4131
rect 18187 4097 18196 4131
rect 18144 4088 18196 4097
rect 18880 4088 18932 4140
rect 13912 4063 13964 4072
rect 13912 4029 13921 4063
rect 13921 4029 13955 4063
rect 13955 4029 13964 4063
rect 13912 4020 13964 4029
rect 14372 4063 14424 4072
rect 14372 4029 14381 4063
rect 14381 4029 14415 4063
rect 14415 4029 14424 4063
rect 14372 4020 14424 4029
rect 14832 4063 14884 4072
rect 14832 4029 14841 4063
rect 14841 4029 14875 4063
rect 14875 4029 14884 4063
rect 14832 4020 14884 4029
rect 14924 4020 14976 4072
rect 19616 4020 19668 4072
rect 6184 3927 6236 3936
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 6644 3884 6696 3936
rect 7840 3927 7892 3936
rect 7840 3893 7849 3927
rect 7849 3893 7883 3927
rect 7883 3893 7892 3927
rect 7840 3884 7892 3893
rect 7932 3884 7984 3936
rect 9588 3884 9640 3936
rect 9864 3927 9916 3936
rect 9864 3893 9873 3927
rect 9873 3893 9907 3927
rect 9907 3893 9916 3927
rect 12624 3952 12676 4004
rect 13544 3952 13596 4004
rect 16304 3995 16356 4004
rect 16304 3961 16313 3995
rect 16313 3961 16347 3995
rect 16347 3961 16356 3995
rect 16304 3952 16356 3961
rect 16396 3995 16448 4004
rect 16396 3961 16405 3995
rect 16405 3961 16439 3995
rect 16439 3961 16448 3995
rect 18236 3995 18288 4004
rect 16396 3952 16448 3961
rect 18236 3961 18245 3995
rect 18245 3961 18279 3995
rect 18279 3961 18288 3995
rect 18236 3952 18288 3961
rect 20168 3952 20220 4004
rect 11244 3927 11296 3936
rect 9864 3884 9916 3893
rect 11244 3893 11253 3927
rect 11253 3893 11287 3927
rect 11287 3893 11296 3927
rect 11244 3884 11296 3893
rect 11704 3884 11756 3936
rect 14832 3884 14884 3936
rect 15384 3884 15436 3936
rect 17408 3884 17460 3936
rect 8315 3782 8367 3834
rect 8379 3782 8431 3834
rect 8443 3782 8495 3834
rect 8507 3782 8559 3834
rect 15648 3782 15700 3834
rect 15712 3782 15764 3834
rect 15776 3782 15828 3834
rect 15840 3782 15892 3834
rect 1860 3680 1912 3732
rect 2964 3680 3016 3732
rect 4344 3680 4396 3732
rect 4896 3723 4948 3732
rect 4896 3689 4905 3723
rect 4905 3689 4939 3723
rect 4939 3689 4948 3723
rect 4896 3680 4948 3689
rect 2320 3655 2372 3664
rect 2320 3621 2323 3655
rect 2323 3621 2357 3655
rect 2357 3621 2372 3655
rect 2320 3612 2372 3621
rect 2780 3612 2832 3664
rect 5172 3680 5224 3732
rect 8944 3680 8996 3732
rect 13268 3680 13320 3732
rect 14004 3680 14056 3732
rect 14372 3680 14424 3732
rect 14924 3723 14976 3732
rect 14924 3689 14933 3723
rect 14933 3689 14967 3723
rect 14967 3689 14976 3723
rect 14924 3680 14976 3689
rect 16396 3723 16448 3732
rect 16396 3689 16405 3723
rect 16405 3689 16439 3723
rect 16439 3689 16448 3723
rect 16396 3680 16448 3689
rect 16672 3723 16724 3732
rect 16672 3689 16681 3723
rect 16681 3689 16715 3723
rect 16715 3689 16724 3723
rect 16672 3680 16724 3689
rect 17684 3680 17736 3732
rect 19616 3680 19668 3732
rect 5080 3544 5132 3596
rect 5264 3587 5316 3596
rect 5264 3553 5273 3587
rect 5273 3553 5307 3587
rect 5307 3553 5316 3587
rect 5264 3544 5316 3553
rect 6000 3587 6052 3596
rect 2044 3476 2096 3528
rect 4528 3476 4580 3528
rect 6000 3553 6009 3587
rect 6009 3553 6043 3587
rect 6043 3553 6052 3587
rect 6000 3544 6052 3553
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 7104 3612 7156 3664
rect 9220 3612 9272 3664
rect 10692 3612 10744 3664
rect 15016 3612 15068 3664
rect 17132 3612 17184 3664
rect 17776 3612 17828 3664
rect 18696 3612 18748 3664
rect 6920 3544 6972 3596
rect 8116 3587 8168 3596
rect 6644 3476 6696 3528
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 8760 3544 8812 3596
rect 9404 3544 9456 3596
rect 10048 3544 10100 3596
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 11336 3587 11388 3596
rect 11336 3553 11345 3587
rect 11345 3553 11379 3587
rect 11379 3553 11388 3587
rect 11336 3544 11388 3553
rect 11704 3587 11756 3596
rect 7012 3408 7064 3460
rect 7748 3408 7800 3460
rect 8208 3476 8260 3528
rect 10968 3476 11020 3528
rect 11704 3553 11713 3587
rect 11713 3553 11747 3587
rect 11747 3553 11756 3587
rect 11704 3544 11756 3553
rect 11796 3544 11848 3596
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 13084 3544 13136 3596
rect 13268 3519 13320 3528
rect 13268 3485 13277 3519
rect 13277 3485 13311 3519
rect 13311 3485 13320 3519
rect 13268 3476 13320 3485
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 15108 3476 15160 3528
rect 1768 3383 1820 3392
rect 1768 3349 1777 3383
rect 1777 3349 1811 3383
rect 1811 3349 1820 3383
rect 1768 3340 1820 3349
rect 4436 3340 4488 3392
rect 4988 3340 5040 3392
rect 9864 3340 9916 3392
rect 11152 3340 11204 3392
rect 12808 3408 12860 3460
rect 13820 3408 13872 3460
rect 15476 3476 15528 3528
rect 17684 3451 17736 3460
rect 17684 3417 17693 3451
rect 17693 3417 17727 3451
rect 17727 3417 17736 3451
rect 17684 3408 17736 3417
rect 17776 3408 17828 3460
rect 11704 3340 11756 3392
rect 17224 3340 17276 3392
rect 17316 3340 17368 3392
rect 17592 3340 17644 3392
rect 18880 3476 18932 3528
rect 4648 3238 4700 3290
rect 4712 3238 4764 3290
rect 4776 3238 4828 3290
rect 4840 3238 4892 3290
rect 11982 3238 12034 3290
rect 12046 3238 12098 3290
rect 12110 3238 12162 3290
rect 12174 3238 12226 3290
rect 19315 3238 19367 3290
rect 19379 3238 19431 3290
rect 19443 3238 19495 3290
rect 19507 3238 19559 3290
rect 1952 3136 2004 3188
rect 3608 3179 3660 3188
rect 3608 3145 3617 3179
rect 3617 3145 3651 3179
rect 3651 3145 3660 3179
rect 3608 3136 3660 3145
rect 3700 3136 3752 3188
rect 2688 3068 2740 3120
rect 6000 3136 6052 3188
rect 8760 3136 8812 3188
rect 10048 3179 10100 3188
rect 4988 3068 5040 3120
rect 6184 3111 6236 3120
rect 6184 3077 6193 3111
rect 6193 3077 6227 3111
rect 6227 3077 6236 3111
rect 6184 3068 6236 3077
rect 1952 2932 2004 2984
rect 2780 2932 2832 2984
rect 4988 2975 5040 2984
rect 2320 2796 2372 2848
rect 4620 2864 4672 2916
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 8024 3000 8076 3052
rect 10048 3145 10057 3179
rect 10057 3145 10091 3179
rect 10091 3145 10100 3179
rect 10048 3136 10100 3145
rect 10968 3136 11020 3188
rect 11336 3136 11388 3188
rect 11152 3068 11204 3120
rect 5264 2864 5316 2916
rect 6552 2932 6604 2984
rect 8208 2932 8260 2984
rect 9036 2932 9088 2984
rect 12348 3000 12400 3052
rect 9496 2975 9548 2984
rect 9496 2941 9505 2975
rect 9505 2941 9539 2975
rect 9539 2941 9548 2975
rect 9496 2932 9548 2941
rect 13268 3136 13320 3188
rect 15016 3179 15068 3188
rect 15016 3145 15025 3179
rect 15025 3145 15059 3179
rect 15059 3145 15068 3179
rect 15016 3136 15068 3145
rect 17132 3179 17184 3188
rect 17132 3145 17141 3179
rect 17141 3145 17175 3179
rect 17175 3145 17184 3179
rect 17132 3136 17184 3145
rect 17224 3136 17276 3188
rect 19156 3136 19208 3188
rect 6000 2864 6052 2916
rect 7104 2864 7156 2916
rect 9772 2907 9824 2916
rect 9772 2873 9781 2907
rect 9781 2873 9815 2907
rect 9815 2873 9824 2907
rect 9772 2864 9824 2873
rect 9864 2864 9916 2916
rect 12256 2864 12308 2916
rect 4528 2839 4580 2848
rect 4528 2805 4537 2839
rect 4537 2805 4571 2839
rect 4571 2805 4580 2839
rect 4528 2796 4580 2805
rect 13084 2932 13136 2984
rect 14004 3000 14056 3052
rect 14188 3043 14240 3052
rect 14188 3009 14197 3043
rect 14197 3009 14231 3043
rect 14231 3009 14240 3043
rect 14188 3000 14240 3009
rect 17316 3000 17368 3052
rect 17684 3000 17736 3052
rect 13728 2975 13780 2984
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13728 2932 13780 2941
rect 13820 2932 13872 2984
rect 14924 2932 14976 2984
rect 17776 2932 17828 2984
rect 18972 2932 19024 2984
rect 13360 2864 13412 2916
rect 14004 2864 14056 2916
rect 15384 2907 15436 2916
rect 15384 2873 15393 2907
rect 15393 2873 15427 2907
rect 15427 2873 15436 2907
rect 15384 2864 15436 2873
rect 17592 2864 17644 2916
rect 17868 2864 17920 2916
rect 16672 2796 16724 2848
rect 17776 2839 17828 2848
rect 17776 2805 17785 2839
rect 17785 2805 17819 2839
rect 17819 2805 17828 2839
rect 18420 2864 18472 2916
rect 18788 2907 18840 2916
rect 18788 2873 18797 2907
rect 18797 2873 18831 2907
rect 18831 2873 18840 2907
rect 18788 2864 18840 2873
rect 21548 2864 21600 2916
rect 19432 2839 19484 2848
rect 17776 2796 17828 2805
rect 19432 2805 19441 2839
rect 19441 2805 19475 2839
rect 19475 2805 19484 2839
rect 19432 2796 19484 2805
rect 8315 2694 8367 2746
rect 8379 2694 8431 2746
rect 8443 2694 8495 2746
rect 8507 2694 8559 2746
rect 15648 2694 15700 2746
rect 15712 2694 15764 2746
rect 15776 2694 15828 2746
rect 15840 2694 15892 2746
rect 1768 2592 1820 2644
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 4620 2635 4672 2644
rect 4620 2601 4629 2635
rect 4629 2601 4663 2635
rect 4663 2601 4672 2635
rect 4620 2592 4672 2601
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 3976 2456 4028 2508
rect 6184 2524 6236 2576
rect 2320 2388 2372 2440
rect 5172 2456 5224 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 7748 2499 7800 2508
rect 7748 2465 7757 2499
rect 7757 2465 7791 2499
rect 7791 2465 7800 2499
rect 7748 2456 7800 2465
rect 11520 2592 11572 2644
rect 9036 2567 9088 2576
rect 9036 2533 9045 2567
rect 9045 2533 9079 2567
rect 9079 2533 9088 2567
rect 9036 2524 9088 2533
rect 9864 2524 9916 2576
rect 10324 2524 10376 2576
rect 13636 2524 13688 2576
rect 14004 2524 14056 2576
rect 15016 2524 15068 2576
rect 17868 2592 17920 2644
rect 16672 2567 16724 2576
rect 10692 2499 10744 2508
rect 10692 2465 10701 2499
rect 10701 2465 10735 2499
rect 10735 2465 10744 2499
rect 10692 2456 10744 2465
rect 8208 2388 8260 2440
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 10140 2388 10192 2440
rect 12256 2456 12308 2508
rect 13360 2499 13412 2508
rect 13360 2465 13369 2499
rect 13369 2465 13403 2499
rect 13403 2465 13412 2499
rect 13360 2456 13412 2465
rect 14188 2456 14240 2508
rect 15384 2456 15436 2508
rect 15568 2499 15620 2508
rect 15568 2465 15586 2499
rect 15586 2465 15620 2499
rect 15568 2456 15620 2465
rect 16212 2456 16264 2508
rect 11152 2388 11204 2440
rect 11796 2388 11848 2440
rect 12348 2388 12400 2440
rect 6460 2320 6512 2372
rect 16672 2533 16681 2567
rect 16681 2533 16715 2567
rect 16715 2533 16724 2567
rect 16672 2524 16724 2533
rect 17684 2524 17736 2576
rect 18512 2567 18564 2576
rect 18512 2533 18521 2567
rect 18521 2533 18555 2567
rect 18555 2533 18564 2567
rect 18512 2524 18564 2533
rect 18880 2524 18932 2576
rect 17316 2456 17368 2508
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 18788 2388 18840 2440
rect 1768 2252 1820 2304
rect 2320 2252 2372 2304
rect 2780 2252 2832 2304
rect 6000 2295 6052 2304
rect 6000 2261 6009 2295
rect 6009 2261 6043 2295
rect 6043 2261 6052 2295
rect 6000 2252 6052 2261
rect 9864 2252 9916 2304
rect 12348 2252 12400 2304
rect 18420 2252 18472 2304
rect 4648 2150 4700 2202
rect 4712 2150 4764 2202
rect 4776 2150 4828 2202
rect 4840 2150 4892 2202
rect 11982 2150 12034 2202
rect 12046 2150 12098 2202
rect 12110 2150 12162 2202
rect 12174 2150 12226 2202
rect 19315 2150 19367 2202
rect 19379 2150 19431 2202
rect 19443 2150 19495 2202
rect 19507 2150 19559 2202
rect 9772 2048 9824 2100
rect 15568 2048 15620 2100
rect 12348 76 12400 128
rect 15108 76 15160 128
<< metal2 >>
rect 1582 21570 1638 22000
rect 4710 21570 4766 22000
rect 7838 21570 7894 22000
rect 10966 21570 11022 22000
rect 14094 21570 14150 22000
rect 1320 21542 1638 21570
rect 1320 18222 1348 21542
rect 1582 21520 1638 21542
rect 4540 21542 4766 21570
rect 1582 20360 1638 20369
rect 1582 20295 1638 20304
rect 1596 18426 1624 20295
rect 4540 18426 4568 21542
rect 4710 21520 4766 21542
rect 7668 21542 7894 21570
rect 4622 19612 4918 19632
rect 4678 19610 4702 19612
rect 4758 19610 4782 19612
rect 4838 19610 4862 19612
rect 4700 19558 4702 19610
rect 4764 19558 4776 19610
rect 4838 19558 4840 19610
rect 4678 19556 4702 19558
rect 4758 19556 4782 19558
rect 4838 19556 4862 19558
rect 4622 19536 4918 19556
rect 4622 18524 4918 18544
rect 4678 18522 4702 18524
rect 4758 18522 4782 18524
rect 4838 18522 4862 18524
rect 4700 18470 4702 18522
rect 4764 18470 4776 18522
rect 4838 18470 4840 18522
rect 4678 18468 4702 18470
rect 4758 18468 4782 18470
rect 4838 18468 4862 18470
rect 4622 18448 4918 18468
rect 7668 18426 7696 21542
rect 7838 21520 7894 21542
rect 10888 21542 11022 21570
rect 8289 19068 8585 19088
rect 8345 19066 8369 19068
rect 8425 19066 8449 19068
rect 8505 19066 8529 19068
rect 8367 19014 8369 19066
rect 8431 19014 8443 19066
rect 8505 19014 8507 19066
rect 8345 19012 8369 19014
rect 8425 19012 8449 19014
rect 8505 19012 8529 19014
rect 8289 18992 8585 19012
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 1308 18216 1360 18222
rect 1308 18158 1360 18164
rect 1858 18184 1914 18193
rect 110 10160 166 10169
rect 110 10095 166 10104
rect 124 9897 152 10095
rect 110 9888 166 9897
rect 110 9823 166 9832
rect 1320 9042 1348 18158
rect 1858 18119 1914 18128
rect 1582 16008 1638 16017
rect 1582 15943 1638 15952
rect 1596 15706 1624 15943
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1412 14822 1440 15506
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 1308 9036 1360 9042
rect 1308 8978 1360 8984
rect 1320 8634 1348 8978
rect 1308 8628 1360 8634
rect 1308 8570 1360 8576
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 1688 6866 1716 7414
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 112 6656 164 6662
rect 112 6598 164 6604
rect 124 3369 152 6598
rect 1872 6458 1900 18119
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 4622 17436 4918 17456
rect 4678 17434 4702 17436
rect 4758 17434 4782 17436
rect 4838 17434 4862 17436
rect 4700 17382 4702 17434
rect 4764 17382 4776 17434
rect 4838 17382 4840 17434
rect 4678 17380 4702 17382
rect 4758 17380 4782 17382
rect 4838 17380 4862 17382
rect 4622 17360 4918 17380
rect 4622 16348 4918 16368
rect 4678 16346 4702 16348
rect 4758 16346 4782 16348
rect 4838 16346 4862 16348
rect 4700 16294 4702 16346
rect 4764 16294 4776 16346
rect 4838 16294 4840 16346
rect 4678 16292 4702 16294
rect 4758 16292 4782 16294
rect 4838 16292 4862 16294
rect 4622 16272 4918 16292
rect 4622 15260 4918 15280
rect 4678 15258 4702 15260
rect 4758 15258 4782 15260
rect 4838 15258 4862 15260
rect 4700 15206 4702 15258
rect 4764 15206 4776 15258
rect 4838 15206 4840 15258
rect 4678 15204 4702 15206
rect 4758 15204 4782 15206
rect 4838 15204 4862 15206
rect 4622 15184 4918 15204
rect 4622 14172 4918 14192
rect 4678 14170 4702 14172
rect 4758 14170 4782 14172
rect 4838 14170 4862 14172
rect 4700 14118 4702 14170
rect 4764 14118 4776 14170
rect 4838 14118 4840 14170
rect 4678 14116 4702 14118
rect 4758 14116 4782 14118
rect 4838 14116 4862 14118
rect 4622 14096 4918 14116
rect 4622 13084 4918 13104
rect 4678 13082 4702 13084
rect 4758 13082 4782 13084
rect 4838 13082 4862 13084
rect 4700 13030 4702 13082
rect 4764 13030 4776 13082
rect 4838 13030 4840 13082
rect 4678 13028 4702 13030
rect 4758 13028 4782 13030
rect 4838 13028 4862 13030
rect 4622 13008 4918 13028
rect 4622 11996 4918 12016
rect 4678 11994 4702 11996
rect 4758 11994 4782 11996
rect 4838 11994 4862 11996
rect 4700 11942 4702 11994
rect 4764 11942 4776 11994
rect 4838 11942 4840 11994
rect 4678 11940 4702 11942
rect 4758 11940 4782 11942
rect 4838 11940 4862 11942
rect 4622 11920 4918 11940
rect 2042 11656 2098 11665
rect 2042 11591 2098 11600
rect 2056 8498 2084 11591
rect 5276 11121 5304 18022
rect 8289 17980 8585 18000
rect 8345 17978 8369 17980
rect 8425 17978 8449 17980
rect 8505 17978 8529 17980
rect 8367 17926 8369 17978
rect 8431 17926 8443 17978
rect 8505 17926 8507 17978
rect 8345 17924 8369 17926
rect 8425 17924 8449 17926
rect 8505 17924 8529 17926
rect 8289 17904 8585 17924
rect 8289 16892 8585 16912
rect 8345 16890 8369 16892
rect 8425 16890 8449 16892
rect 8505 16890 8529 16892
rect 8367 16838 8369 16890
rect 8431 16838 8443 16890
rect 8505 16838 8507 16890
rect 8345 16836 8369 16838
rect 8425 16836 8449 16838
rect 8505 16836 8529 16838
rect 8289 16816 8585 16836
rect 8289 15804 8585 15824
rect 8345 15802 8369 15804
rect 8425 15802 8449 15804
rect 8505 15802 8529 15804
rect 8367 15750 8369 15802
rect 8431 15750 8443 15802
rect 8505 15750 8507 15802
rect 8345 15748 8369 15750
rect 8425 15748 8449 15750
rect 8505 15748 8529 15750
rect 8289 15728 8585 15748
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5262 11112 5318 11121
rect 5262 11047 5318 11056
rect 4622 10908 4918 10928
rect 4678 10906 4702 10908
rect 4758 10906 4782 10908
rect 4838 10906 4862 10908
rect 4700 10854 4702 10906
rect 4764 10854 4776 10906
rect 4838 10854 4840 10906
rect 4678 10852 4702 10854
rect 4758 10852 4782 10854
rect 4838 10852 4862 10854
rect 4622 10832 4918 10852
rect 4622 9820 4918 9840
rect 4678 9818 4702 9820
rect 4758 9818 4782 9820
rect 4838 9818 4862 9820
rect 4700 9766 4702 9818
rect 4764 9766 4776 9818
rect 4838 9766 4840 9818
rect 4678 9764 4702 9766
rect 4758 9764 4782 9766
rect 4838 9764 4862 9766
rect 4622 9744 4918 9764
rect 5276 9654 5304 11047
rect 5264 9648 5316 9654
rect 5264 9590 5316 9596
rect 5368 9518 5396 14758
rect 8289 14716 8585 14736
rect 8345 14714 8369 14716
rect 8425 14714 8449 14716
rect 8505 14714 8529 14716
rect 8367 14662 8369 14714
rect 8431 14662 8443 14714
rect 8505 14662 8507 14714
rect 8345 14660 8369 14662
rect 8425 14660 8449 14662
rect 8505 14660 8529 14662
rect 8289 14640 8585 14660
rect 8289 13628 8585 13648
rect 8345 13626 8369 13628
rect 8425 13626 8449 13628
rect 8505 13626 8529 13628
rect 8367 13574 8369 13626
rect 8431 13574 8443 13626
rect 8505 13574 8507 13626
rect 8345 13572 8369 13574
rect 8425 13572 8449 13574
rect 8505 13572 8529 13574
rect 8289 13552 8585 13572
rect 8289 12540 8585 12560
rect 8345 12538 8369 12540
rect 8425 12538 8449 12540
rect 8505 12538 8529 12540
rect 8367 12486 8369 12538
rect 8431 12486 8443 12538
rect 8505 12486 8507 12538
rect 8345 12484 8369 12486
rect 8425 12484 8449 12486
rect 8505 12484 8529 12486
rect 8289 12464 8585 12484
rect 8289 11452 8585 11472
rect 8345 11450 8369 11452
rect 8425 11450 8449 11452
rect 8505 11450 8529 11452
rect 8367 11398 8369 11450
rect 8431 11398 8443 11450
rect 8505 11398 8507 11450
rect 8345 11396 8369 11398
rect 8425 11396 8449 11398
rect 8505 11396 8529 11398
rect 8289 11376 8585 11396
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 10538 6960 10950
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 6012 9042 6040 10406
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 4622 8732 4918 8752
rect 4678 8730 4702 8732
rect 4758 8730 4782 8732
rect 4838 8730 4862 8732
rect 4700 8678 4702 8730
rect 4764 8678 4776 8730
rect 4838 8678 4840 8730
rect 4678 8676 4702 8678
rect 4758 8676 4782 8678
rect 4838 8676 4862 8678
rect 4622 8656 4918 8676
rect 6012 8634 6040 8978
rect 6288 8906 6316 9930
rect 6380 9722 6408 9998
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6564 9382 6592 10134
rect 6932 9654 6960 10474
rect 7576 10266 7604 10474
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7576 9654 7604 10202
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7760 9450 7788 10474
rect 8128 10198 8156 11086
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 8220 10198 8248 10542
rect 8289 10364 8585 10384
rect 8345 10362 8369 10364
rect 8425 10362 8449 10364
rect 8505 10362 8529 10364
rect 8367 10310 8369 10362
rect 8431 10310 8443 10362
rect 8505 10310 8507 10362
rect 8345 10308 8369 10310
rect 8425 10308 8449 10310
rect 8505 10308 8529 10310
rect 8289 10288 8585 10308
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 9402 10160 9458 10169
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2056 8276 2084 8434
rect 1964 8248 2084 8276
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 6089 1440 6190
rect 1768 6112 1820 6118
rect 1398 6080 1454 6089
rect 1768 6054 1820 6060
rect 1398 6015 1454 6024
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1596 4826 1624 5102
rect 848 4820 900 4826
rect 848 4762 900 4768
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 110 3360 166 3369
rect 110 3295 166 3304
rect 478 82 534 480
rect 860 82 888 4762
rect 1780 4146 1808 6054
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1872 5574 1900 5714
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1872 4010 1900 5510
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1872 3738 1900 3946
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1780 2650 1808 3334
rect 1964 3194 1992 8248
rect 3896 8090 3924 8502
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 2056 3534 2084 7142
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2148 5778 2176 6598
rect 2332 6254 2360 6598
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2424 6118 2452 7142
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2240 4826 2268 5306
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2424 4758 2452 5510
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2424 4282 2452 4694
rect 2700 4622 2728 7142
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 1964 2990 1992 3130
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 2332 2854 2360 3606
rect 2700 3126 2728 4558
rect 2792 3670 2820 6598
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 2976 5030 3004 5782
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2976 4282 3004 4966
rect 3068 4758 3096 7142
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3344 5098 3372 5646
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3528 5166 3556 5510
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3620 5098 3648 6598
rect 3712 5098 3740 7278
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3700 5092 3752 5098
rect 3700 5034 3752 5040
rect 3344 4826 3372 5034
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2976 3738 3004 4218
rect 3068 4010 3096 4694
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2688 3120 2740 3126
rect 2688 3062 2740 3068
rect 2792 2990 2820 3606
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 2332 2446 2360 2790
rect 3528 2650 3556 4966
rect 3620 4010 3648 5034
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3620 3194 3648 3946
rect 3712 3194 3740 5034
rect 3896 5030 3924 5510
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 3942 3924 4966
rect 3988 4010 4016 8230
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 4080 4282 4108 5578
rect 4172 4622 4200 8502
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4540 6730 4568 8366
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 4622 7644 4918 7664
rect 4678 7642 4702 7644
rect 4758 7642 4782 7644
rect 4838 7642 4862 7644
rect 4700 7590 4702 7642
rect 4764 7590 4776 7642
rect 4838 7590 4840 7642
rect 4678 7588 4702 7590
rect 4758 7588 4782 7590
rect 4838 7588 4862 7590
rect 4622 7568 4918 7588
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4356 5370 4384 6122
rect 4448 5574 4476 6190
rect 4540 5710 4568 6666
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 4622 6556 4918 6576
rect 4678 6554 4702 6556
rect 4758 6554 4782 6556
rect 4838 6554 4862 6556
rect 4700 6502 4702 6554
rect 4764 6502 4776 6554
rect 4838 6502 4840 6554
rect 4678 6500 4702 6502
rect 4758 6500 4782 6502
rect 4838 6500 4862 6502
rect 4622 6480 4918 6500
rect 5000 5778 5028 6598
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4264 4758 4292 5306
rect 4448 5030 4476 5510
rect 4540 5302 4568 5646
rect 4622 5468 4918 5488
rect 4678 5466 4702 5468
rect 4758 5466 4782 5468
rect 4838 5466 4862 5468
rect 4700 5414 4702 5466
rect 4764 5414 4776 5466
rect 4838 5414 4840 5466
rect 4678 5412 4702 5414
rect 4758 5412 4782 5414
rect 4838 5412 4862 5414
rect 4622 5392 4918 5412
rect 4528 5296 4580 5302
rect 4528 5238 4580 5244
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2332 2310 2360 2382
rect 1768 2304 1820 2310
rect 1768 2246 1820 2252
rect 2320 2304 2372 2310
rect 2320 2246 2372 2252
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 478 54 888 82
rect 1490 82 1546 480
rect 1780 82 1808 2246
rect 1490 54 1808 82
rect 2502 82 2558 480
rect 2792 82 2820 2246
rect 2502 54 2820 82
rect 3606 82 3662 480
rect 3896 82 3924 3878
rect 3988 2514 4016 3946
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4080 1737 4108 4218
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4356 3738 4384 3946
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4448 3398 4476 4966
rect 4540 4826 4568 5238
rect 5000 5098 5028 5714
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4622 4380 4918 4400
rect 4678 4378 4702 4380
rect 4758 4378 4782 4380
rect 4838 4378 4862 4380
rect 4700 4326 4702 4378
rect 4764 4326 4776 4378
rect 4838 4326 4840 4378
rect 4678 4324 4702 4326
rect 4758 4324 4782 4326
rect 4838 4324 4862 4326
rect 4622 4304 4918 4324
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4908 3738 4936 4150
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5092 3602 5120 8298
rect 6380 7993 6408 9318
rect 6564 9110 6592 9318
rect 7760 9178 7788 9386
rect 8128 9178 8156 10134
rect 8220 9722 8248 10134
rect 9402 10095 9458 10104
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8404 9586 8432 9998
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9232 9586 9260 9862
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 8289 9276 8585 9296
rect 8345 9274 8369 9276
rect 8425 9274 8449 9276
rect 8505 9274 8529 9276
rect 8367 9222 8369 9274
rect 8431 9222 8443 9274
rect 8505 9222 8507 9274
rect 8345 9220 8369 9222
rect 8425 9220 8449 9222
rect 8505 9220 8529 9222
rect 8289 9200 8585 9220
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6366 7984 6422 7993
rect 6366 7919 6422 7928
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5184 3738 5212 7686
rect 5276 7410 5304 7822
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5368 7274 5396 7686
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5552 7002 5580 7822
rect 6092 7200 6144 7206
rect 6144 7160 6224 7188
rect 6092 7142 6144 7148
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 6196 6866 6224 7160
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 5276 6118 5304 6802
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5368 5642 5396 6190
rect 5736 6186 5764 6802
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 6012 6118 6040 6802
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5828 5302 5856 6054
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5354 5128 5410 5137
rect 5354 5063 5410 5072
rect 5368 4690 5396 5063
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5552 4486 5580 5238
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5644 4826 5672 5170
rect 6012 5030 6040 5578
rect 6196 5234 6224 6802
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 4146 5580 4422
rect 5736 4282 5764 4626
rect 6380 4622 6408 6054
rect 6472 4826 6500 8774
rect 6840 8430 6868 8774
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 8022 6684 8230
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6748 6458 6776 6666
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6564 6118 6592 6258
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6000 4616 6052 4622
rect 5828 4576 6000 4604
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4540 2854 4568 3470
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4622 3292 4918 3312
rect 4678 3290 4702 3292
rect 4758 3290 4782 3292
rect 4838 3290 4862 3292
rect 4700 3238 4702 3290
rect 4764 3238 4776 3290
rect 4838 3238 4840 3290
rect 4678 3236 4702 3238
rect 4758 3236 4782 3238
rect 4838 3236 4862 3238
rect 4622 3216 4918 3236
rect 5000 3126 5028 3334
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 5000 2990 5028 3062
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4632 2650 4660 2858
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4622 2204 4918 2224
rect 4678 2202 4702 2204
rect 4758 2202 4782 2204
rect 4838 2202 4862 2204
rect 4700 2150 4702 2202
rect 4764 2150 4776 2202
rect 4838 2150 4840 2202
rect 4678 2148 4702 2150
rect 4758 2148 4782 2150
rect 4838 2148 4862 2150
rect 4622 2128 4918 2148
rect 4066 1728 4122 1737
rect 4066 1663 4122 1672
rect 3606 54 3924 82
rect 4618 82 4674 480
rect 5000 82 5028 2926
rect 5184 2514 5212 3674
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5276 2922 5304 3538
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 4618 54 5028 82
rect 5630 82 5686 480
rect 5736 82 5764 4218
rect 5828 4214 5856 4576
rect 6000 4558 6052 4564
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 6000 4004 6052 4010
rect 6000 3946 6052 3952
rect 6012 3602 6040 3946
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 6012 3194 6040 3538
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6012 2922 6040 3130
rect 6196 3126 6224 3878
rect 6380 3602 6408 4558
rect 6564 4078 6592 6054
rect 6840 5914 6868 8366
rect 7300 8362 7328 9114
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7944 7954 7972 8774
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 8036 8022 8064 8298
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7208 7274 7236 7686
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 6254 6960 6598
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6656 5030 6684 5646
rect 6932 5370 6960 6190
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6656 4690 6684 4966
rect 6932 4758 6960 5306
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 7024 4690 7052 5782
rect 7116 5098 7144 6326
rect 7208 5642 7236 7210
rect 7484 7206 7512 7278
rect 7944 7206 7972 7890
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7484 6866 7512 7142
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7484 6390 7512 6802
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 7208 5098 7236 5578
rect 7484 5574 7512 6326
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 6196 2582 6224 3062
rect 6380 2650 6408 3538
rect 6564 2990 6592 4014
rect 6656 3942 6684 4626
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6656 3534 6684 3878
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6184 2576 6236 2582
rect 6184 2518 6236 2524
rect 6932 2514 6960 3538
rect 7024 3466 7052 4626
rect 7116 3670 7144 5034
rect 7300 4826 7328 5510
rect 7484 5302 7512 5510
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7484 4214 7512 5238
rect 7576 4729 7604 6122
rect 7852 6118 7880 6666
rect 7944 6254 7972 6802
rect 8024 6792 8076 6798
rect 8128 6780 8156 8842
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9232 8566 9260 8774
rect 9220 8560 9272 8566
rect 9034 8528 9090 8537
rect 9220 8502 9272 8508
rect 9034 8463 9090 8472
rect 9048 8430 9076 8463
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8289 8188 8585 8208
rect 8345 8186 8369 8188
rect 8425 8186 8449 8188
rect 8505 8186 8529 8188
rect 8367 8134 8369 8186
rect 8431 8134 8443 8186
rect 8505 8134 8507 8186
rect 8345 8132 8369 8134
rect 8425 8132 8449 8134
rect 8505 8132 8529 8134
rect 8289 8112 8585 8132
rect 8680 7750 8708 8230
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8220 7342 8248 7686
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8496 7342 8524 7414
rect 8680 7342 8708 7686
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8076 6752 8156 6780
rect 8024 6734 8076 6740
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7944 6118 7972 6190
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7852 5778 7880 6054
rect 8128 5846 8156 6752
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7852 5302 7880 5714
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 8220 5166 8248 7278
rect 8289 7100 8585 7120
rect 8345 7098 8369 7100
rect 8425 7098 8449 7100
rect 8505 7098 8529 7100
rect 8367 7046 8369 7098
rect 8431 7046 8443 7098
rect 8505 7046 8507 7098
rect 8345 7044 8369 7046
rect 8425 7044 8449 7046
rect 8505 7044 8529 7046
rect 8289 7024 8585 7044
rect 8680 6866 8708 7278
rect 8772 6934 8800 7278
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8289 6012 8585 6032
rect 8345 6010 8369 6012
rect 8425 6010 8449 6012
rect 8505 6010 8529 6012
rect 8367 5958 8369 6010
rect 8431 5958 8443 6010
rect 8505 5958 8507 6010
rect 8345 5956 8369 5958
rect 8425 5956 8449 5958
rect 8505 5956 8529 5958
rect 8289 5936 8585 5956
rect 8772 5846 8800 6122
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8772 5370 8800 5782
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 7562 4720 7618 4729
rect 7562 4655 7618 4664
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7852 3942 7880 5102
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7944 3942 7972 4626
rect 8036 4010 8064 5102
rect 8289 4924 8585 4944
rect 8345 4922 8369 4924
rect 8425 4922 8449 4924
rect 8505 4922 8529 4924
rect 8367 4870 8369 4922
rect 8431 4870 8443 4922
rect 8505 4870 8507 4922
rect 8345 4868 8369 4870
rect 8425 4868 8449 4870
rect 8505 4868 8529 4870
rect 8289 4848 8585 4868
rect 8680 4808 8708 5238
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8588 4780 8708 4808
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7104 3664 7156 3670
rect 7104 3606 7156 3612
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 7116 2922 7144 3606
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 7760 2514 7788 3402
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 5998 2408 6054 2417
rect 5998 2343 6054 2352
rect 6460 2372 6512 2378
rect 6012 2310 6040 2343
rect 6460 2314 6512 2320
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 5630 54 5764 82
rect 6472 82 6500 2314
rect 6734 82 6790 480
rect 6472 54 6790 82
rect 478 0 534 54
rect 1490 0 1546 54
rect 2502 0 2558 54
rect 3606 0 3662 54
rect 4618 0 4674 54
rect 5630 0 5686 54
rect 6734 0 6790 54
rect 7746 82 7802 480
rect 7944 82 7972 3878
rect 8036 3058 8064 3946
rect 8128 3602 8156 4558
rect 8588 4486 8616 4780
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8220 3534 8248 4150
rect 8588 4078 8616 4422
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8289 3836 8585 3856
rect 8345 3834 8369 3836
rect 8425 3834 8449 3836
rect 8505 3834 8529 3836
rect 8367 3782 8369 3834
rect 8431 3782 8443 3834
rect 8505 3782 8507 3834
rect 8345 3780 8369 3782
rect 8425 3780 8449 3782
rect 8505 3780 8529 3782
rect 8289 3760 8585 3780
rect 8772 3602 8800 5170
rect 8864 4554 8892 5850
rect 9048 5166 9076 6802
rect 9140 5914 9168 7414
rect 9232 6322 9260 8502
rect 9324 7546 9352 9386
rect 9416 7834 9444 10095
rect 9600 10062 9628 10542
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9692 9178 9720 10950
rect 9784 10470 9812 11154
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 9784 10062 9812 10134
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9784 9722 9812 9998
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9508 8498 9536 8978
rect 9692 8498 9720 9114
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9784 8090 9812 8298
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9772 7880 9824 7886
rect 9416 7806 9536 7834
rect 9772 7822 9824 7828
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9220 6180 9272 6186
rect 9220 6122 9272 6128
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9140 5302 9168 5850
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9036 5160 9088 5166
rect 8956 5120 9036 5148
rect 8956 4690 8984 5120
rect 9232 5137 9260 6122
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9036 5102 9088 5108
rect 9218 5128 9274 5137
rect 9218 5063 9274 5072
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8864 4146 8892 4490
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8956 3738 8984 4422
rect 9048 4010 9076 4966
rect 9232 4865 9260 5063
rect 9218 4856 9274 4865
rect 9128 4820 9180 4826
rect 9218 4791 9274 4800
rect 9128 4762 9180 4768
rect 9140 4078 9168 4762
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9232 3670 9260 4626
rect 9324 4554 9352 6054
rect 9416 5846 9444 7686
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5166 9444 5510
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9312 4548 9364 4554
rect 9312 4490 9364 4496
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9508 4154 9536 7806
rect 9784 7002 9812 7822
rect 9876 7410 9904 9386
rect 10152 9382 10180 10134
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9968 7342 9996 8774
rect 10060 8090 10088 9046
rect 10152 8362 10180 9318
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 10060 7274 10088 8026
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 10060 6118 10088 7210
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9784 5166 9812 6054
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 8220 2990 8248 3470
rect 8772 3194 8800 3538
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 8220 2446 8248 2926
rect 8289 2748 8585 2768
rect 8345 2746 8369 2748
rect 8425 2746 8449 2748
rect 8505 2746 8529 2748
rect 8367 2694 8369 2746
rect 8431 2694 8443 2746
rect 8505 2694 8507 2746
rect 8345 2692 8369 2694
rect 8425 2692 8449 2694
rect 8505 2692 8529 2694
rect 8289 2672 8585 2692
rect 9048 2582 9076 2926
rect 9036 2576 9088 2582
rect 9036 2518 9088 2524
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 7746 54 7972 82
rect 8850 82 8906 480
rect 9324 116 9352 4150
rect 9416 4126 9536 4154
rect 9416 3602 9444 4126
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9508 2990 9536 4014
rect 9600 3942 9628 4966
rect 10152 4826 10180 5102
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10244 4154 10272 18022
rect 10322 16552 10378 16561
rect 10322 16487 10378 16496
rect 10336 10810 10364 16487
rect 10888 13814 10916 21542
rect 10966 21520 11022 21542
rect 13832 21542 14150 21570
rect 11956 19612 12252 19632
rect 12012 19610 12036 19612
rect 12092 19610 12116 19612
rect 12172 19610 12196 19612
rect 12034 19558 12036 19610
rect 12098 19558 12110 19610
rect 12172 19558 12174 19610
rect 12012 19556 12036 19558
rect 12092 19556 12116 19558
rect 12172 19556 12196 19558
rect 11956 19536 12252 19556
rect 11956 18524 12252 18544
rect 12012 18522 12036 18524
rect 12092 18522 12116 18524
rect 12172 18522 12196 18524
rect 12034 18470 12036 18522
rect 12098 18470 12110 18522
rect 12172 18470 12174 18522
rect 12012 18468 12036 18470
rect 12092 18468 12116 18470
rect 12172 18468 12196 18470
rect 11956 18448 12252 18468
rect 11956 17436 12252 17456
rect 12012 17434 12036 17436
rect 12092 17434 12116 17436
rect 12172 17434 12196 17436
rect 12034 17382 12036 17434
rect 12098 17382 12110 17434
rect 12172 17382 12174 17434
rect 12012 17380 12036 17382
rect 12092 17380 12116 17382
rect 12172 17380 12196 17382
rect 11956 17360 12252 17380
rect 11956 16348 12252 16368
rect 12012 16346 12036 16348
rect 12092 16346 12116 16348
rect 12172 16346 12196 16348
rect 12034 16294 12036 16346
rect 12098 16294 12110 16346
rect 12172 16294 12174 16346
rect 12012 16292 12036 16294
rect 12092 16292 12116 16294
rect 12172 16292 12196 16294
rect 11956 16272 12252 16292
rect 11956 15260 12252 15280
rect 12012 15258 12036 15260
rect 12092 15258 12116 15260
rect 12172 15258 12196 15260
rect 12034 15206 12036 15258
rect 12098 15206 12110 15258
rect 12172 15206 12174 15258
rect 12012 15204 12036 15206
rect 12092 15204 12116 15206
rect 12172 15204 12196 15206
rect 11956 15184 12252 15204
rect 11956 14172 12252 14192
rect 12012 14170 12036 14172
rect 12092 14170 12116 14172
rect 12172 14170 12196 14172
rect 12034 14118 12036 14170
rect 12098 14118 12110 14170
rect 12172 14118 12174 14170
rect 12012 14116 12036 14118
rect 12092 14116 12116 14118
rect 12172 14116 12196 14118
rect 11956 14096 12252 14116
rect 10888 13786 11008 13814
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10796 9994 10824 10406
rect 10888 10033 10916 10542
rect 10874 10024 10930 10033
rect 10784 9988 10836 9994
rect 10874 9959 10930 9968
rect 10784 9930 10836 9936
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10428 6254 10456 6802
rect 10520 6458 10548 8774
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10428 5574 10456 6190
rect 10520 5710 10548 6394
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10152 4126 10272 4154
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9876 3398 9904 3878
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9876 2922 9904 3334
rect 10060 3194 10088 3538
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 9784 2446 9812 2858
rect 9876 2582 9904 2858
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9876 2310 9904 2518
rect 10152 2446 10180 4126
rect 10336 2582 10364 4558
rect 10612 4486 10640 8842
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10704 5914 10732 6802
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10796 5370 10824 9930
rect 10980 9518 11008 13786
rect 13832 13394 13860 21542
rect 14094 21520 14150 21542
rect 16580 21548 16632 21554
rect 17222 21548 17278 22000
rect 20350 21570 20406 22000
rect 17222 21520 17224 21548
rect 16580 21490 16632 21496
rect 17276 21520 17278 21548
rect 20088 21542 20406 21570
rect 17224 21490 17276 21496
rect 15622 19068 15918 19088
rect 15678 19066 15702 19068
rect 15758 19066 15782 19068
rect 15838 19066 15862 19068
rect 15700 19014 15702 19066
rect 15764 19014 15776 19066
rect 15838 19014 15840 19066
rect 15678 19012 15702 19014
rect 15758 19012 15782 19014
rect 15838 19012 15862 19014
rect 15622 18992 15918 19012
rect 15622 17980 15918 18000
rect 15678 17978 15702 17980
rect 15758 17978 15782 17980
rect 15838 17978 15862 17980
rect 15700 17926 15702 17978
rect 15764 17926 15776 17978
rect 15838 17926 15840 17978
rect 15678 17924 15702 17926
rect 15758 17924 15782 17926
rect 15838 17924 15862 17926
rect 15622 17904 15918 17924
rect 15622 16892 15918 16912
rect 15678 16890 15702 16892
rect 15758 16890 15782 16892
rect 15838 16890 15862 16892
rect 15700 16838 15702 16890
rect 15764 16838 15776 16890
rect 15838 16838 15840 16890
rect 15678 16836 15702 16838
rect 15758 16836 15782 16838
rect 15838 16836 15862 16838
rect 15622 16816 15918 16836
rect 15622 15804 15918 15824
rect 15678 15802 15702 15804
rect 15758 15802 15782 15804
rect 15838 15802 15862 15804
rect 15700 15750 15702 15802
rect 15764 15750 15776 15802
rect 15838 15750 15840 15802
rect 15678 15748 15702 15750
rect 15758 15748 15782 15750
rect 15838 15748 15862 15750
rect 15622 15728 15918 15748
rect 15106 15056 15162 15065
rect 15106 14991 15162 15000
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 11956 13084 12252 13104
rect 12012 13082 12036 13084
rect 12092 13082 12116 13084
rect 12172 13082 12196 13084
rect 12034 13030 12036 13082
rect 12098 13030 12110 13082
rect 12172 13030 12174 13082
rect 12012 13028 12036 13030
rect 12092 13028 12116 13030
rect 12172 13028 12196 13030
rect 11956 13008 12252 13028
rect 11956 11996 12252 12016
rect 12012 11994 12036 11996
rect 12092 11994 12116 11996
rect 12172 11994 12196 11996
rect 12034 11942 12036 11994
rect 12098 11942 12110 11994
rect 12172 11942 12174 11994
rect 12012 11940 12036 11942
rect 12092 11940 12116 11942
rect 12172 11940 12196 11942
rect 11956 11920 12252 11940
rect 11956 10908 12252 10928
rect 12012 10906 12036 10908
rect 12092 10906 12116 10908
rect 12172 10906 12196 10908
rect 12034 10854 12036 10906
rect 12098 10854 12110 10906
rect 12172 10854 12174 10906
rect 12012 10852 12036 10854
rect 12092 10852 12116 10854
rect 12172 10852 12196 10854
rect 11956 10832 12252 10852
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10888 7857 10916 8366
rect 11072 8294 11100 8910
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10874 7848 10930 7857
rect 10874 7783 10930 7792
rect 10888 7478 10916 7783
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10888 6866 10916 7142
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 11072 6390 11100 8230
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10888 4826 10916 5782
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 10980 5370 11008 5510
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11072 5114 11100 5510
rect 10980 5086 11100 5114
rect 10980 5030 11008 5086
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 10704 2514 10732 3606
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10980 3194 11008 3470
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 9772 2100 9824 2106
rect 9772 2042 9824 2048
rect 9232 88 9352 116
rect 9232 82 9260 88
rect 8850 54 9260 82
rect 9784 82 9812 2042
rect 9862 82 9918 480
rect 9784 54 9918 82
rect 7746 0 7802 54
rect 8850 0 8906 54
rect 9862 0 9918 54
rect 10874 82 10930 480
rect 11072 82 11100 4966
rect 11164 4214 11192 9318
rect 11348 8974 11376 10406
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 11956 9820 12252 9840
rect 12012 9818 12036 9820
rect 12092 9818 12116 9820
rect 12172 9818 12196 9820
rect 12034 9766 12036 9818
rect 12098 9766 12110 9818
rect 12172 9766 12174 9818
rect 12012 9764 12036 9766
rect 12092 9764 12116 9766
rect 12172 9764 12196 9766
rect 11956 9744 12252 9764
rect 12360 9722 12388 10066
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11440 8566 11468 9386
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11624 8022 11652 8230
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11532 7750 11560 7822
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11532 7002 11560 7686
rect 11624 7342 11652 7958
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11256 6254 11284 6734
rect 11808 6254 11836 9454
rect 11956 8732 12252 8752
rect 12012 8730 12036 8732
rect 12092 8730 12116 8732
rect 12172 8730 12196 8732
rect 12034 8678 12036 8730
rect 12098 8678 12110 8730
rect 12172 8678 12174 8730
rect 12012 8676 12036 8678
rect 12092 8676 12116 8678
rect 12172 8676 12196 8678
rect 11956 8656 12252 8676
rect 12360 7750 12388 9658
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 11956 7644 12252 7664
rect 12012 7642 12036 7644
rect 12092 7642 12116 7644
rect 12172 7642 12196 7644
rect 12034 7590 12036 7642
rect 12098 7590 12110 7642
rect 12172 7590 12174 7642
rect 12012 7588 12036 7590
rect 12092 7588 12116 7590
rect 12172 7588 12196 7590
rect 11956 7568 12252 7588
rect 12452 7426 12480 9862
rect 12728 9586 12756 10406
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 12636 9110 12664 9386
rect 12912 9382 12940 10406
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12636 7818 12664 8298
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 13004 7546 13032 13330
rect 15120 11121 15148 14991
rect 15622 14716 15918 14736
rect 15678 14714 15702 14716
rect 15758 14714 15782 14716
rect 15838 14714 15862 14716
rect 15700 14662 15702 14714
rect 15764 14662 15776 14714
rect 15838 14662 15840 14714
rect 15678 14660 15702 14662
rect 15758 14660 15782 14662
rect 15838 14660 15862 14662
rect 15622 14640 15918 14660
rect 15622 13628 15918 13648
rect 15678 13626 15702 13628
rect 15758 13626 15782 13628
rect 15838 13626 15862 13628
rect 15700 13574 15702 13626
rect 15764 13574 15776 13626
rect 15838 13574 15840 13626
rect 15678 13572 15702 13574
rect 15758 13572 15782 13574
rect 15838 13572 15862 13574
rect 15622 13552 15918 13572
rect 15622 12540 15918 12560
rect 15678 12538 15702 12540
rect 15758 12538 15782 12540
rect 15838 12538 15862 12540
rect 15700 12486 15702 12538
rect 15764 12486 15776 12538
rect 15838 12486 15840 12538
rect 15678 12484 15702 12486
rect 15758 12484 15782 12486
rect 15838 12484 15862 12486
rect 15622 12464 15918 12484
rect 15622 11452 15918 11472
rect 15678 11450 15702 11452
rect 15758 11450 15782 11452
rect 15838 11450 15862 11452
rect 15700 11398 15702 11450
rect 15764 11398 15776 11450
rect 15838 11398 15840 11450
rect 15678 11396 15702 11398
rect 15758 11396 15782 11398
rect 15838 11396 15862 11398
rect 15622 11376 15918 11396
rect 15106 11112 15162 11121
rect 15106 11047 15162 11056
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13188 8498 13216 9386
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13464 8634 13492 9046
rect 13556 8906 13584 9998
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13740 9586 13768 9930
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13556 7886 13584 8842
rect 14108 8362 14136 9114
rect 15120 9042 15148 11047
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15120 8634 15148 8978
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 8022 13952 8230
rect 13912 8016 13964 8022
rect 13912 7958 13964 7964
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12360 7398 12480 7426
rect 12360 6866 12388 7398
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12728 6866 12756 7142
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11256 4758 11284 6054
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11256 3942 11284 4694
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11348 3602 11376 4490
rect 11624 3924 11652 6054
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11716 4690 11744 5850
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11808 4214 11836 5782
rect 11900 5778 11928 6802
rect 11956 6556 12252 6576
rect 12012 6554 12036 6556
rect 12092 6554 12116 6556
rect 12172 6554 12196 6556
rect 12034 6502 12036 6554
rect 12098 6502 12110 6554
rect 12172 6502 12174 6554
rect 12012 6500 12036 6502
rect 12092 6500 12116 6502
rect 12172 6500 12196 6502
rect 11956 6480 12252 6500
rect 12728 6322 12756 6802
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 11992 5778 12020 6258
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11992 5658 12020 5714
rect 11900 5630 12020 5658
rect 11900 5302 11928 5630
rect 11956 5468 12252 5488
rect 12012 5466 12036 5468
rect 12092 5466 12116 5468
rect 12172 5466 12196 5468
rect 12034 5414 12036 5466
rect 12098 5414 12110 5466
rect 12172 5414 12174 5466
rect 12012 5412 12036 5414
rect 12092 5412 12116 5414
rect 12172 5412 12196 5414
rect 11956 5392 12252 5412
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 12360 4758 12388 5782
rect 12544 5778 12572 5850
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 11956 4380 12252 4400
rect 12012 4378 12036 4380
rect 12092 4378 12116 4380
rect 12172 4378 12196 4380
rect 12034 4326 12036 4378
rect 12098 4326 12110 4378
rect 12172 4326 12174 4378
rect 12012 4324 12036 4326
rect 12092 4324 12116 4326
rect 12172 4324 12196 4326
rect 11956 4304 12252 4324
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12176 4049 12204 4082
rect 12162 4040 12218 4049
rect 12636 4010 12664 5646
rect 12728 5302 12756 6258
rect 12912 6118 12940 6802
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12820 5574 12848 5714
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12716 5296 12768 5302
rect 12716 5238 12768 5244
rect 12162 3975 12218 3984
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 11704 3936 11756 3942
rect 11624 3896 11704 3924
rect 11704 3878 11756 3884
rect 11716 3602 11744 3878
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 11164 3398 11192 3538
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11164 3126 11192 3334
rect 11348 3194 11376 3538
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 11164 2446 11192 3062
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11532 2553 11560 2586
rect 11518 2544 11574 2553
rect 11518 2479 11574 2488
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 10874 54 11100 82
rect 11716 82 11744 3334
rect 11808 2446 11836 3538
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 11956 3292 12252 3312
rect 12012 3290 12036 3292
rect 12092 3290 12116 3292
rect 12172 3290 12196 3292
rect 12034 3238 12036 3290
rect 12098 3238 12110 3290
rect 12172 3238 12174 3290
rect 12012 3236 12036 3238
rect 12092 3236 12116 3238
rect 12172 3236 12196 3238
rect 11956 3216 12252 3236
rect 12360 3058 12388 3470
rect 12820 3466 12848 5510
rect 13004 5370 13032 7482
rect 13464 7342 13492 7822
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 13648 7546 13676 7686
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13648 7342 13676 7482
rect 15120 7342 15148 7686
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 13464 7002 13492 7278
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 14016 6254 14044 7278
rect 14660 6866 14688 7278
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14016 5846 14044 6190
rect 14660 5914 14688 6802
rect 15120 6254 15148 7278
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15120 5914 15148 6190
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 14004 5840 14056 5846
rect 13924 5800 14004 5828
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 13188 5098 13216 5714
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13740 5166 13768 5646
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12256 2916 12308 2922
rect 12256 2858 12308 2864
rect 12268 2514 12296 2858
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12360 2446 12388 2994
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 11956 2204 12252 2224
rect 12012 2202 12036 2204
rect 12092 2202 12116 2204
rect 12172 2202 12196 2204
rect 12034 2150 12036 2202
rect 12098 2150 12110 2202
rect 12172 2150 12174 2202
rect 12012 2148 12036 2150
rect 12092 2148 12116 2150
rect 12172 2148 12196 2150
rect 11956 2128 12252 2148
rect 11978 82 12034 480
rect 12360 134 12388 2246
rect 11716 54 12034 82
rect 12348 128 12400 134
rect 12348 70 12400 76
rect 12912 82 12940 4966
rect 13924 4758 13952 5800
rect 14004 5782 14056 5788
rect 14660 5166 14688 5850
rect 15120 5166 15148 5850
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 15108 5160 15160 5166
rect 15108 5102 15160 5108
rect 14660 4758 14688 5102
rect 13912 4752 13964 4758
rect 14648 4752 14700 4758
rect 13912 4694 13964 4700
rect 14002 4720 14058 4729
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13360 4684 13412 4690
rect 13360 4626 13412 4632
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13096 4214 13124 4626
rect 13372 4554 13400 4626
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13360 4548 13412 4554
rect 13360 4490 13412 4496
rect 13648 4282 13676 4558
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 13096 3602 13124 4150
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13096 2990 13124 3538
rect 13280 3534 13308 3674
rect 13556 3534 13584 3946
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13280 3194 13308 3470
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13740 2990 13768 4626
rect 13924 4078 13952 4694
rect 14648 4694 14700 4700
rect 15120 4690 15148 5102
rect 14096 4684 14148 4690
rect 14058 4664 14096 4672
rect 14002 4655 14096 4664
rect 14016 4644 14096 4655
rect 14096 4626 14148 4632
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 13832 2990 13860 3402
rect 14016 3058 14044 3674
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 13372 2514 13400 2858
rect 13636 2576 13688 2582
rect 13740 2564 13768 2926
rect 14004 2916 14056 2922
rect 14004 2858 14056 2864
rect 14016 2582 14044 2858
rect 13688 2536 13768 2564
rect 14004 2576 14056 2582
rect 13636 2518 13688 2524
rect 14004 2518 14056 2524
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 12990 82 13046 480
rect 12912 54 13046 82
rect 10874 0 10930 54
rect 11978 0 12034 54
rect 12990 0 13046 54
rect 14002 82 14058 480
rect 14108 82 14136 4150
rect 14936 4078 14964 4626
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14384 3738 14412 4014
rect 14844 3942 14872 4014
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14200 2514 14228 2994
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14844 1465 14872 3878
rect 14936 3738 14964 4014
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 15016 3664 15068 3670
rect 15016 3606 15068 3612
rect 15028 3194 15056 3606
rect 15120 3534 15148 4422
rect 15212 4049 15240 9318
rect 15396 8838 15424 10406
rect 15622 10364 15918 10384
rect 15678 10362 15702 10364
rect 15758 10362 15782 10364
rect 15838 10362 15862 10364
rect 15700 10310 15702 10362
rect 15764 10310 15776 10362
rect 15838 10310 15840 10362
rect 15678 10308 15702 10310
rect 15758 10308 15782 10310
rect 15838 10308 15862 10310
rect 15622 10288 15918 10308
rect 16592 9722 16620 21490
rect 17236 21459 17264 21490
rect 19154 20496 19210 20505
rect 19154 20431 19210 20440
rect 19062 18728 19118 18737
rect 19062 18663 19118 18672
rect 17774 16824 17830 16833
rect 17774 16759 17830 16768
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 17788 9586 17816 16759
rect 19076 13394 19104 18663
rect 19064 13388 19116 13394
rect 19064 13330 19116 13336
rect 19076 12646 19104 13330
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 18524 9518 18552 12582
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 19076 10470 19104 11154
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 17776 9444 17828 9450
rect 17776 9386 17828 9392
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 15622 9276 15918 9296
rect 15678 9274 15702 9276
rect 15758 9274 15782 9276
rect 15838 9274 15862 9276
rect 15700 9222 15702 9274
rect 15764 9222 15776 9274
rect 15838 9222 15840 9274
rect 15678 9220 15702 9222
rect 15758 9220 15782 9222
rect 15838 9220 15862 9222
rect 15622 9200 15918 9220
rect 15948 9110 15976 9318
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 16580 9104 16632 9110
rect 16580 9046 16632 9052
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 8634 16252 8774
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 15622 8188 15918 8208
rect 15678 8186 15702 8188
rect 15758 8186 15782 8188
rect 15838 8186 15862 8188
rect 15700 8134 15702 8186
rect 15764 8134 15776 8186
rect 15838 8134 15840 8186
rect 15678 8132 15702 8134
rect 15758 8132 15782 8134
rect 15838 8132 15862 8134
rect 15622 8112 15918 8132
rect 15948 8090 15976 8230
rect 16316 8090 16344 9046
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 8498 16528 8774
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16592 8022 16620 9046
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16960 8090 16988 8298
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15304 7002 15332 7822
rect 16040 7206 16068 7958
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 7410 16528 7686
rect 16960 7546 16988 8026
rect 17236 7886 17264 9318
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 15622 7100 15918 7120
rect 15678 7098 15702 7100
rect 15758 7098 15782 7100
rect 15838 7098 15862 7100
rect 15700 7046 15702 7098
rect 15764 7046 15776 7098
rect 15838 7046 15840 7098
rect 15678 7044 15702 7046
rect 15758 7044 15782 7046
rect 15838 7044 15862 7046
rect 15622 7024 15918 7044
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15488 5914 15516 6802
rect 15764 6458 15792 6802
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15948 6118 15976 6802
rect 16040 6168 16068 7142
rect 16224 6866 16252 7278
rect 17236 7002 17264 7822
rect 17328 7546 17356 7958
rect 17420 7886 17448 8298
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16224 6322 16252 6598
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16120 6180 16172 6186
rect 16040 6140 16120 6168
rect 16120 6122 16172 6128
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15622 6012 15918 6032
rect 15678 6010 15702 6012
rect 15758 6010 15782 6012
rect 15838 6010 15862 6012
rect 15700 5958 15702 6010
rect 15764 5958 15776 6010
rect 15838 5958 15840 6010
rect 15678 5956 15702 5958
rect 15758 5956 15782 5958
rect 15838 5956 15862 5958
rect 15622 5936 15918 5956
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15488 5710 15516 5850
rect 16132 5846 16160 6122
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16120 5840 16172 5846
rect 16120 5782 16172 5788
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15672 5234 15700 5646
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15304 4214 15332 4762
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15198 4040 15254 4049
rect 15198 3975 15254 3984
rect 15396 3942 15424 4966
rect 15622 4924 15918 4944
rect 15678 4922 15702 4924
rect 15758 4922 15782 4924
rect 15838 4922 15862 4924
rect 15700 4870 15702 4922
rect 15764 4870 15776 4922
rect 15838 4870 15840 4922
rect 15678 4868 15702 4870
rect 15758 4868 15782 4870
rect 15838 4868 15862 4870
rect 15474 4856 15530 4865
rect 15622 4848 15918 4868
rect 15474 4791 15530 4800
rect 15488 4214 15516 4791
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15016 3188 15068 3194
rect 15016 3130 15068 3136
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14936 2553 14964 2926
rect 15028 2582 15056 3130
rect 15396 2922 15424 3878
rect 15488 3534 15516 4150
rect 15622 3836 15918 3856
rect 15678 3834 15702 3836
rect 15758 3834 15782 3836
rect 15838 3834 15862 3836
rect 15700 3782 15702 3834
rect 15764 3782 15776 3834
rect 15838 3782 15840 3834
rect 15678 3780 15702 3782
rect 15758 3780 15782 3782
rect 15838 3780 15862 3782
rect 15622 3760 15918 3780
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 15622 2748 15918 2768
rect 15678 2746 15702 2748
rect 15758 2746 15782 2748
rect 15838 2746 15862 2748
rect 15700 2694 15702 2746
rect 15764 2694 15776 2746
rect 15838 2694 15840 2746
rect 15678 2692 15702 2694
rect 15758 2692 15782 2694
rect 15838 2692 15862 2694
rect 15622 2672 15918 2692
rect 15016 2576 15068 2582
rect 14922 2544 14978 2553
rect 15016 2518 15068 2524
rect 15474 2544 15530 2553
rect 14922 2479 14978 2488
rect 15384 2508 15436 2514
rect 15436 2488 15474 2496
rect 15436 2479 15530 2488
rect 15568 2508 15620 2514
rect 15436 2468 15516 2479
rect 15384 2450 15436 2456
rect 15568 2450 15620 2456
rect 15580 2106 15608 2450
rect 15568 2100 15620 2106
rect 15568 2042 15620 2048
rect 14830 1456 14886 1465
rect 14830 1391 14886 1400
rect 14002 54 14136 82
rect 15106 128 15162 480
rect 15106 76 15108 128
rect 15160 76 15162 128
rect 14002 0 14058 54
rect 15106 0 15162 76
rect 15948 82 15976 5578
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 16040 4826 16068 5102
rect 16132 5030 16160 5782
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16132 4758 16160 4966
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 16224 2514 16252 6054
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17420 5370 17448 5850
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 16316 4010 16344 4694
rect 16776 4690 16804 5170
rect 17408 4752 17460 4758
rect 17328 4712 17408 4740
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16408 4010 16436 4626
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16408 3738 16436 3946
rect 16684 3738 16712 4558
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17144 3194 17172 3606
rect 17328 3398 17356 4712
rect 17408 4694 17460 4700
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17420 4214 17448 4558
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17420 3942 17448 4150
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17236 3194 17264 3334
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 16684 2689 16712 2790
rect 16670 2680 16726 2689
rect 16670 2615 16726 2624
rect 16684 2582 16712 2615
rect 16672 2576 16724 2582
rect 16672 2518 16724 2524
rect 17328 2514 17356 2994
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 16118 82 16174 480
rect 15948 54 16174 82
rect 16118 0 16174 54
rect 17222 82 17278 480
rect 17512 82 17540 7482
rect 17788 7410 17816 9386
rect 17880 9042 17908 9454
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18340 9178 18368 9318
rect 19168 9178 19196 20431
rect 19289 19612 19585 19632
rect 19345 19610 19369 19612
rect 19425 19610 19449 19612
rect 19505 19610 19529 19612
rect 19367 19558 19369 19610
rect 19431 19558 19443 19610
rect 19505 19558 19507 19610
rect 19345 19556 19369 19558
rect 19425 19556 19449 19558
rect 19505 19556 19529 19558
rect 19289 19536 19585 19556
rect 19289 18524 19585 18544
rect 19345 18522 19369 18524
rect 19425 18522 19449 18524
rect 19505 18522 19529 18524
rect 19367 18470 19369 18522
rect 19431 18470 19443 18522
rect 19505 18470 19507 18522
rect 19345 18468 19369 18470
rect 19425 18468 19449 18470
rect 19505 18468 19529 18470
rect 19289 18448 19585 18468
rect 19289 17436 19585 17456
rect 19345 17434 19369 17436
rect 19425 17434 19449 17436
rect 19505 17434 19529 17436
rect 19367 17382 19369 17434
rect 19431 17382 19443 17434
rect 19505 17382 19507 17434
rect 19345 17380 19369 17382
rect 19425 17380 19449 17382
rect 19505 17380 19529 17382
rect 19289 17360 19585 17380
rect 20088 16561 20116 21542
rect 20350 21520 20406 21542
rect 20074 16552 20130 16561
rect 20074 16487 20130 16496
rect 19289 16348 19585 16368
rect 19345 16346 19369 16348
rect 19425 16346 19449 16348
rect 19505 16346 19529 16348
rect 19367 16294 19369 16346
rect 19431 16294 19443 16346
rect 19505 16294 19507 16346
rect 19345 16292 19369 16294
rect 19425 16292 19449 16294
rect 19505 16292 19529 16294
rect 19289 16272 19585 16292
rect 19289 15260 19585 15280
rect 19345 15258 19369 15260
rect 19425 15258 19449 15260
rect 19505 15258 19529 15260
rect 19367 15206 19369 15258
rect 19431 15206 19443 15258
rect 19505 15206 19507 15258
rect 19345 15204 19369 15206
rect 19425 15204 19449 15206
rect 19505 15204 19529 15206
rect 19289 15184 19585 15204
rect 19289 14172 19585 14192
rect 19345 14170 19369 14172
rect 19425 14170 19449 14172
rect 19505 14170 19529 14172
rect 19367 14118 19369 14170
rect 19431 14118 19443 14170
rect 19505 14118 19507 14170
rect 19345 14116 19369 14118
rect 19425 14116 19449 14118
rect 19505 14116 19529 14118
rect 19289 14096 19585 14116
rect 19246 13560 19302 13569
rect 19246 13495 19302 13504
rect 19260 13258 19288 13495
rect 19248 13252 19300 13258
rect 19248 13194 19300 13200
rect 19289 13084 19585 13104
rect 19345 13082 19369 13084
rect 19425 13082 19449 13084
rect 19505 13082 19529 13084
rect 19367 13030 19369 13082
rect 19431 13030 19443 13082
rect 19505 13030 19507 13082
rect 19345 13028 19369 13030
rect 19425 13028 19449 13030
rect 19505 13028 19529 13030
rect 19289 13008 19585 13028
rect 19289 11996 19585 12016
rect 19345 11994 19369 11996
rect 19425 11994 19449 11996
rect 19505 11994 19529 11996
rect 19367 11942 19369 11994
rect 19431 11942 19443 11994
rect 19505 11942 19507 11994
rect 19345 11940 19369 11942
rect 19425 11940 19449 11942
rect 19505 11940 19529 11942
rect 19289 11920 19585 11940
rect 19338 11520 19394 11529
rect 19338 11455 19394 11464
rect 19352 11354 19380 11455
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19289 10908 19585 10928
rect 19345 10906 19369 10908
rect 19425 10906 19449 10908
rect 19505 10906 19529 10908
rect 19367 10854 19369 10906
rect 19431 10854 19443 10906
rect 19505 10854 19507 10906
rect 19345 10852 19369 10854
rect 19425 10852 19449 10854
rect 19505 10852 19529 10854
rect 19289 10832 19585 10852
rect 21546 10024 21602 10033
rect 21546 9959 21602 9968
rect 19289 9820 19585 9840
rect 19345 9818 19369 9820
rect 19425 9818 19449 9820
rect 19505 9818 19529 9820
rect 19367 9766 19369 9818
rect 19431 9766 19443 9818
rect 19505 9766 19507 9818
rect 19345 9764 19369 9766
rect 19425 9764 19449 9766
rect 19505 9764 19529 9766
rect 19289 9744 19585 9764
rect 21560 9654 21588 9959
rect 21548 9648 21600 9654
rect 21548 9590 21600 9596
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 19156 9036 19208 9042
rect 19260 9024 19288 9454
rect 19208 8996 19288 9024
rect 19156 8978 19208 8984
rect 17880 8362 17908 8978
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18432 8498 18460 8910
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 17880 8265 17908 8298
rect 17866 8256 17922 8265
rect 17866 8191 17922 8200
rect 18248 8090 18276 8298
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17776 6928 17828 6934
rect 17776 6870 17828 6876
rect 17788 6458 17816 6870
rect 18156 6798 18184 7686
rect 18432 6934 18460 8434
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18602 7984 18658 7993
rect 18602 7919 18604 7928
rect 18656 7919 18658 7928
rect 18604 7890 18656 7896
rect 18616 7274 18644 7890
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18604 7268 18656 7274
rect 18604 7210 18656 7216
rect 18420 6928 18472 6934
rect 18420 6870 18472 6876
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17788 6186 17816 6394
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 18156 5914 18184 6734
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18432 5710 18460 6870
rect 18604 6724 18656 6730
rect 18604 6666 18656 6672
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17776 4616 17828 4622
rect 17776 4558 17828 4564
rect 17696 4146 17724 4558
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17696 3738 17724 4082
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17788 3670 17816 4558
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18156 4146 18184 4218
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18248 4010 18276 4490
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 17684 3460 17736 3466
rect 17684 3402 17736 3408
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17604 2922 17632 3334
rect 17696 3058 17724 3402
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 17592 2916 17644 2922
rect 17592 2858 17644 2864
rect 17696 2582 17724 2994
rect 17788 2990 17816 3402
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 18432 2922 18460 5306
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 18420 2916 18472 2922
rect 18420 2858 18472 2864
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17684 2576 17736 2582
rect 17684 2518 17736 2524
rect 17788 2417 17816 2790
rect 17880 2650 17908 2858
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 18524 2582 18552 5646
rect 18512 2576 18564 2582
rect 18512 2518 18564 2524
rect 18420 2440 18472 2446
rect 17774 2408 17830 2417
rect 18420 2382 18472 2388
rect 17774 2343 17830 2352
rect 18432 2310 18460 2382
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 17222 54 17540 82
rect 18234 82 18290 480
rect 18616 82 18644 6666
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18708 6458 18736 6598
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18800 6322 18828 7822
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18800 5914 18828 6258
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18800 5234 18828 5850
rect 18892 5778 18920 8366
rect 19168 8294 19196 8978
rect 19289 8732 19585 8752
rect 19345 8730 19369 8732
rect 19425 8730 19449 8732
rect 19505 8730 19529 8732
rect 19367 8678 19369 8730
rect 19431 8678 19443 8730
rect 19505 8678 19507 8730
rect 19345 8676 19369 8678
rect 19425 8676 19449 8678
rect 19505 8676 19529 8678
rect 19289 8656 19585 8676
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18892 5302 18920 5714
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 18708 2553 18736 3606
rect 18800 3040 18828 4218
rect 18892 4146 18920 5238
rect 18984 4154 19012 7142
rect 19168 6905 19196 8230
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19289 7644 19585 7664
rect 19345 7642 19369 7644
rect 19425 7642 19449 7644
rect 19505 7642 19529 7644
rect 19367 7590 19369 7642
rect 19431 7590 19443 7642
rect 19505 7590 19507 7642
rect 19345 7588 19369 7590
rect 19425 7588 19449 7590
rect 19505 7588 19529 7590
rect 19289 7568 19585 7588
rect 19154 6896 19210 6905
rect 19064 6860 19116 6866
rect 19154 6831 19210 6840
rect 19064 6802 19116 6808
rect 19076 6118 19104 6802
rect 19289 6556 19585 6576
rect 19345 6554 19369 6556
rect 19425 6554 19449 6556
rect 19505 6554 19529 6556
rect 19367 6502 19369 6554
rect 19431 6502 19443 6554
rect 19505 6502 19507 6554
rect 19345 6500 19369 6502
rect 19425 6500 19449 6502
rect 19505 6500 19529 6502
rect 19289 6480 19585 6500
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 19076 5370 19104 5714
rect 19289 5468 19585 5488
rect 19345 5466 19369 5468
rect 19425 5466 19449 5468
rect 19505 5466 19529 5468
rect 19367 5414 19369 5466
rect 19431 5414 19443 5466
rect 19505 5414 19507 5466
rect 19345 5412 19369 5414
rect 19425 5412 19449 5414
rect 19505 5412 19529 5414
rect 19289 5392 19585 5412
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 19076 4282 19104 4626
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 18880 4140 18932 4146
rect 18984 4126 19104 4154
rect 18880 4082 18932 4088
rect 18878 4040 18934 4049
rect 18878 3975 18934 3984
rect 18892 3534 18920 3975
rect 18880 3528 18932 3534
rect 18932 3488 19012 3516
rect 18880 3470 18932 3476
rect 18800 3012 18920 3040
rect 18788 2916 18840 2922
rect 18788 2858 18840 2864
rect 18694 2544 18750 2553
rect 18694 2479 18750 2488
rect 18800 2446 18828 2858
rect 18892 2689 18920 3012
rect 18984 2990 19012 3488
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 18878 2680 18934 2689
rect 18878 2615 18934 2624
rect 18892 2582 18920 2615
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 18234 54 18644 82
rect 19076 82 19104 4126
rect 19168 3194 19196 4966
rect 19289 4380 19585 4400
rect 19345 4378 19369 4380
rect 19425 4378 19449 4380
rect 19505 4378 19529 4380
rect 19367 4326 19369 4378
rect 19431 4326 19443 4378
rect 19505 4326 19507 4378
rect 19345 4324 19369 4326
rect 19425 4324 19449 4326
rect 19505 4324 19529 4326
rect 19289 4304 19585 4324
rect 19628 4214 19656 7822
rect 19720 6254 19748 9522
rect 21456 8356 21508 8362
rect 21456 8298 21508 8304
rect 19800 7268 19852 7274
rect 19800 7210 19852 7216
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19812 5137 19840 7210
rect 19798 5128 19854 5137
rect 19798 5063 19854 5072
rect 19616 4208 19668 4214
rect 19616 4150 19668 4156
rect 19616 4072 19668 4078
rect 19616 4014 19668 4020
rect 19628 3738 19656 4014
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 19289 3292 19585 3312
rect 19345 3290 19369 3292
rect 19425 3290 19449 3292
rect 19505 3290 19529 3292
rect 19367 3238 19369 3290
rect 19431 3238 19443 3290
rect 19505 3238 19507 3290
rect 19345 3236 19369 3238
rect 19425 3236 19449 3238
rect 19505 3236 19529 3238
rect 19289 3216 19585 3236
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19444 2553 19472 2790
rect 19430 2544 19486 2553
rect 19430 2479 19486 2488
rect 19289 2204 19585 2224
rect 19345 2202 19369 2204
rect 19425 2202 19449 2204
rect 19505 2202 19529 2204
rect 19367 2150 19369 2202
rect 19431 2150 19443 2202
rect 19505 2150 19507 2202
rect 19345 2148 19369 2150
rect 19425 2148 19449 2150
rect 19505 2148 19529 2150
rect 19289 2128 19585 2148
rect 19246 82 19302 480
rect 19076 54 19302 82
rect 20180 82 20208 3946
rect 20350 82 20406 480
rect 20180 54 20406 82
rect 17222 0 17278 54
rect 18234 0 18290 54
rect 19246 0 19302 54
rect 20350 0 20406 54
rect 21362 82 21418 480
rect 21468 82 21496 8298
rect 21548 2916 21600 2922
rect 21548 2858 21600 2864
rect 21560 2689 21588 2858
rect 21546 2680 21602 2689
rect 21546 2615 21602 2624
rect 21362 54 21496 82
rect 21362 0 21418 54
<< via2 >>
rect 1582 20304 1638 20360
rect 4622 19610 4678 19612
rect 4702 19610 4758 19612
rect 4782 19610 4838 19612
rect 4862 19610 4918 19612
rect 4622 19558 4648 19610
rect 4648 19558 4678 19610
rect 4702 19558 4712 19610
rect 4712 19558 4758 19610
rect 4782 19558 4828 19610
rect 4828 19558 4838 19610
rect 4862 19558 4892 19610
rect 4892 19558 4918 19610
rect 4622 19556 4678 19558
rect 4702 19556 4758 19558
rect 4782 19556 4838 19558
rect 4862 19556 4918 19558
rect 4622 18522 4678 18524
rect 4702 18522 4758 18524
rect 4782 18522 4838 18524
rect 4862 18522 4918 18524
rect 4622 18470 4648 18522
rect 4648 18470 4678 18522
rect 4702 18470 4712 18522
rect 4712 18470 4758 18522
rect 4782 18470 4828 18522
rect 4828 18470 4838 18522
rect 4862 18470 4892 18522
rect 4892 18470 4918 18522
rect 4622 18468 4678 18470
rect 4702 18468 4758 18470
rect 4782 18468 4838 18470
rect 4862 18468 4918 18470
rect 8289 19066 8345 19068
rect 8369 19066 8425 19068
rect 8449 19066 8505 19068
rect 8529 19066 8585 19068
rect 8289 19014 8315 19066
rect 8315 19014 8345 19066
rect 8369 19014 8379 19066
rect 8379 19014 8425 19066
rect 8449 19014 8495 19066
rect 8495 19014 8505 19066
rect 8529 19014 8559 19066
rect 8559 19014 8585 19066
rect 8289 19012 8345 19014
rect 8369 19012 8425 19014
rect 8449 19012 8505 19014
rect 8529 19012 8585 19014
rect 110 10104 166 10160
rect 110 9832 166 9888
rect 1858 18128 1914 18184
rect 1582 15952 1638 16008
rect 4622 17434 4678 17436
rect 4702 17434 4758 17436
rect 4782 17434 4838 17436
rect 4862 17434 4918 17436
rect 4622 17382 4648 17434
rect 4648 17382 4678 17434
rect 4702 17382 4712 17434
rect 4712 17382 4758 17434
rect 4782 17382 4828 17434
rect 4828 17382 4838 17434
rect 4862 17382 4892 17434
rect 4892 17382 4918 17434
rect 4622 17380 4678 17382
rect 4702 17380 4758 17382
rect 4782 17380 4838 17382
rect 4862 17380 4918 17382
rect 4622 16346 4678 16348
rect 4702 16346 4758 16348
rect 4782 16346 4838 16348
rect 4862 16346 4918 16348
rect 4622 16294 4648 16346
rect 4648 16294 4678 16346
rect 4702 16294 4712 16346
rect 4712 16294 4758 16346
rect 4782 16294 4828 16346
rect 4828 16294 4838 16346
rect 4862 16294 4892 16346
rect 4892 16294 4918 16346
rect 4622 16292 4678 16294
rect 4702 16292 4758 16294
rect 4782 16292 4838 16294
rect 4862 16292 4918 16294
rect 4622 15258 4678 15260
rect 4702 15258 4758 15260
rect 4782 15258 4838 15260
rect 4862 15258 4918 15260
rect 4622 15206 4648 15258
rect 4648 15206 4678 15258
rect 4702 15206 4712 15258
rect 4712 15206 4758 15258
rect 4782 15206 4828 15258
rect 4828 15206 4838 15258
rect 4862 15206 4892 15258
rect 4892 15206 4918 15258
rect 4622 15204 4678 15206
rect 4702 15204 4758 15206
rect 4782 15204 4838 15206
rect 4862 15204 4918 15206
rect 4622 14170 4678 14172
rect 4702 14170 4758 14172
rect 4782 14170 4838 14172
rect 4862 14170 4918 14172
rect 4622 14118 4648 14170
rect 4648 14118 4678 14170
rect 4702 14118 4712 14170
rect 4712 14118 4758 14170
rect 4782 14118 4828 14170
rect 4828 14118 4838 14170
rect 4862 14118 4892 14170
rect 4892 14118 4918 14170
rect 4622 14116 4678 14118
rect 4702 14116 4758 14118
rect 4782 14116 4838 14118
rect 4862 14116 4918 14118
rect 4622 13082 4678 13084
rect 4702 13082 4758 13084
rect 4782 13082 4838 13084
rect 4862 13082 4918 13084
rect 4622 13030 4648 13082
rect 4648 13030 4678 13082
rect 4702 13030 4712 13082
rect 4712 13030 4758 13082
rect 4782 13030 4828 13082
rect 4828 13030 4838 13082
rect 4862 13030 4892 13082
rect 4892 13030 4918 13082
rect 4622 13028 4678 13030
rect 4702 13028 4758 13030
rect 4782 13028 4838 13030
rect 4862 13028 4918 13030
rect 4622 11994 4678 11996
rect 4702 11994 4758 11996
rect 4782 11994 4838 11996
rect 4862 11994 4918 11996
rect 4622 11942 4648 11994
rect 4648 11942 4678 11994
rect 4702 11942 4712 11994
rect 4712 11942 4758 11994
rect 4782 11942 4828 11994
rect 4828 11942 4838 11994
rect 4862 11942 4892 11994
rect 4892 11942 4918 11994
rect 4622 11940 4678 11942
rect 4702 11940 4758 11942
rect 4782 11940 4838 11942
rect 4862 11940 4918 11942
rect 2042 11600 2098 11656
rect 8289 17978 8345 17980
rect 8369 17978 8425 17980
rect 8449 17978 8505 17980
rect 8529 17978 8585 17980
rect 8289 17926 8315 17978
rect 8315 17926 8345 17978
rect 8369 17926 8379 17978
rect 8379 17926 8425 17978
rect 8449 17926 8495 17978
rect 8495 17926 8505 17978
rect 8529 17926 8559 17978
rect 8559 17926 8585 17978
rect 8289 17924 8345 17926
rect 8369 17924 8425 17926
rect 8449 17924 8505 17926
rect 8529 17924 8585 17926
rect 8289 16890 8345 16892
rect 8369 16890 8425 16892
rect 8449 16890 8505 16892
rect 8529 16890 8585 16892
rect 8289 16838 8315 16890
rect 8315 16838 8345 16890
rect 8369 16838 8379 16890
rect 8379 16838 8425 16890
rect 8449 16838 8495 16890
rect 8495 16838 8505 16890
rect 8529 16838 8559 16890
rect 8559 16838 8585 16890
rect 8289 16836 8345 16838
rect 8369 16836 8425 16838
rect 8449 16836 8505 16838
rect 8529 16836 8585 16838
rect 8289 15802 8345 15804
rect 8369 15802 8425 15804
rect 8449 15802 8505 15804
rect 8529 15802 8585 15804
rect 8289 15750 8315 15802
rect 8315 15750 8345 15802
rect 8369 15750 8379 15802
rect 8379 15750 8425 15802
rect 8449 15750 8495 15802
rect 8495 15750 8505 15802
rect 8529 15750 8559 15802
rect 8559 15750 8585 15802
rect 8289 15748 8345 15750
rect 8369 15748 8425 15750
rect 8449 15748 8505 15750
rect 8529 15748 8585 15750
rect 5262 11056 5318 11112
rect 4622 10906 4678 10908
rect 4702 10906 4758 10908
rect 4782 10906 4838 10908
rect 4862 10906 4918 10908
rect 4622 10854 4648 10906
rect 4648 10854 4678 10906
rect 4702 10854 4712 10906
rect 4712 10854 4758 10906
rect 4782 10854 4828 10906
rect 4828 10854 4838 10906
rect 4862 10854 4892 10906
rect 4892 10854 4918 10906
rect 4622 10852 4678 10854
rect 4702 10852 4758 10854
rect 4782 10852 4838 10854
rect 4862 10852 4918 10854
rect 4622 9818 4678 9820
rect 4702 9818 4758 9820
rect 4782 9818 4838 9820
rect 4862 9818 4918 9820
rect 4622 9766 4648 9818
rect 4648 9766 4678 9818
rect 4702 9766 4712 9818
rect 4712 9766 4758 9818
rect 4782 9766 4828 9818
rect 4828 9766 4838 9818
rect 4862 9766 4892 9818
rect 4892 9766 4918 9818
rect 4622 9764 4678 9766
rect 4702 9764 4758 9766
rect 4782 9764 4838 9766
rect 4862 9764 4918 9766
rect 8289 14714 8345 14716
rect 8369 14714 8425 14716
rect 8449 14714 8505 14716
rect 8529 14714 8585 14716
rect 8289 14662 8315 14714
rect 8315 14662 8345 14714
rect 8369 14662 8379 14714
rect 8379 14662 8425 14714
rect 8449 14662 8495 14714
rect 8495 14662 8505 14714
rect 8529 14662 8559 14714
rect 8559 14662 8585 14714
rect 8289 14660 8345 14662
rect 8369 14660 8425 14662
rect 8449 14660 8505 14662
rect 8529 14660 8585 14662
rect 8289 13626 8345 13628
rect 8369 13626 8425 13628
rect 8449 13626 8505 13628
rect 8529 13626 8585 13628
rect 8289 13574 8315 13626
rect 8315 13574 8345 13626
rect 8369 13574 8379 13626
rect 8379 13574 8425 13626
rect 8449 13574 8495 13626
rect 8495 13574 8505 13626
rect 8529 13574 8559 13626
rect 8559 13574 8585 13626
rect 8289 13572 8345 13574
rect 8369 13572 8425 13574
rect 8449 13572 8505 13574
rect 8529 13572 8585 13574
rect 8289 12538 8345 12540
rect 8369 12538 8425 12540
rect 8449 12538 8505 12540
rect 8529 12538 8585 12540
rect 8289 12486 8315 12538
rect 8315 12486 8345 12538
rect 8369 12486 8379 12538
rect 8379 12486 8425 12538
rect 8449 12486 8495 12538
rect 8495 12486 8505 12538
rect 8529 12486 8559 12538
rect 8559 12486 8585 12538
rect 8289 12484 8345 12486
rect 8369 12484 8425 12486
rect 8449 12484 8505 12486
rect 8529 12484 8585 12486
rect 8289 11450 8345 11452
rect 8369 11450 8425 11452
rect 8449 11450 8505 11452
rect 8529 11450 8585 11452
rect 8289 11398 8315 11450
rect 8315 11398 8345 11450
rect 8369 11398 8379 11450
rect 8379 11398 8425 11450
rect 8449 11398 8495 11450
rect 8495 11398 8505 11450
rect 8529 11398 8559 11450
rect 8559 11398 8585 11450
rect 8289 11396 8345 11398
rect 8369 11396 8425 11398
rect 8449 11396 8505 11398
rect 8529 11396 8585 11398
rect 4622 8730 4678 8732
rect 4702 8730 4758 8732
rect 4782 8730 4838 8732
rect 4862 8730 4918 8732
rect 4622 8678 4648 8730
rect 4648 8678 4678 8730
rect 4702 8678 4712 8730
rect 4712 8678 4758 8730
rect 4782 8678 4828 8730
rect 4828 8678 4838 8730
rect 4862 8678 4892 8730
rect 4892 8678 4918 8730
rect 4622 8676 4678 8678
rect 4702 8676 4758 8678
rect 4782 8676 4838 8678
rect 4862 8676 4918 8678
rect 8289 10362 8345 10364
rect 8369 10362 8425 10364
rect 8449 10362 8505 10364
rect 8529 10362 8585 10364
rect 8289 10310 8315 10362
rect 8315 10310 8345 10362
rect 8369 10310 8379 10362
rect 8379 10310 8425 10362
rect 8449 10310 8495 10362
rect 8495 10310 8505 10362
rect 8529 10310 8559 10362
rect 8559 10310 8585 10362
rect 8289 10308 8345 10310
rect 8369 10308 8425 10310
rect 8449 10308 8505 10310
rect 8529 10308 8585 10310
rect 1398 6024 1454 6080
rect 110 3304 166 3360
rect 4622 7642 4678 7644
rect 4702 7642 4758 7644
rect 4782 7642 4838 7644
rect 4862 7642 4918 7644
rect 4622 7590 4648 7642
rect 4648 7590 4678 7642
rect 4702 7590 4712 7642
rect 4712 7590 4758 7642
rect 4782 7590 4828 7642
rect 4828 7590 4838 7642
rect 4862 7590 4892 7642
rect 4892 7590 4918 7642
rect 4622 7588 4678 7590
rect 4702 7588 4758 7590
rect 4782 7588 4838 7590
rect 4862 7588 4918 7590
rect 4622 6554 4678 6556
rect 4702 6554 4758 6556
rect 4782 6554 4838 6556
rect 4862 6554 4918 6556
rect 4622 6502 4648 6554
rect 4648 6502 4678 6554
rect 4702 6502 4712 6554
rect 4712 6502 4758 6554
rect 4782 6502 4828 6554
rect 4828 6502 4838 6554
rect 4862 6502 4892 6554
rect 4892 6502 4918 6554
rect 4622 6500 4678 6502
rect 4702 6500 4758 6502
rect 4782 6500 4838 6502
rect 4862 6500 4918 6502
rect 4622 5466 4678 5468
rect 4702 5466 4758 5468
rect 4782 5466 4838 5468
rect 4862 5466 4918 5468
rect 4622 5414 4648 5466
rect 4648 5414 4678 5466
rect 4702 5414 4712 5466
rect 4712 5414 4758 5466
rect 4782 5414 4828 5466
rect 4828 5414 4838 5466
rect 4862 5414 4892 5466
rect 4892 5414 4918 5466
rect 4622 5412 4678 5414
rect 4702 5412 4758 5414
rect 4782 5412 4838 5414
rect 4862 5412 4918 5414
rect 4622 4378 4678 4380
rect 4702 4378 4758 4380
rect 4782 4378 4838 4380
rect 4862 4378 4918 4380
rect 4622 4326 4648 4378
rect 4648 4326 4678 4378
rect 4702 4326 4712 4378
rect 4712 4326 4758 4378
rect 4782 4326 4828 4378
rect 4828 4326 4838 4378
rect 4862 4326 4892 4378
rect 4892 4326 4918 4378
rect 4622 4324 4678 4326
rect 4702 4324 4758 4326
rect 4782 4324 4838 4326
rect 4862 4324 4918 4326
rect 9402 10104 9458 10160
rect 8289 9274 8345 9276
rect 8369 9274 8425 9276
rect 8449 9274 8505 9276
rect 8529 9274 8585 9276
rect 8289 9222 8315 9274
rect 8315 9222 8345 9274
rect 8369 9222 8379 9274
rect 8379 9222 8425 9274
rect 8449 9222 8495 9274
rect 8495 9222 8505 9274
rect 8529 9222 8559 9274
rect 8559 9222 8585 9274
rect 8289 9220 8345 9222
rect 8369 9220 8425 9222
rect 8449 9220 8505 9222
rect 8529 9220 8585 9222
rect 6366 7928 6422 7984
rect 5354 5072 5410 5128
rect 4622 3290 4678 3292
rect 4702 3290 4758 3292
rect 4782 3290 4838 3292
rect 4862 3290 4918 3292
rect 4622 3238 4648 3290
rect 4648 3238 4678 3290
rect 4702 3238 4712 3290
rect 4712 3238 4758 3290
rect 4782 3238 4828 3290
rect 4828 3238 4838 3290
rect 4862 3238 4892 3290
rect 4892 3238 4918 3290
rect 4622 3236 4678 3238
rect 4702 3236 4758 3238
rect 4782 3236 4838 3238
rect 4862 3236 4918 3238
rect 4622 2202 4678 2204
rect 4702 2202 4758 2204
rect 4782 2202 4838 2204
rect 4862 2202 4918 2204
rect 4622 2150 4648 2202
rect 4648 2150 4678 2202
rect 4702 2150 4712 2202
rect 4712 2150 4758 2202
rect 4782 2150 4828 2202
rect 4828 2150 4838 2202
rect 4862 2150 4892 2202
rect 4892 2150 4918 2202
rect 4622 2148 4678 2150
rect 4702 2148 4758 2150
rect 4782 2148 4838 2150
rect 4862 2148 4918 2150
rect 4066 1672 4122 1728
rect 9034 8472 9090 8528
rect 8289 8186 8345 8188
rect 8369 8186 8425 8188
rect 8449 8186 8505 8188
rect 8529 8186 8585 8188
rect 8289 8134 8315 8186
rect 8315 8134 8345 8186
rect 8369 8134 8379 8186
rect 8379 8134 8425 8186
rect 8449 8134 8495 8186
rect 8495 8134 8505 8186
rect 8529 8134 8559 8186
rect 8559 8134 8585 8186
rect 8289 8132 8345 8134
rect 8369 8132 8425 8134
rect 8449 8132 8505 8134
rect 8529 8132 8585 8134
rect 8289 7098 8345 7100
rect 8369 7098 8425 7100
rect 8449 7098 8505 7100
rect 8529 7098 8585 7100
rect 8289 7046 8315 7098
rect 8315 7046 8345 7098
rect 8369 7046 8379 7098
rect 8379 7046 8425 7098
rect 8449 7046 8495 7098
rect 8495 7046 8505 7098
rect 8529 7046 8559 7098
rect 8559 7046 8585 7098
rect 8289 7044 8345 7046
rect 8369 7044 8425 7046
rect 8449 7044 8505 7046
rect 8529 7044 8585 7046
rect 8289 6010 8345 6012
rect 8369 6010 8425 6012
rect 8449 6010 8505 6012
rect 8529 6010 8585 6012
rect 8289 5958 8315 6010
rect 8315 5958 8345 6010
rect 8369 5958 8379 6010
rect 8379 5958 8425 6010
rect 8449 5958 8495 6010
rect 8495 5958 8505 6010
rect 8529 5958 8559 6010
rect 8559 5958 8585 6010
rect 8289 5956 8345 5958
rect 8369 5956 8425 5958
rect 8449 5956 8505 5958
rect 8529 5956 8585 5958
rect 7562 4664 7618 4720
rect 8289 4922 8345 4924
rect 8369 4922 8425 4924
rect 8449 4922 8505 4924
rect 8529 4922 8585 4924
rect 8289 4870 8315 4922
rect 8315 4870 8345 4922
rect 8369 4870 8379 4922
rect 8379 4870 8425 4922
rect 8449 4870 8495 4922
rect 8495 4870 8505 4922
rect 8529 4870 8559 4922
rect 8559 4870 8585 4922
rect 8289 4868 8345 4870
rect 8369 4868 8425 4870
rect 8449 4868 8505 4870
rect 8529 4868 8585 4870
rect 5998 2352 6054 2408
rect 8289 3834 8345 3836
rect 8369 3834 8425 3836
rect 8449 3834 8505 3836
rect 8529 3834 8585 3836
rect 8289 3782 8315 3834
rect 8315 3782 8345 3834
rect 8369 3782 8379 3834
rect 8379 3782 8425 3834
rect 8449 3782 8495 3834
rect 8495 3782 8505 3834
rect 8529 3782 8559 3834
rect 8559 3782 8585 3834
rect 8289 3780 8345 3782
rect 8369 3780 8425 3782
rect 8449 3780 8505 3782
rect 8529 3780 8585 3782
rect 9218 5072 9274 5128
rect 9218 4800 9274 4856
rect 8289 2746 8345 2748
rect 8369 2746 8425 2748
rect 8449 2746 8505 2748
rect 8529 2746 8585 2748
rect 8289 2694 8315 2746
rect 8315 2694 8345 2746
rect 8369 2694 8379 2746
rect 8379 2694 8425 2746
rect 8449 2694 8495 2746
rect 8495 2694 8505 2746
rect 8529 2694 8559 2746
rect 8559 2694 8585 2746
rect 8289 2692 8345 2694
rect 8369 2692 8425 2694
rect 8449 2692 8505 2694
rect 8529 2692 8585 2694
rect 10322 16496 10378 16552
rect 11956 19610 12012 19612
rect 12036 19610 12092 19612
rect 12116 19610 12172 19612
rect 12196 19610 12252 19612
rect 11956 19558 11982 19610
rect 11982 19558 12012 19610
rect 12036 19558 12046 19610
rect 12046 19558 12092 19610
rect 12116 19558 12162 19610
rect 12162 19558 12172 19610
rect 12196 19558 12226 19610
rect 12226 19558 12252 19610
rect 11956 19556 12012 19558
rect 12036 19556 12092 19558
rect 12116 19556 12172 19558
rect 12196 19556 12252 19558
rect 11956 18522 12012 18524
rect 12036 18522 12092 18524
rect 12116 18522 12172 18524
rect 12196 18522 12252 18524
rect 11956 18470 11982 18522
rect 11982 18470 12012 18522
rect 12036 18470 12046 18522
rect 12046 18470 12092 18522
rect 12116 18470 12162 18522
rect 12162 18470 12172 18522
rect 12196 18470 12226 18522
rect 12226 18470 12252 18522
rect 11956 18468 12012 18470
rect 12036 18468 12092 18470
rect 12116 18468 12172 18470
rect 12196 18468 12252 18470
rect 11956 17434 12012 17436
rect 12036 17434 12092 17436
rect 12116 17434 12172 17436
rect 12196 17434 12252 17436
rect 11956 17382 11982 17434
rect 11982 17382 12012 17434
rect 12036 17382 12046 17434
rect 12046 17382 12092 17434
rect 12116 17382 12162 17434
rect 12162 17382 12172 17434
rect 12196 17382 12226 17434
rect 12226 17382 12252 17434
rect 11956 17380 12012 17382
rect 12036 17380 12092 17382
rect 12116 17380 12172 17382
rect 12196 17380 12252 17382
rect 11956 16346 12012 16348
rect 12036 16346 12092 16348
rect 12116 16346 12172 16348
rect 12196 16346 12252 16348
rect 11956 16294 11982 16346
rect 11982 16294 12012 16346
rect 12036 16294 12046 16346
rect 12046 16294 12092 16346
rect 12116 16294 12162 16346
rect 12162 16294 12172 16346
rect 12196 16294 12226 16346
rect 12226 16294 12252 16346
rect 11956 16292 12012 16294
rect 12036 16292 12092 16294
rect 12116 16292 12172 16294
rect 12196 16292 12252 16294
rect 11956 15258 12012 15260
rect 12036 15258 12092 15260
rect 12116 15258 12172 15260
rect 12196 15258 12252 15260
rect 11956 15206 11982 15258
rect 11982 15206 12012 15258
rect 12036 15206 12046 15258
rect 12046 15206 12092 15258
rect 12116 15206 12162 15258
rect 12162 15206 12172 15258
rect 12196 15206 12226 15258
rect 12226 15206 12252 15258
rect 11956 15204 12012 15206
rect 12036 15204 12092 15206
rect 12116 15204 12172 15206
rect 12196 15204 12252 15206
rect 11956 14170 12012 14172
rect 12036 14170 12092 14172
rect 12116 14170 12172 14172
rect 12196 14170 12252 14172
rect 11956 14118 11982 14170
rect 11982 14118 12012 14170
rect 12036 14118 12046 14170
rect 12046 14118 12092 14170
rect 12116 14118 12162 14170
rect 12162 14118 12172 14170
rect 12196 14118 12226 14170
rect 12226 14118 12252 14170
rect 11956 14116 12012 14118
rect 12036 14116 12092 14118
rect 12116 14116 12172 14118
rect 12196 14116 12252 14118
rect 10874 9968 10930 10024
rect 15622 19066 15678 19068
rect 15702 19066 15758 19068
rect 15782 19066 15838 19068
rect 15862 19066 15918 19068
rect 15622 19014 15648 19066
rect 15648 19014 15678 19066
rect 15702 19014 15712 19066
rect 15712 19014 15758 19066
rect 15782 19014 15828 19066
rect 15828 19014 15838 19066
rect 15862 19014 15892 19066
rect 15892 19014 15918 19066
rect 15622 19012 15678 19014
rect 15702 19012 15758 19014
rect 15782 19012 15838 19014
rect 15862 19012 15918 19014
rect 15622 17978 15678 17980
rect 15702 17978 15758 17980
rect 15782 17978 15838 17980
rect 15862 17978 15918 17980
rect 15622 17926 15648 17978
rect 15648 17926 15678 17978
rect 15702 17926 15712 17978
rect 15712 17926 15758 17978
rect 15782 17926 15828 17978
rect 15828 17926 15838 17978
rect 15862 17926 15892 17978
rect 15892 17926 15918 17978
rect 15622 17924 15678 17926
rect 15702 17924 15758 17926
rect 15782 17924 15838 17926
rect 15862 17924 15918 17926
rect 15622 16890 15678 16892
rect 15702 16890 15758 16892
rect 15782 16890 15838 16892
rect 15862 16890 15918 16892
rect 15622 16838 15648 16890
rect 15648 16838 15678 16890
rect 15702 16838 15712 16890
rect 15712 16838 15758 16890
rect 15782 16838 15828 16890
rect 15828 16838 15838 16890
rect 15862 16838 15892 16890
rect 15892 16838 15918 16890
rect 15622 16836 15678 16838
rect 15702 16836 15758 16838
rect 15782 16836 15838 16838
rect 15862 16836 15918 16838
rect 15622 15802 15678 15804
rect 15702 15802 15758 15804
rect 15782 15802 15838 15804
rect 15862 15802 15918 15804
rect 15622 15750 15648 15802
rect 15648 15750 15678 15802
rect 15702 15750 15712 15802
rect 15712 15750 15758 15802
rect 15782 15750 15828 15802
rect 15828 15750 15838 15802
rect 15862 15750 15892 15802
rect 15892 15750 15918 15802
rect 15622 15748 15678 15750
rect 15702 15748 15758 15750
rect 15782 15748 15838 15750
rect 15862 15748 15918 15750
rect 15106 15000 15162 15056
rect 11956 13082 12012 13084
rect 12036 13082 12092 13084
rect 12116 13082 12172 13084
rect 12196 13082 12252 13084
rect 11956 13030 11982 13082
rect 11982 13030 12012 13082
rect 12036 13030 12046 13082
rect 12046 13030 12092 13082
rect 12116 13030 12162 13082
rect 12162 13030 12172 13082
rect 12196 13030 12226 13082
rect 12226 13030 12252 13082
rect 11956 13028 12012 13030
rect 12036 13028 12092 13030
rect 12116 13028 12172 13030
rect 12196 13028 12252 13030
rect 11956 11994 12012 11996
rect 12036 11994 12092 11996
rect 12116 11994 12172 11996
rect 12196 11994 12252 11996
rect 11956 11942 11982 11994
rect 11982 11942 12012 11994
rect 12036 11942 12046 11994
rect 12046 11942 12092 11994
rect 12116 11942 12162 11994
rect 12162 11942 12172 11994
rect 12196 11942 12226 11994
rect 12226 11942 12252 11994
rect 11956 11940 12012 11942
rect 12036 11940 12092 11942
rect 12116 11940 12172 11942
rect 12196 11940 12252 11942
rect 11956 10906 12012 10908
rect 12036 10906 12092 10908
rect 12116 10906 12172 10908
rect 12196 10906 12252 10908
rect 11956 10854 11982 10906
rect 11982 10854 12012 10906
rect 12036 10854 12046 10906
rect 12046 10854 12092 10906
rect 12116 10854 12162 10906
rect 12162 10854 12172 10906
rect 12196 10854 12226 10906
rect 12226 10854 12252 10906
rect 11956 10852 12012 10854
rect 12036 10852 12092 10854
rect 12116 10852 12172 10854
rect 12196 10852 12252 10854
rect 10874 7792 10930 7848
rect 11956 9818 12012 9820
rect 12036 9818 12092 9820
rect 12116 9818 12172 9820
rect 12196 9818 12252 9820
rect 11956 9766 11982 9818
rect 11982 9766 12012 9818
rect 12036 9766 12046 9818
rect 12046 9766 12092 9818
rect 12116 9766 12162 9818
rect 12162 9766 12172 9818
rect 12196 9766 12226 9818
rect 12226 9766 12252 9818
rect 11956 9764 12012 9766
rect 12036 9764 12092 9766
rect 12116 9764 12172 9766
rect 12196 9764 12252 9766
rect 11956 8730 12012 8732
rect 12036 8730 12092 8732
rect 12116 8730 12172 8732
rect 12196 8730 12252 8732
rect 11956 8678 11982 8730
rect 11982 8678 12012 8730
rect 12036 8678 12046 8730
rect 12046 8678 12092 8730
rect 12116 8678 12162 8730
rect 12162 8678 12172 8730
rect 12196 8678 12226 8730
rect 12226 8678 12252 8730
rect 11956 8676 12012 8678
rect 12036 8676 12092 8678
rect 12116 8676 12172 8678
rect 12196 8676 12252 8678
rect 11956 7642 12012 7644
rect 12036 7642 12092 7644
rect 12116 7642 12172 7644
rect 12196 7642 12252 7644
rect 11956 7590 11982 7642
rect 11982 7590 12012 7642
rect 12036 7590 12046 7642
rect 12046 7590 12092 7642
rect 12116 7590 12162 7642
rect 12162 7590 12172 7642
rect 12196 7590 12226 7642
rect 12226 7590 12252 7642
rect 11956 7588 12012 7590
rect 12036 7588 12092 7590
rect 12116 7588 12172 7590
rect 12196 7588 12252 7590
rect 15622 14714 15678 14716
rect 15702 14714 15758 14716
rect 15782 14714 15838 14716
rect 15862 14714 15918 14716
rect 15622 14662 15648 14714
rect 15648 14662 15678 14714
rect 15702 14662 15712 14714
rect 15712 14662 15758 14714
rect 15782 14662 15828 14714
rect 15828 14662 15838 14714
rect 15862 14662 15892 14714
rect 15892 14662 15918 14714
rect 15622 14660 15678 14662
rect 15702 14660 15758 14662
rect 15782 14660 15838 14662
rect 15862 14660 15918 14662
rect 15622 13626 15678 13628
rect 15702 13626 15758 13628
rect 15782 13626 15838 13628
rect 15862 13626 15918 13628
rect 15622 13574 15648 13626
rect 15648 13574 15678 13626
rect 15702 13574 15712 13626
rect 15712 13574 15758 13626
rect 15782 13574 15828 13626
rect 15828 13574 15838 13626
rect 15862 13574 15892 13626
rect 15892 13574 15918 13626
rect 15622 13572 15678 13574
rect 15702 13572 15758 13574
rect 15782 13572 15838 13574
rect 15862 13572 15918 13574
rect 15622 12538 15678 12540
rect 15702 12538 15758 12540
rect 15782 12538 15838 12540
rect 15862 12538 15918 12540
rect 15622 12486 15648 12538
rect 15648 12486 15678 12538
rect 15702 12486 15712 12538
rect 15712 12486 15758 12538
rect 15782 12486 15828 12538
rect 15828 12486 15838 12538
rect 15862 12486 15892 12538
rect 15892 12486 15918 12538
rect 15622 12484 15678 12486
rect 15702 12484 15758 12486
rect 15782 12484 15838 12486
rect 15862 12484 15918 12486
rect 15622 11450 15678 11452
rect 15702 11450 15758 11452
rect 15782 11450 15838 11452
rect 15862 11450 15918 11452
rect 15622 11398 15648 11450
rect 15648 11398 15678 11450
rect 15702 11398 15712 11450
rect 15712 11398 15758 11450
rect 15782 11398 15828 11450
rect 15828 11398 15838 11450
rect 15862 11398 15892 11450
rect 15892 11398 15918 11450
rect 15622 11396 15678 11398
rect 15702 11396 15758 11398
rect 15782 11396 15838 11398
rect 15862 11396 15918 11398
rect 15106 11056 15162 11112
rect 11956 6554 12012 6556
rect 12036 6554 12092 6556
rect 12116 6554 12172 6556
rect 12196 6554 12252 6556
rect 11956 6502 11982 6554
rect 11982 6502 12012 6554
rect 12036 6502 12046 6554
rect 12046 6502 12092 6554
rect 12116 6502 12162 6554
rect 12162 6502 12172 6554
rect 12196 6502 12226 6554
rect 12226 6502 12252 6554
rect 11956 6500 12012 6502
rect 12036 6500 12092 6502
rect 12116 6500 12172 6502
rect 12196 6500 12252 6502
rect 11956 5466 12012 5468
rect 12036 5466 12092 5468
rect 12116 5466 12172 5468
rect 12196 5466 12252 5468
rect 11956 5414 11982 5466
rect 11982 5414 12012 5466
rect 12036 5414 12046 5466
rect 12046 5414 12092 5466
rect 12116 5414 12162 5466
rect 12162 5414 12172 5466
rect 12196 5414 12226 5466
rect 12226 5414 12252 5466
rect 11956 5412 12012 5414
rect 12036 5412 12092 5414
rect 12116 5412 12172 5414
rect 12196 5412 12252 5414
rect 11956 4378 12012 4380
rect 12036 4378 12092 4380
rect 12116 4378 12172 4380
rect 12196 4378 12252 4380
rect 11956 4326 11982 4378
rect 11982 4326 12012 4378
rect 12036 4326 12046 4378
rect 12046 4326 12092 4378
rect 12116 4326 12162 4378
rect 12162 4326 12172 4378
rect 12196 4326 12226 4378
rect 12226 4326 12252 4378
rect 11956 4324 12012 4326
rect 12036 4324 12092 4326
rect 12116 4324 12172 4326
rect 12196 4324 12252 4326
rect 12162 3984 12218 4040
rect 11518 2488 11574 2544
rect 11956 3290 12012 3292
rect 12036 3290 12092 3292
rect 12116 3290 12172 3292
rect 12196 3290 12252 3292
rect 11956 3238 11982 3290
rect 11982 3238 12012 3290
rect 12036 3238 12046 3290
rect 12046 3238 12092 3290
rect 12116 3238 12162 3290
rect 12162 3238 12172 3290
rect 12196 3238 12226 3290
rect 12226 3238 12252 3290
rect 11956 3236 12012 3238
rect 12036 3236 12092 3238
rect 12116 3236 12172 3238
rect 12196 3236 12252 3238
rect 11956 2202 12012 2204
rect 12036 2202 12092 2204
rect 12116 2202 12172 2204
rect 12196 2202 12252 2204
rect 11956 2150 11982 2202
rect 11982 2150 12012 2202
rect 12036 2150 12046 2202
rect 12046 2150 12092 2202
rect 12116 2150 12162 2202
rect 12162 2150 12172 2202
rect 12196 2150 12226 2202
rect 12226 2150 12252 2202
rect 11956 2148 12012 2150
rect 12036 2148 12092 2150
rect 12116 2148 12172 2150
rect 12196 2148 12252 2150
rect 14002 4664 14058 4720
rect 15622 10362 15678 10364
rect 15702 10362 15758 10364
rect 15782 10362 15838 10364
rect 15862 10362 15918 10364
rect 15622 10310 15648 10362
rect 15648 10310 15678 10362
rect 15702 10310 15712 10362
rect 15712 10310 15758 10362
rect 15782 10310 15828 10362
rect 15828 10310 15838 10362
rect 15862 10310 15892 10362
rect 15892 10310 15918 10362
rect 15622 10308 15678 10310
rect 15702 10308 15758 10310
rect 15782 10308 15838 10310
rect 15862 10308 15918 10310
rect 19154 20440 19210 20496
rect 19062 18672 19118 18728
rect 17774 16768 17830 16824
rect 15622 9274 15678 9276
rect 15702 9274 15758 9276
rect 15782 9274 15838 9276
rect 15862 9274 15918 9276
rect 15622 9222 15648 9274
rect 15648 9222 15678 9274
rect 15702 9222 15712 9274
rect 15712 9222 15758 9274
rect 15782 9222 15828 9274
rect 15828 9222 15838 9274
rect 15862 9222 15892 9274
rect 15892 9222 15918 9274
rect 15622 9220 15678 9222
rect 15702 9220 15758 9222
rect 15782 9220 15838 9222
rect 15862 9220 15918 9222
rect 15622 8186 15678 8188
rect 15702 8186 15758 8188
rect 15782 8186 15838 8188
rect 15862 8186 15918 8188
rect 15622 8134 15648 8186
rect 15648 8134 15678 8186
rect 15702 8134 15712 8186
rect 15712 8134 15758 8186
rect 15782 8134 15828 8186
rect 15828 8134 15838 8186
rect 15862 8134 15892 8186
rect 15892 8134 15918 8186
rect 15622 8132 15678 8134
rect 15702 8132 15758 8134
rect 15782 8132 15838 8134
rect 15862 8132 15918 8134
rect 15622 7098 15678 7100
rect 15702 7098 15758 7100
rect 15782 7098 15838 7100
rect 15862 7098 15918 7100
rect 15622 7046 15648 7098
rect 15648 7046 15678 7098
rect 15702 7046 15712 7098
rect 15712 7046 15758 7098
rect 15782 7046 15828 7098
rect 15828 7046 15838 7098
rect 15862 7046 15892 7098
rect 15892 7046 15918 7098
rect 15622 7044 15678 7046
rect 15702 7044 15758 7046
rect 15782 7044 15838 7046
rect 15862 7044 15918 7046
rect 15622 6010 15678 6012
rect 15702 6010 15758 6012
rect 15782 6010 15838 6012
rect 15862 6010 15918 6012
rect 15622 5958 15648 6010
rect 15648 5958 15678 6010
rect 15702 5958 15712 6010
rect 15712 5958 15758 6010
rect 15782 5958 15828 6010
rect 15828 5958 15838 6010
rect 15862 5958 15892 6010
rect 15892 5958 15918 6010
rect 15622 5956 15678 5958
rect 15702 5956 15758 5958
rect 15782 5956 15838 5958
rect 15862 5956 15918 5958
rect 15198 3984 15254 4040
rect 15622 4922 15678 4924
rect 15702 4922 15758 4924
rect 15782 4922 15838 4924
rect 15862 4922 15918 4924
rect 15622 4870 15648 4922
rect 15648 4870 15678 4922
rect 15702 4870 15712 4922
rect 15712 4870 15758 4922
rect 15782 4870 15828 4922
rect 15828 4870 15838 4922
rect 15862 4870 15892 4922
rect 15892 4870 15918 4922
rect 15622 4868 15678 4870
rect 15702 4868 15758 4870
rect 15782 4868 15838 4870
rect 15862 4868 15918 4870
rect 15474 4800 15530 4856
rect 15622 3834 15678 3836
rect 15702 3834 15758 3836
rect 15782 3834 15838 3836
rect 15862 3834 15918 3836
rect 15622 3782 15648 3834
rect 15648 3782 15678 3834
rect 15702 3782 15712 3834
rect 15712 3782 15758 3834
rect 15782 3782 15828 3834
rect 15828 3782 15838 3834
rect 15862 3782 15892 3834
rect 15892 3782 15918 3834
rect 15622 3780 15678 3782
rect 15702 3780 15758 3782
rect 15782 3780 15838 3782
rect 15862 3780 15918 3782
rect 15622 2746 15678 2748
rect 15702 2746 15758 2748
rect 15782 2746 15838 2748
rect 15862 2746 15918 2748
rect 15622 2694 15648 2746
rect 15648 2694 15678 2746
rect 15702 2694 15712 2746
rect 15712 2694 15758 2746
rect 15782 2694 15828 2746
rect 15828 2694 15838 2746
rect 15862 2694 15892 2746
rect 15892 2694 15918 2746
rect 15622 2692 15678 2694
rect 15702 2692 15758 2694
rect 15782 2692 15838 2694
rect 15862 2692 15918 2694
rect 14922 2488 14978 2544
rect 15474 2488 15530 2544
rect 14830 1400 14886 1456
rect 16670 2624 16726 2680
rect 19289 19610 19345 19612
rect 19369 19610 19425 19612
rect 19449 19610 19505 19612
rect 19529 19610 19585 19612
rect 19289 19558 19315 19610
rect 19315 19558 19345 19610
rect 19369 19558 19379 19610
rect 19379 19558 19425 19610
rect 19449 19558 19495 19610
rect 19495 19558 19505 19610
rect 19529 19558 19559 19610
rect 19559 19558 19585 19610
rect 19289 19556 19345 19558
rect 19369 19556 19425 19558
rect 19449 19556 19505 19558
rect 19529 19556 19585 19558
rect 19289 18522 19345 18524
rect 19369 18522 19425 18524
rect 19449 18522 19505 18524
rect 19529 18522 19585 18524
rect 19289 18470 19315 18522
rect 19315 18470 19345 18522
rect 19369 18470 19379 18522
rect 19379 18470 19425 18522
rect 19449 18470 19495 18522
rect 19495 18470 19505 18522
rect 19529 18470 19559 18522
rect 19559 18470 19585 18522
rect 19289 18468 19345 18470
rect 19369 18468 19425 18470
rect 19449 18468 19505 18470
rect 19529 18468 19585 18470
rect 19289 17434 19345 17436
rect 19369 17434 19425 17436
rect 19449 17434 19505 17436
rect 19529 17434 19585 17436
rect 19289 17382 19315 17434
rect 19315 17382 19345 17434
rect 19369 17382 19379 17434
rect 19379 17382 19425 17434
rect 19449 17382 19495 17434
rect 19495 17382 19505 17434
rect 19529 17382 19559 17434
rect 19559 17382 19585 17434
rect 19289 17380 19345 17382
rect 19369 17380 19425 17382
rect 19449 17380 19505 17382
rect 19529 17380 19585 17382
rect 20074 16496 20130 16552
rect 19289 16346 19345 16348
rect 19369 16346 19425 16348
rect 19449 16346 19505 16348
rect 19529 16346 19585 16348
rect 19289 16294 19315 16346
rect 19315 16294 19345 16346
rect 19369 16294 19379 16346
rect 19379 16294 19425 16346
rect 19449 16294 19495 16346
rect 19495 16294 19505 16346
rect 19529 16294 19559 16346
rect 19559 16294 19585 16346
rect 19289 16292 19345 16294
rect 19369 16292 19425 16294
rect 19449 16292 19505 16294
rect 19529 16292 19585 16294
rect 19289 15258 19345 15260
rect 19369 15258 19425 15260
rect 19449 15258 19505 15260
rect 19529 15258 19585 15260
rect 19289 15206 19315 15258
rect 19315 15206 19345 15258
rect 19369 15206 19379 15258
rect 19379 15206 19425 15258
rect 19449 15206 19495 15258
rect 19495 15206 19505 15258
rect 19529 15206 19559 15258
rect 19559 15206 19585 15258
rect 19289 15204 19345 15206
rect 19369 15204 19425 15206
rect 19449 15204 19505 15206
rect 19529 15204 19585 15206
rect 19289 14170 19345 14172
rect 19369 14170 19425 14172
rect 19449 14170 19505 14172
rect 19529 14170 19585 14172
rect 19289 14118 19315 14170
rect 19315 14118 19345 14170
rect 19369 14118 19379 14170
rect 19379 14118 19425 14170
rect 19449 14118 19495 14170
rect 19495 14118 19505 14170
rect 19529 14118 19559 14170
rect 19559 14118 19585 14170
rect 19289 14116 19345 14118
rect 19369 14116 19425 14118
rect 19449 14116 19505 14118
rect 19529 14116 19585 14118
rect 19246 13504 19302 13560
rect 19289 13082 19345 13084
rect 19369 13082 19425 13084
rect 19449 13082 19505 13084
rect 19529 13082 19585 13084
rect 19289 13030 19315 13082
rect 19315 13030 19345 13082
rect 19369 13030 19379 13082
rect 19379 13030 19425 13082
rect 19449 13030 19495 13082
rect 19495 13030 19505 13082
rect 19529 13030 19559 13082
rect 19559 13030 19585 13082
rect 19289 13028 19345 13030
rect 19369 13028 19425 13030
rect 19449 13028 19505 13030
rect 19529 13028 19585 13030
rect 19289 11994 19345 11996
rect 19369 11994 19425 11996
rect 19449 11994 19505 11996
rect 19529 11994 19585 11996
rect 19289 11942 19315 11994
rect 19315 11942 19345 11994
rect 19369 11942 19379 11994
rect 19379 11942 19425 11994
rect 19449 11942 19495 11994
rect 19495 11942 19505 11994
rect 19529 11942 19559 11994
rect 19559 11942 19585 11994
rect 19289 11940 19345 11942
rect 19369 11940 19425 11942
rect 19449 11940 19505 11942
rect 19529 11940 19585 11942
rect 19338 11464 19394 11520
rect 19289 10906 19345 10908
rect 19369 10906 19425 10908
rect 19449 10906 19505 10908
rect 19529 10906 19585 10908
rect 19289 10854 19315 10906
rect 19315 10854 19345 10906
rect 19369 10854 19379 10906
rect 19379 10854 19425 10906
rect 19449 10854 19495 10906
rect 19495 10854 19505 10906
rect 19529 10854 19559 10906
rect 19559 10854 19585 10906
rect 19289 10852 19345 10854
rect 19369 10852 19425 10854
rect 19449 10852 19505 10854
rect 19529 10852 19585 10854
rect 21546 9968 21602 10024
rect 19289 9818 19345 9820
rect 19369 9818 19425 9820
rect 19449 9818 19505 9820
rect 19529 9818 19585 9820
rect 19289 9766 19315 9818
rect 19315 9766 19345 9818
rect 19369 9766 19379 9818
rect 19379 9766 19425 9818
rect 19449 9766 19495 9818
rect 19495 9766 19505 9818
rect 19529 9766 19559 9818
rect 19559 9766 19585 9818
rect 19289 9764 19345 9766
rect 19369 9764 19425 9766
rect 19449 9764 19505 9766
rect 19529 9764 19585 9766
rect 17866 8200 17922 8256
rect 18602 7948 18658 7984
rect 18602 7928 18604 7948
rect 18604 7928 18656 7948
rect 18656 7928 18658 7948
rect 17774 2352 17830 2408
rect 19289 8730 19345 8732
rect 19369 8730 19425 8732
rect 19449 8730 19505 8732
rect 19529 8730 19585 8732
rect 19289 8678 19315 8730
rect 19315 8678 19345 8730
rect 19369 8678 19379 8730
rect 19379 8678 19425 8730
rect 19449 8678 19495 8730
rect 19495 8678 19505 8730
rect 19529 8678 19559 8730
rect 19559 8678 19585 8730
rect 19289 8676 19345 8678
rect 19369 8676 19425 8678
rect 19449 8676 19505 8678
rect 19529 8676 19585 8678
rect 19289 7642 19345 7644
rect 19369 7642 19425 7644
rect 19449 7642 19505 7644
rect 19529 7642 19585 7644
rect 19289 7590 19315 7642
rect 19315 7590 19345 7642
rect 19369 7590 19379 7642
rect 19379 7590 19425 7642
rect 19449 7590 19495 7642
rect 19495 7590 19505 7642
rect 19529 7590 19559 7642
rect 19559 7590 19585 7642
rect 19289 7588 19345 7590
rect 19369 7588 19425 7590
rect 19449 7588 19505 7590
rect 19529 7588 19585 7590
rect 19154 6840 19210 6896
rect 19289 6554 19345 6556
rect 19369 6554 19425 6556
rect 19449 6554 19505 6556
rect 19529 6554 19585 6556
rect 19289 6502 19315 6554
rect 19315 6502 19345 6554
rect 19369 6502 19379 6554
rect 19379 6502 19425 6554
rect 19449 6502 19495 6554
rect 19495 6502 19505 6554
rect 19529 6502 19559 6554
rect 19559 6502 19585 6554
rect 19289 6500 19345 6502
rect 19369 6500 19425 6502
rect 19449 6500 19505 6502
rect 19529 6500 19585 6502
rect 19289 5466 19345 5468
rect 19369 5466 19425 5468
rect 19449 5466 19505 5468
rect 19529 5466 19585 5468
rect 19289 5414 19315 5466
rect 19315 5414 19345 5466
rect 19369 5414 19379 5466
rect 19379 5414 19425 5466
rect 19449 5414 19495 5466
rect 19495 5414 19505 5466
rect 19529 5414 19559 5466
rect 19559 5414 19585 5466
rect 19289 5412 19345 5414
rect 19369 5412 19425 5414
rect 19449 5412 19505 5414
rect 19529 5412 19585 5414
rect 18878 3984 18934 4040
rect 18694 2488 18750 2544
rect 18878 2624 18934 2680
rect 19289 4378 19345 4380
rect 19369 4378 19425 4380
rect 19449 4378 19505 4380
rect 19529 4378 19585 4380
rect 19289 4326 19315 4378
rect 19315 4326 19345 4378
rect 19369 4326 19379 4378
rect 19379 4326 19425 4378
rect 19449 4326 19495 4378
rect 19495 4326 19505 4378
rect 19529 4326 19559 4378
rect 19559 4326 19585 4378
rect 19289 4324 19345 4326
rect 19369 4324 19425 4326
rect 19449 4324 19505 4326
rect 19529 4324 19585 4326
rect 19798 5072 19854 5128
rect 19289 3290 19345 3292
rect 19369 3290 19425 3292
rect 19449 3290 19505 3292
rect 19529 3290 19585 3292
rect 19289 3238 19315 3290
rect 19315 3238 19345 3290
rect 19369 3238 19379 3290
rect 19379 3238 19425 3290
rect 19449 3238 19495 3290
rect 19495 3238 19505 3290
rect 19529 3238 19559 3290
rect 19559 3238 19585 3290
rect 19289 3236 19345 3238
rect 19369 3236 19425 3238
rect 19449 3236 19505 3238
rect 19529 3236 19585 3238
rect 19430 2488 19486 2544
rect 19289 2202 19345 2204
rect 19369 2202 19425 2204
rect 19449 2202 19505 2204
rect 19529 2202 19585 2204
rect 19289 2150 19315 2202
rect 19315 2150 19345 2202
rect 19369 2150 19379 2202
rect 19379 2150 19425 2202
rect 19449 2150 19495 2202
rect 19495 2150 19505 2202
rect 19529 2150 19559 2202
rect 19559 2150 19585 2202
rect 19289 2148 19345 2150
rect 19369 2148 19425 2150
rect 19449 2148 19505 2150
rect 19529 2148 19585 2150
rect 21546 2624 21602 2680
<< metal3 >>
rect 21520 20952 22000 21072
rect 0 20816 480 20936
rect 62 20362 122 20816
rect 19149 20498 19215 20501
rect 21590 20498 21650 20952
rect 19149 20496 21650 20498
rect 19149 20440 19154 20496
rect 19210 20440 21650 20496
rect 19149 20438 21650 20440
rect 19149 20435 19215 20438
rect 1577 20362 1643 20365
rect 62 20360 1643 20362
rect 62 20304 1582 20360
rect 1638 20304 1643 20360
rect 62 20302 1643 20304
rect 1577 20299 1643 20302
rect 4610 19616 4930 19617
rect 4610 19552 4618 19616
rect 4682 19552 4698 19616
rect 4762 19552 4778 19616
rect 4842 19552 4858 19616
rect 4922 19552 4930 19616
rect 4610 19551 4930 19552
rect 11944 19616 12264 19617
rect 11944 19552 11952 19616
rect 12016 19552 12032 19616
rect 12096 19552 12112 19616
rect 12176 19552 12192 19616
rect 12256 19552 12264 19616
rect 11944 19551 12264 19552
rect 19277 19616 19597 19617
rect 19277 19552 19285 19616
rect 19349 19552 19365 19616
rect 19429 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19597 19616
rect 19277 19551 19597 19552
rect 21520 19184 22000 19304
rect 8277 19072 8597 19073
rect 8277 19008 8285 19072
rect 8349 19008 8365 19072
rect 8429 19008 8445 19072
rect 8509 19008 8525 19072
rect 8589 19008 8597 19072
rect 8277 19007 8597 19008
rect 15610 19072 15930 19073
rect 15610 19008 15618 19072
rect 15682 19008 15698 19072
rect 15762 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15930 19072
rect 15610 19007 15930 19008
rect 0 18640 480 18760
rect 19057 18730 19123 18733
rect 21590 18730 21650 19184
rect 19057 18728 21650 18730
rect 19057 18672 19062 18728
rect 19118 18672 21650 18728
rect 19057 18670 21650 18672
rect 19057 18667 19123 18670
rect 62 18186 122 18640
rect 4610 18528 4930 18529
rect 4610 18464 4618 18528
rect 4682 18464 4698 18528
rect 4762 18464 4778 18528
rect 4842 18464 4858 18528
rect 4922 18464 4930 18528
rect 4610 18463 4930 18464
rect 11944 18528 12264 18529
rect 11944 18464 11952 18528
rect 12016 18464 12032 18528
rect 12096 18464 12112 18528
rect 12176 18464 12192 18528
rect 12256 18464 12264 18528
rect 11944 18463 12264 18464
rect 19277 18528 19597 18529
rect 19277 18464 19285 18528
rect 19349 18464 19365 18528
rect 19429 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19597 18528
rect 19277 18463 19597 18464
rect 1853 18186 1919 18189
rect 62 18184 1919 18186
rect 62 18128 1858 18184
rect 1914 18128 1919 18184
rect 62 18126 1919 18128
rect 1853 18123 1919 18126
rect 8277 17984 8597 17985
rect 8277 17920 8285 17984
rect 8349 17920 8365 17984
rect 8429 17920 8445 17984
rect 8509 17920 8525 17984
rect 8589 17920 8597 17984
rect 8277 17919 8597 17920
rect 15610 17984 15930 17985
rect 15610 17920 15618 17984
rect 15682 17920 15698 17984
rect 15762 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15930 17984
rect 15610 17919 15930 17920
rect 4610 17440 4930 17441
rect 4610 17376 4618 17440
rect 4682 17376 4698 17440
rect 4762 17376 4778 17440
rect 4842 17376 4858 17440
rect 4922 17376 4930 17440
rect 4610 17375 4930 17376
rect 11944 17440 12264 17441
rect 11944 17376 11952 17440
rect 12016 17376 12032 17440
rect 12096 17376 12112 17440
rect 12176 17376 12192 17440
rect 12256 17376 12264 17440
rect 11944 17375 12264 17376
rect 19277 17440 19597 17441
rect 19277 17376 19285 17440
rect 19349 17376 19365 17440
rect 19429 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19597 17440
rect 19277 17375 19597 17376
rect 21520 17280 22000 17400
rect 8277 16896 8597 16897
rect 8277 16832 8285 16896
rect 8349 16832 8365 16896
rect 8429 16832 8445 16896
rect 8509 16832 8525 16896
rect 8589 16832 8597 16896
rect 8277 16831 8597 16832
rect 15610 16896 15930 16897
rect 15610 16832 15618 16896
rect 15682 16832 15698 16896
rect 15762 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15930 16896
rect 15610 16831 15930 16832
rect 17769 16826 17835 16829
rect 21590 16826 21650 17280
rect 17769 16824 21650 16826
rect 17769 16768 17774 16824
rect 17830 16768 21650 16824
rect 17769 16766 21650 16768
rect 17769 16763 17835 16766
rect 0 16464 480 16584
rect 10317 16554 10383 16557
rect 20069 16554 20135 16557
rect 10317 16552 20135 16554
rect 10317 16496 10322 16552
rect 10378 16496 20074 16552
rect 20130 16496 20135 16552
rect 10317 16494 20135 16496
rect 10317 16491 10383 16494
rect 20069 16491 20135 16494
rect 62 16010 122 16464
rect 4610 16352 4930 16353
rect 4610 16288 4618 16352
rect 4682 16288 4698 16352
rect 4762 16288 4778 16352
rect 4842 16288 4858 16352
rect 4922 16288 4930 16352
rect 4610 16287 4930 16288
rect 11944 16352 12264 16353
rect 11944 16288 11952 16352
rect 12016 16288 12032 16352
rect 12096 16288 12112 16352
rect 12176 16288 12192 16352
rect 12256 16288 12264 16352
rect 11944 16287 12264 16288
rect 19277 16352 19597 16353
rect 19277 16288 19285 16352
rect 19349 16288 19365 16352
rect 19429 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19597 16352
rect 19277 16287 19597 16288
rect 1577 16010 1643 16013
rect 62 16008 1643 16010
rect 62 15952 1582 16008
rect 1638 15952 1643 16008
rect 62 15950 1643 15952
rect 1577 15947 1643 15950
rect 8277 15808 8597 15809
rect 8277 15744 8285 15808
rect 8349 15744 8365 15808
rect 8429 15744 8445 15808
rect 8509 15744 8525 15808
rect 8589 15744 8597 15808
rect 8277 15743 8597 15744
rect 15610 15808 15930 15809
rect 15610 15744 15618 15808
rect 15682 15744 15698 15808
rect 15762 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15930 15808
rect 15610 15743 15930 15744
rect 21520 15512 22000 15632
rect 4610 15264 4930 15265
rect 4610 15200 4618 15264
rect 4682 15200 4698 15264
rect 4762 15200 4778 15264
rect 4842 15200 4858 15264
rect 4922 15200 4930 15264
rect 4610 15199 4930 15200
rect 11944 15264 12264 15265
rect 11944 15200 11952 15264
rect 12016 15200 12032 15264
rect 12096 15200 12112 15264
rect 12176 15200 12192 15264
rect 12256 15200 12264 15264
rect 11944 15199 12264 15200
rect 19277 15264 19597 15265
rect 19277 15200 19285 15264
rect 19349 15200 19365 15264
rect 19429 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19597 15264
rect 19277 15199 19597 15200
rect 15101 15058 15167 15061
rect 21590 15058 21650 15512
rect 15101 15056 21650 15058
rect 15101 15000 15106 15056
rect 15162 15000 21650 15056
rect 15101 14998 21650 15000
rect 15101 14995 15167 14998
rect 8277 14720 8597 14721
rect 8277 14656 8285 14720
rect 8349 14656 8365 14720
rect 8429 14656 8445 14720
rect 8509 14656 8525 14720
rect 8589 14656 8597 14720
rect 8277 14655 8597 14656
rect 15610 14720 15930 14721
rect 15610 14656 15618 14720
rect 15682 14656 15698 14720
rect 15762 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15930 14720
rect 15610 14655 15930 14656
rect 0 14288 480 14408
rect 62 13834 122 14288
rect 4610 14176 4930 14177
rect 4610 14112 4618 14176
rect 4682 14112 4698 14176
rect 4762 14112 4778 14176
rect 4842 14112 4858 14176
rect 4922 14112 4930 14176
rect 4610 14111 4930 14112
rect 11944 14176 12264 14177
rect 11944 14112 11952 14176
rect 12016 14112 12032 14176
rect 12096 14112 12112 14176
rect 12176 14112 12192 14176
rect 12256 14112 12264 14176
rect 11944 14111 12264 14112
rect 19277 14176 19597 14177
rect 19277 14112 19285 14176
rect 19349 14112 19365 14176
rect 19429 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19597 14176
rect 19277 14111 19597 14112
rect 7966 13834 7972 13836
rect 62 13774 7972 13834
rect 7966 13772 7972 13774
rect 8036 13772 8042 13836
rect 21520 13700 22000 13728
rect 21520 13698 21588 13700
rect 21460 13638 21588 13698
rect 21520 13636 21588 13638
rect 21652 13636 22000 13700
rect 8277 13632 8597 13633
rect 8277 13568 8285 13632
rect 8349 13568 8365 13632
rect 8429 13568 8445 13632
rect 8509 13568 8525 13632
rect 8589 13568 8597 13632
rect 8277 13567 8597 13568
rect 15610 13632 15930 13633
rect 15610 13568 15618 13632
rect 15682 13568 15698 13632
rect 15762 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15930 13632
rect 21520 13608 22000 13636
rect 15610 13567 15930 13568
rect 19241 13562 19307 13565
rect 19241 13560 19350 13562
rect 19241 13504 19246 13560
rect 19302 13504 19350 13560
rect 19241 13499 19350 13504
rect 19290 13426 19350 13499
rect 21582 13426 21588 13428
rect 19290 13366 21588 13426
rect 21582 13364 21588 13366
rect 21652 13364 21658 13428
rect 4610 13088 4930 13089
rect 4610 13024 4618 13088
rect 4682 13024 4698 13088
rect 4762 13024 4778 13088
rect 4842 13024 4858 13088
rect 4922 13024 4930 13088
rect 4610 13023 4930 13024
rect 11944 13088 12264 13089
rect 11944 13024 11952 13088
rect 12016 13024 12032 13088
rect 12096 13024 12112 13088
rect 12176 13024 12192 13088
rect 12256 13024 12264 13088
rect 11944 13023 12264 13024
rect 19277 13088 19597 13089
rect 19277 13024 19285 13088
rect 19349 13024 19365 13088
rect 19429 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19597 13088
rect 19277 13023 19597 13024
rect 8277 12544 8597 12545
rect 8277 12480 8285 12544
rect 8349 12480 8365 12544
rect 8429 12480 8445 12544
rect 8509 12480 8525 12544
rect 8589 12480 8597 12544
rect 8277 12479 8597 12480
rect 15610 12544 15930 12545
rect 15610 12480 15618 12544
rect 15682 12480 15698 12544
rect 15762 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15930 12544
rect 15610 12479 15930 12480
rect 0 12112 480 12232
rect 62 11658 122 12112
rect 4610 12000 4930 12001
rect 4610 11936 4618 12000
rect 4682 11936 4698 12000
rect 4762 11936 4778 12000
rect 4842 11936 4858 12000
rect 4922 11936 4930 12000
rect 4610 11935 4930 11936
rect 11944 12000 12264 12001
rect 11944 11936 11952 12000
rect 12016 11936 12032 12000
rect 12096 11936 12112 12000
rect 12176 11936 12192 12000
rect 12256 11936 12264 12000
rect 11944 11935 12264 11936
rect 19277 12000 19597 12001
rect 19277 11936 19285 12000
rect 19349 11936 19365 12000
rect 19429 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19597 12000
rect 19277 11935 19597 11936
rect 21520 11840 22000 11960
rect 2037 11658 2103 11661
rect 62 11656 2103 11658
rect 62 11600 2042 11656
rect 2098 11600 2103 11656
rect 62 11598 2103 11600
rect 2037 11595 2103 11598
rect 19333 11522 19399 11525
rect 21590 11522 21650 11840
rect 19333 11520 21650 11522
rect 19333 11464 19338 11520
rect 19394 11464 21650 11520
rect 19333 11462 21650 11464
rect 19333 11459 19399 11462
rect 8277 11456 8597 11457
rect 8277 11392 8285 11456
rect 8349 11392 8365 11456
rect 8429 11392 8445 11456
rect 8509 11392 8525 11456
rect 8589 11392 8597 11456
rect 8277 11391 8597 11392
rect 15610 11456 15930 11457
rect 15610 11392 15618 11456
rect 15682 11392 15698 11456
rect 15762 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15930 11456
rect 15610 11391 15930 11392
rect 5257 11114 5323 11117
rect 15101 11114 15167 11117
rect 5257 11112 15167 11114
rect 5257 11056 5262 11112
rect 5318 11056 15106 11112
rect 15162 11056 15167 11112
rect 5257 11054 15167 11056
rect 5257 11051 5323 11054
rect 15101 11051 15167 11054
rect 4610 10912 4930 10913
rect 4610 10848 4618 10912
rect 4682 10848 4698 10912
rect 4762 10848 4778 10912
rect 4842 10848 4858 10912
rect 4922 10848 4930 10912
rect 4610 10847 4930 10848
rect 11944 10912 12264 10913
rect 11944 10848 11952 10912
rect 12016 10848 12032 10912
rect 12096 10848 12112 10912
rect 12176 10848 12192 10912
rect 12256 10848 12264 10912
rect 11944 10847 12264 10848
rect 19277 10912 19597 10913
rect 19277 10848 19285 10912
rect 19349 10848 19365 10912
rect 19429 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19597 10912
rect 19277 10847 19597 10848
rect 8277 10368 8597 10369
rect 8277 10304 8285 10368
rect 8349 10304 8365 10368
rect 8429 10304 8445 10368
rect 8509 10304 8525 10368
rect 8589 10304 8597 10368
rect 8277 10303 8597 10304
rect 15610 10368 15930 10369
rect 15610 10304 15618 10368
rect 15682 10304 15698 10368
rect 15762 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15930 10368
rect 15610 10303 15930 10304
rect 105 10162 171 10165
rect 9397 10162 9463 10165
rect 105 10160 9690 10162
rect 105 10104 110 10160
rect 166 10104 9402 10160
rect 9458 10104 9690 10160
rect 105 10102 9690 10104
rect 105 10099 171 10102
rect 9397 10099 9463 10102
rect 9630 10026 9690 10102
rect 10869 10026 10935 10029
rect 21520 10026 22000 10056
rect 9630 10024 10935 10026
rect 9630 9968 10874 10024
rect 10930 9968 10935 10024
rect 9630 9966 10935 9968
rect 21460 10024 22000 10026
rect 21460 9968 21546 10024
rect 21602 9968 22000 10024
rect 21460 9966 22000 9968
rect 10869 9963 10935 9966
rect 21520 9936 22000 9966
rect 0 9888 480 9920
rect 0 9832 110 9888
rect 166 9832 480 9888
rect 0 9800 480 9832
rect 4610 9824 4930 9825
rect 4610 9760 4618 9824
rect 4682 9760 4698 9824
rect 4762 9760 4778 9824
rect 4842 9760 4858 9824
rect 4922 9760 4930 9824
rect 4610 9759 4930 9760
rect 11944 9824 12264 9825
rect 11944 9760 11952 9824
rect 12016 9760 12032 9824
rect 12096 9760 12112 9824
rect 12176 9760 12192 9824
rect 12256 9760 12264 9824
rect 11944 9759 12264 9760
rect 19277 9824 19597 9825
rect 19277 9760 19285 9824
rect 19349 9760 19365 9824
rect 19429 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19597 9824
rect 19277 9759 19597 9760
rect 8277 9280 8597 9281
rect 8277 9216 8285 9280
rect 8349 9216 8365 9280
rect 8429 9216 8445 9280
rect 8509 9216 8525 9280
rect 8589 9216 8597 9280
rect 8277 9215 8597 9216
rect 15610 9280 15930 9281
rect 15610 9216 15618 9280
rect 15682 9216 15698 9280
rect 15762 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15930 9280
rect 15610 9215 15930 9216
rect 4610 8736 4930 8737
rect 4610 8672 4618 8736
rect 4682 8672 4698 8736
rect 4762 8672 4778 8736
rect 4842 8672 4858 8736
rect 4922 8672 4930 8736
rect 4610 8671 4930 8672
rect 11944 8736 12264 8737
rect 11944 8672 11952 8736
rect 12016 8672 12032 8736
rect 12096 8672 12112 8736
rect 12176 8672 12192 8736
rect 12256 8672 12264 8736
rect 11944 8671 12264 8672
rect 19277 8736 19597 8737
rect 19277 8672 19285 8736
rect 19349 8672 19365 8736
rect 19429 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19597 8736
rect 19277 8671 19597 8672
rect 7966 8468 7972 8532
rect 8036 8530 8042 8532
rect 9029 8530 9095 8533
rect 9254 8530 9260 8532
rect 8036 8528 9260 8530
rect 8036 8472 9034 8528
rect 9090 8472 9260 8528
rect 8036 8470 9260 8472
rect 8036 8468 8042 8470
rect 9029 8467 9095 8470
rect 9254 8468 9260 8470
rect 9324 8468 9330 8532
rect 17861 8258 17927 8261
rect 21520 8258 22000 8288
rect 17861 8256 22000 8258
rect 17861 8200 17866 8256
rect 17922 8200 22000 8256
rect 17861 8198 22000 8200
rect 17861 8195 17927 8198
rect 8277 8192 8597 8193
rect 8277 8128 8285 8192
rect 8349 8128 8365 8192
rect 8429 8128 8445 8192
rect 8509 8128 8525 8192
rect 8589 8128 8597 8192
rect 8277 8127 8597 8128
rect 15610 8192 15930 8193
rect 15610 8128 15618 8192
rect 15682 8128 15698 8192
rect 15762 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15930 8192
rect 21520 8168 22000 8198
rect 15610 8127 15930 8128
rect 54 7924 60 7988
rect 124 7986 130 7988
rect 6361 7986 6427 7989
rect 18597 7986 18663 7989
rect 124 7926 674 7986
rect 124 7924 130 7926
rect 614 7850 674 7926
rect 6361 7984 18663 7986
rect 6361 7928 6366 7984
rect 6422 7928 18602 7984
rect 18658 7928 18663 7984
rect 6361 7926 18663 7928
rect 6361 7923 6427 7926
rect 18597 7923 18663 7926
rect 10869 7850 10935 7853
rect 614 7848 10935 7850
rect 614 7792 10874 7848
rect 10930 7792 10935 7848
rect 614 7790 10935 7792
rect 10869 7787 10935 7790
rect 0 7716 480 7744
rect 0 7652 60 7716
rect 124 7652 480 7716
rect 0 7624 480 7652
rect 4610 7648 4930 7649
rect 4610 7584 4618 7648
rect 4682 7584 4698 7648
rect 4762 7584 4778 7648
rect 4842 7584 4858 7648
rect 4922 7584 4930 7648
rect 4610 7583 4930 7584
rect 11944 7648 12264 7649
rect 11944 7584 11952 7648
rect 12016 7584 12032 7648
rect 12096 7584 12112 7648
rect 12176 7584 12192 7648
rect 12256 7584 12264 7648
rect 11944 7583 12264 7584
rect 19277 7648 19597 7649
rect 19277 7584 19285 7648
rect 19349 7584 19365 7648
rect 19429 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19597 7648
rect 19277 7583 19597 7584
rect 8277 7104 8597 7105
rect 8277 7040 8285 7104
rect 8349 7040 8365 7104
rect 8429 7040 8445 7104
rect 8509 7040 8525 7104
rect 8589 7040 8597 7104
rect 8277 7039 8597 7040
rect 15610 7104 15930 7105
rect 15610 7040 15618 7104
rect 15682 7040 15698 7104
rect 15762 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15930 7104
rect 15610 7039 15930 7040
rect 19149 6898 19215 6901
rect 19149 6896 21650 6898
rect 19149 6840 19154 6896
rect 19210 6840 21650 6896
rect 19149 6838 21650 6840
rect 19149 6835 19215 6838
rect 4610 6560 4930 6561
rect 4610 6496 4618 6560
rect 4682 6496 4698 6560
rect 4762 6496 4778 6560
rect 4842 6496 4858 6560
rect 4922 6496 4930 6560
rect 4610 6495 4930 6496
rect 11944 6560 12264 6561
rect 11944 6496 11952 6560
rect 12016 6496 12032 6560
rect 12096 6496 12112 6560
rect 12176 6496 12192 6560
rect 12256 6496 12264 6560
rect 11944 6495 12264 6496
rect 19277 6560 19597 6561
rect 19277 6496 19285 6560
rect 19349 6496 19365 6560
rect 19429 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19597 6560
rect 19277 6495 19597 6496
rect 21590 6384 21650 6838
rect 21520 6264 22000 6384
rect 1393 6082 1459 6085
rect 62 6080 1459 6082
rect 62 6024 1398 6080
rect 1454 6024 1459 6080
rect 62 6022 1459 6024
rect 62 5568 122 6022
rect 1393 6019 1459 6022
rect 8277 6016 8597 6017
rect 8277 5952 8285 6016
rect 8349 5952 8365 6016
rect 8429 5952 8445 6016
rect 8509 5952 8525 6016
rect 8589 5952 8597 6016
rect 8277 5951 8597 5952
rect 15610 6016 15930 6017
rect 15610 5952 15618 6016
rect 15682 5952 15698 6016
rect 15762 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15930 6016
rect 15610 5951 15930 5952
rect 0 5448 480 5568
rect 4610 5472 4930 5473
rect 4610 5408 4618 5472
rect 4682 5408 4698 5472
rect 4762 5408 4778 5472
rect 4842 5408 4858 5472
rect 4922 5408 4930 5472
rect 4610 5407 4930 5408
rect 11944 5472 12264 5473
rect 11944 5408 11952 5472
rect 12016 5408 12032 5472
rect 12096 5408 12112 5472
rect 12176 5408 12192 5472
rect 12256 5408 12264 5472
rect 11944 5407 12264 5408
rect 19277 5472 19597 5473
rect 19277 5408 19285 5472
rect 19349 5408 19365 5472
rect 19429 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19597 5472
rect 19277 5407 19597 5408
rect 5349 5130 5415 5133
rect 9213 5130 9279 5133
rect 5349 5128 9279 5130
rect 5349 5072 5354 5128
rect 5410 5072 9218 5128
rect 9274 5072 9279 5128
rect 5349 5070 9279 5072
rect 5349 5067 5415 5070
rect 9213 5067 9279 5070
rect 19793 5130 19859 5133
rect 19793 5128 21650 5130
rect 19793 5072 19798 5128
rect 19854 5072 21650 5128
rect 19793 5070 21650 5072
rect 19793 5067 19859 5070
rect 8277 4928 8597 4929
rect 8277 4864 8285 4928
rect 8349 4864 8365 4928
rect 8429 4864 8445 4928
rect 8509 4864 8525 4928
rect 8589 4864 8597 4928
rect 8277 4863 8597 4864
rect 15610 4928 15930 4929
rect 15610 4864 15618 4928
rect 15682 4864 15698 4928
rect 15762 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15930 4928
rect 15610 4863 15930 4864
rect 9213 4858 9279 4861
rect 15469 4858 15535 4861
rect 9213 4856 15535 4858
rect 9213 4800 9218 4856
rect 9274 4800 15474 4856
rect 15530 4800 15535 4856
rect 9213 4798 15535 4800
rect 9213 4795 9279 4798
rect 15469 4795 15535 4798
rect 7557 4722 7623 4725
rect 13997 4722 14063 4725
rect 7557 4720 14063 4722
rect 7557 4664 7562 4720
rect 7618 4664 14002 4720
rect 14058 4664 14063 4720
rect 7557 4662 14063 4664
rect 7557 4659 7623 4662
rect 13997 4659 14063 4662
rect 21590 4616 21650 5070
rect 21520 4496 22000 4616
rect 4610 4384 4930 4385
rect 4610 4320 4618 4384
rect 4682 4320 4698 4384
rect 4762 4320 4778 4384
rect 4842 4320 4858 4384
rect 4922 4320 4930 4384
rect 4610 4319 4930 4320
rect 11944 4384 12264 4385
rect 11944 4320 11952 4384
rect 12016 4320 12032 4384
rect 12096 4320 12112 4384
rect 12176 4320 12192 4384
rect 12256 4320 12264 4384
rect 11944 4319 12264 4320
rect 19277 4384 19597 4385
rect 19277 4320 19285 4384
rect 19349 4320 19365 4384
rect 19429 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19597 4384
rect 19277 4319 19597 4320
rect 9254 3980 9260 4044
rect 9324 4042 9330 4044
rect 12157 4042 12223 4045
rect 9324 4040 12223 4042
rect 9324 3984 12162 4040
rect 12218 3984 12223 4040
rect 9324 3982 12223 3984
rect 9324 3980 9330 3982
rect 12157 3979 12223 3982
rect 15193 4042 15259 4045
rect 18873 4042 18939 4045
rect 15193 4040 18939 4042
rect 15193 3984 15198 4040
rect 15254 3984 18878 4040
rect 18934 3984 18939 4040
rect 15193 3982 18939 3984
rect 15193 3979 15259 3982
rect 18873 3979 18939 3982
rect 8277 3840 8597 3841
rect 8277 3776 8285 3840
rect 8349 3776 8365 3840
rect 8429 3776 8445 3840
rect 8509 3776 8525 3840
rect 8589 3776 8597 3840
rect 8277 3775 8597 3776
rect 15610 3840 15930 3841
rect 15610 3776 15618 3840
rect 15682 3776 15698 3840
rect 15762 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15930 3840
rect 15610 3775 15930 3776
rect 0 3360 480 3392
rect 0 3304 110 3360
rect 166 3304 480 3360
rect 0 3272 480 3304
rect 4610 3296 4930 3297
rect 4610 3232 4618 3296
rect 4682 3232 4698 3296
rect 4762 3232 4778 3296
rect 4842 3232 4858 3296
rect 4922 3232 4930 3296
rect 4610 3231 4930 3232
rect 11944 3296 12264 3297
rect 11944 3232 11952 3296
rect 12016 3232 12032 3296
rect 12096 3232 12112 3296
rect 12176 3232 12192 3296
rect 12256 3232 12264 3296
rect 11944 3231 12264 3232
rect 19277 3296 19597 3297
rect 19277 3232 19285 3296
rect 19349 3232 19365 3296
rect 19429 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19597 3296
rect 19277 3231 19597 3232
rect 8277 2752 8597 2753
rect 8277 2688 8285 2752
rect 8349 2688 8365 2752
rect 8429 2688 8445 2752
rect 8509 2688 8525 2752
rect 8589 2688 8597 2752
rect 8277 2687 8597 2688
rect 15610 2752 15930 2753
rect 15610 2688 15618 2752
rect 15682 2688 15698 2752
rect 15762 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15930 2752
rect 15610 2687 15930 2688
rect 16665 2682 16731 2685
rect 18873 2682 18939 2685
rect 21520 2682 22000 2712
rect 16665 2680 18939 2682
rect 16665 2624 16670 2680
rect 16726 2624 18878 2680
rect 18934 2624 18939 2680
rect 16665 2622 18939 2624
rect 21460 2680 22000 2682
rect 21460 2624 21546 2680
rect 21602 2624 22000 2680
rect 21460 2622 22000 2624
rect 16665 2619 16731 2622
rect 18873 2619 18939 2622
rect 21520 2592 22000 2622
rect 11513 2546 11579 2549
rect 14917 2546 14983 2549
rect 11513 2544 14983 2546
rect 11513 2488 11518 2544
rect 11574 2488 14922 2544
rect 14978 2488 14983 2544
rect 11513 2486 14983 2488
rect 11513 2483 11579 2486
rect 14917 2483 14983 2486
rect 15469 2546 15535 2549
rect 18689 2546 18755 2549
rect 19425 2546 19491 2549
rect 15469 2544 19491 2546
rect 15469 2488 15474 2544
rect 15530 2488 18694 2544
rect 18750 2488 19430 2544
rect 19486 2488 19491 2544
rect 15469 2486 19491 2488
rect 15469 2483 15535 2486
rect 18689 2483 18755 2486
rect 19425 2483 19491 2486
rect 5993 2410 6059 2413
rect 17769 2410 17835 2413
rect 5993 2408 17835 2410
rect 5993 2352 5998 2408
rect 6054 2352 17774 2408
rect 17830 2352 17835 2408
rect 5993 2350 17835 2352
rect 5993 2347 6059 2350
rect 17769 2347 17835 2350
rect 4610 2208 4930 2209
rect 4610 2144 4618 2208
rect 4682 2144 4698 2208
rect 4762 2144 4778 2208
rect 4842 2144 4858 2208
rect 4922 2144 4930 2208
rect 4610 2143 4930 2144
rect 11944 2208 12264 2209
rect 11944 2144 11952 2208
rect 12016 2144 12032 2208
rect 12096 2144 12112 2208
rect 12176 2144 12192 2208
rect 12256 2144 12264 2208
rect 11944 2143 12264 2144
rect 19277 2208 19597 2209
rect 19277 2144 19285 2208
rect 19349 2144 19365 2208
rect 19429 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19597 2208
rect 19277 2143 19597 2144
rect 4061 1730 4127 1733
rect 62 1728 4127 1730
rect 62 1672 4066 1728
rect 4122 1672 4127 1728
rect 62 1670 4127 1672
rect 62 1216 122 1670
rect 4061 1667 4127 1670
rect 14825 1458 14891 1461
rect 14825 1456 21650 1458
rect 14825 1400 14830 1456
rect 14886 1400 21650 1456
rect 14825 1398 21650 1400
rect 14825 1395 14891 1398
rect 0 1096 480 1216
rect 21590 944 21650 1398
rect 21520 824 22000 944
<< via3 >>
rect 4618 19612 4682 19616
rect 4618 19556 4622 19612
rect 4622 19556 4678 19612
rect 4678 19556 4682 19612
rect 4618 19552 4682 19556
rect 4698 19612 4762 19616
rect 4698 19556 4702 19612
rect 4702 19556 4758 19612
rect 4758 19556 4762 19612
rect 4698 19552 4762 19556
rect 4778 19612 4842 19616
rect 4778 19556 4782 19612
rect 4782 19556 4838 19612
rect 4838 19556 4842 19612
rect 4778 19552 4842 19556
rect 4858 19612 4922 19616
rect 4858 19556 4862 19612
rect 4862 19556 4918 19612
rect 4918 19556 4922 19612
rect 4858 19552 4922 19556
rect 11952 19612 12016 19616
rect 11952 19556 11956 19612
rect 11956 19556 12012 19612
rect 12012 19556 12016 19612
rect 11952 19552 12016 19556
rect 12032 19612 12096 19616
rect 12032 19556 12036 19612
rect 12036 19556 12092 19612
rect 12092 19556 12096 19612
rect 12032 19552 12096 19556
rect 12112 19612 12176 19616
rect 12112 19556 12116 19612
rect 12116 19556 12172 19612
rect 12172 19556 12176 19612
rect 12112 19552 12176 19556
rect 12192 19612 12256 19616
rect 12192 19556 12196 19612
rect 12196 19556 12252 19612
rect 12252 19556 12256 19612
rect 12192 19552 12256 19556
rect 19285 19612 19349 19616
rect 19285 19556 19289 19612
rect 19289 19556 19345 19612
rect 19345 19556 19349 19612
rect 19285 19552 19349 19556
rect 19365 19612 19429 19616
rect 19365 19556 19369 19612
rect 19369 19556 19425 19612
rect 19425 19556 19429 19612
rect 19365 19552 19429 19556
rect 19445 19612 19509 19616
rect 19445 19556 19449 19612
rect 19449 19556 19505 19612
rect 19505 19556 19509 19612
rect 19445 19552 19509 19556
rect 19525 19612 19589 19616
rect 19525 19556 19529 19612
rect 19529 19556 19585 19612
rect 19585 19556 19589 19612
rect 19525 19552 19589 19556
rect 8285 19068 8349 19072
rect 8285 19012 8289 19068
rect 8289 19012 8345 19068
rect 8345 19012 8349 19068
rect 8285 19008 8349 19012
rect 8365 19068 8429 19072
rect 8365 19012 8369 19068
rect 8369 19012 8425 19068
rect 8425 19012 8429 19068
rect 8365 19008 8429 19012
rect 8445 19068 8509 19072
rect 8445 19012 8449 19068
rect 8449 19012 8505 19068
rect 8505 19012 8509 19068
rect 8445 19008 8509 19012
rect 8525 19068 8589 19072
rect 8525 19012 8529 19068
rect 8529 19012 8585 19068
rect 8585 19012 8589 19068
rect 8525 19008 8589 19012
rect 15618 19068 15682 19072
rect 15618 19012 15622 19068
rect 15622 19012 15678 19068
rect 15678 19012 15682 19068
rect 15618 19008 15682 19012
rect 15698 19068 15762 19072
rect 15698 19012 15702 19068
rect 15702 19012 15758 19068
rect 15758 19012 15762 19068
rect 15698 19008 15762 19012
rect 15778 19068 15842 19072
rect 15778 19012 15782 19068
rect 15782 19012 15838 19068
rect 15838 19012 15842 19068
rect 15778 19008 15842 19012
rect 15858 19068 15922 19072
rect 15858 19012 15862 19068
rect 15862 19012 15918 19068
rect 15918 19012 15922 19068
rect 15858 19008 15922 19012
rect 4618 18524 4682 18528
rect 4618 18468 4622 18524
rect 4622 18468 4678 18524
rect 4678 18468 4682 18524
rect 4618 18464 4682 18468
rect 4698 18524 4762 18528
rect 4698 18468 4702 18524
rect 4702 18468 4758 18524
rect 4758 18468 4762 18524
rect 4698 18464 4762 18468
rect 4778 18524 4842 18528
rect 4778 18468 4782 18524
rect 4782 18468 4838 18524
rect 4838 18468 4842 18524
rect 4778 18464 4842 18468
rect 4858 18524 4922 18528
rect 4858 18468 4862 18524
rect 4862 18468 4918 18524
rect 4918 18468 4922 18524
rect 4858 18464 4922 18468
rect 11952 18524 12016 18528
rect 11952 18468 11956 18524
rect 11956 18468 12012 18524
rect 12012 18468 12016 18524
rect 11952 18464 12016 18468
rect 12032 18524 12096 18528
rect 12032 18468 12036 18524
rect 12036 18468 12092 18524
rect 12092 18468 12096 18524
rect 12032 18464 12096 18468
rect 12112 18524 12176 18528
rect 12112 18468 12116 18524
rect 12116 18468 12172 18524
rect 12172 18468 12176 18524
rect 12112 18464 12176 18468
rect 12192 18524 12256 18528
rect 12192 18468 12196 18524
rect 12196 18468 12252 18524
rect 12252 18468 12256 18524
rect 12192 18464 12256 18468
rect 19285 18524 19349 18528
rect 19285 18468 19289 18524
rect 19289 18468 19345 18524
rect 19345 18468 19349 18524
rect 19285 18464 19349 18468
rect 19365 18524 19429 18528
rect 19365 18468 19369 18524
rect 19369 18468 19425 18524
rect 19425 18468 19429 18524
rect 19365 18464 19429 18468
rect 19445 18524 19509 18528
rect 19445 18468 19449 18524
rect 19449 18468 19505 18524
rect 19505 18468 19509 18524
rect 19445 18464 19509 18468
rect 19525 18524 19589 18528
rect 19525 18468 19529 18524
rect 19529 18468 19585 18524
rect 19585 18468 19589 18524
rect 19525 18464 19589 18468
rect 8285 17980 8349 17984
rect 8285 17924 8289 17980
rect 8289 17924 8345 17980
rect 8345 17924 8349 17980
rect 8285 17920 8349 17924
rect 8365 17980 8429 17984
rect 8365 17924 8369 17980
rect 8369 17924 8425 17980
rect 8425 17924 8429 17980
rect 8365 17920 8429 17924
rect 8445 17980 8509 17984
rect 8445 17924 8449 17980
rect 8449 17924 8505 17980
rect 8505 17924 8509 17980
rect 8445 17920 8509 17924
rect 8525 17980 8589 17984
rect 8525 17924 8529 17980
rect 8529 17924 8585 17980
rect 8585 17924 8589 17980
rect 8525 17920 8589 17924
rect 15618 17980 15682 17984
rect 15618 17924 15622 17980
rect 15622 17924 15678 17980
rect 15678 17924 15682 17980
rect 15618 17920 15682 17924
rect 15698 17980 15762 17984
rect 15698 17924 15702 17980
rect 15702 17924 15758 17980
rect 15758 17924 15762 17980
rect 15698 17920 15762 17924
rect 15778 17980 15842 17984
rect 15778 17924 15782 17980
rect 15782 17924 15838 17980
rect 15838 17924 15842 17980
rect 15778 17920 15842 17924
rect 15858 17980 15922 17984
rect 15858 17924 15862 17980
rect 15862 17924 15918 17980
rect 15918 17924 15922 17980
rect 15858 17920 15922 17924
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 4698 17436 4762 17440
rect 4698 17380 4702 17436
rect 4702 17380 4758 17436
rect 4758 17380 4762 17436
rect 4698 17376 4762 17380
rect 4778 17436 4842 17440
rect 4778 17380 4782 17436
rect 4782 17380 4838 17436
rect 4838 17380 4842 17436
rect 4778 17376 4842 17380
rect 4858 17436 4922 17440
rect 4858 17380 4862 17436
rect 4862 17380 4918 17436
rect 4918 17380 4922 17436
rect 4858 17376 4922 17380
rect 11952 17436 12016 17440
rect 11952 17380 11956 17436
rect 11956 17380 12012 17436
rect 12012 17380 12016 17436
rect 11952 17376 12016 17380
rect 12032 17436 12096 17440
rect 12032 17380 12036 17436
rect 12036 17380 12092 17436
rect 12092 17380 12096 17436
rect 12032 17376 12096 17380
rect 12112 17436 12176 17440
rect 12112 17380 12116 17436
rect 12116 17380 12172 17436
rect 12172 17380 12176 17436
rect 12112 17376 12176 17380
rect 12192 17436 12256 17440
rect 12192 17380 12196 17436
rect 12196 17380 12252 17436
rect 12252 17380 12256 17436
rect 12192 17376 12256 17380
rect 19285 17436 19349 17440
rect 19285 17380 19289 17436
rect 19289 17380 19345 17436
rect 19345 17380 19349 17436
rect 19285 17376 19349 17380
rect 19365 17436 19429 17440
rect 19365 17380 19369 17436
rect 19369 17380 19425 17436
rect 19425 17380 19429 17436
rect 19365 17376 19429 17380
rect 19445 17436 19509 17440
rect 19445 17380 19449 17436
rect 19449 17380 19505 17436
rect 19505 17380 19509 17436
rect 19445 17376 19509 17380
rect 19525 17436 19589 17440
rect 19525 17380 19529 17436
rect 19529 17380 19585 17436
rect 19585 17380 19589 17436
rect 19525 17376 19589 17380
rect 8285 16892 8349 16896
rect 8285 16836 8289 16892
rect 8289 16836 8345 16892
rect 8345 16836 8349 16892
rect 8285 16832 8349 16836
rect 8365 16892 8429 16896
rect 8365 16836 8369 16892
rect 8369 16836 8425 16892
rect 8425 16836 8429 16892
rect 8365 16832 8429 16836
rect 8445 16892 8509 16896
rect 8445 16836 8449 16892
rect 8449 16836 8505 16892
rect 8505 16836 8509 16892
rect 8445 16832 8509 16836
rect 8525 16892 8589 16896
rect 8525 16836 8529 16892
rect 8529 16836 8585 16892
rect 8585 16836 8589 16892
rect 8525 16832 8589 16836
rect 15618 16892 15682 16896
rect 15618 16836 15622 16892
rect 15622 16836 15678 16892
rect 15678 16836 15682 16892
rect 15618 16832 15682 16836
rect 15698 16892 15762 16896
rect 15698 16836 15702 16892
rect 15702 16836 15758 16892
rect 15758 16836 15762 16892
rect 15698 16832 15762 16836
rect 15778 16892 15842 16896
rect 15778 16836 15782 16892
rect 15782 16836 15838 16892
rect 15838 16836 15842 16892
rect 15778 16832 15842 16836
rect 15858 16892 15922 16896
rect 15858 16836 15862 16892
rect 15862 16836 15918 16892
rect 15918 16836 15922 16892
rect 15858 16832 15922 16836
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 4698 16348 4762 16352
rect 4698 16292 4702 16348
rect 4702 16292 4758 16348
rect 4758 16292 4762 16348
rect 4698 16288 4762 16292
rect 4778 16348 4842 16352
rect 4778 16292 4782 16348
rect 4782 16292 4838 16348
rect 4838 16292 4842 16348
rect 4778 16288 4842 16292
rect 4858 16348 4922 16352
rect 4858 16292 4862 16348
rect 4862 16292 4918 16348
rect 4918 16292 4922 16348
rect 4858 16288 4922 16292
rect 11952 16348 12016 16352
rect 11952 16292 11956 16348
rect 11956 16292 12012 16348
rect 12012 16292 12016 16348
rect 11952 16288 12016 16292
rect 12032 16348 12096 16352
rect 12032 16292 12036 16348
rect 12036 16292 12092 16348
rect 12092 16292 12096 16348
rect 12032 16288 12096 16292
rect 12112 16348 12176 16352
rect 12112 16292 12116 16348
rect 12116 16292 12172 16348
rect 12172 16292 12176 16348
rect 12112 16288 12176 16292
rect 12192 16348 12256 16352
rect 12192 16292 12196 16348
rect 12196 16292 12252 16348
rect 12252 16292 12256 16348
rect 12192 16288 12256 16292
rect 19285 16348 19349 16352
rect 19285 16292 19289 16348
rect 19289 16292 19345 16348
rect 19345 16292 19349 16348
rect 19285 16288 19349 16292
rect 19365 16348 19429 16352
rect 19365 16292 19369 16348
rect 19369 16292 19425 16348
rect 19425 16292 19429 16348
rect 19365 16288 19429 16292
rect 19445 16348 19509 16352
rect 19445 16292 19449 16348
rect 19449 16292 19505 16348
rect 19505 16292 19509 16348
rect 19445 16288 19509 16292
rect 19525 16348 19589 16352
rect 19525 16292 19529 16348
rect 19529 16292 19585 16348
rect 19585 16292 19589 16348
rect 19525 16288 19589 16292
rect 8285 15804 8349 15808
rect 8285 15748 8289 15804
rect 8289 15748 8345 15804
rect 8345 15748 8349 15804
rect 8285 15744 8349 15748
rect 8365 15804 8429 15808
rect 8365 15748 8369 15804
rect 8369 15748 8425 15804
rect 8425 15748 8429 15804
rect 8365 15744 8429 15748
rect 8445 15804 8509 15808
rect 8445 15748 8449 15804
rect 8449 15748 8505 15804
rect 8505 15748 8509 15804
rect 8445 15744 8509 15748
rect 8525 15804 8589 15808
rect 8525 15748 8529 15804
rect 8529 15748 8585 15804
rect 8585 15748 8589 15804
rect 8525 15744 8589 15748
rect 15618 15804 15682 15808
rect 15618 15748 15622 15804
rect 15622 15748 15678 15804
rect 15678 15748 15682 15804
rect 15618 15744 15682 15748
rect 15698 15804 15762 15808
rect 15698 15748 15702 15804
rect 15702 15748 15758 15804
rect 15758 15748 15762 15804
rect 15698 15744 15762 15748
rect 15778 15804 15842 15808
rect 15778 15748 15782 15804
rect 15782 15748 15838 15804
rect 15838 15748 15842 15804
rect 15778 15744 15842 15748
rect 15858 15804 15922 15808
rect 15858 15748 15862 15804
rect 15862 15748 15918 15804
rect 15918 15748 15922 15804
rect 15858 15744 15922 15748
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 4698 15260 4762 15264
rect 4698 15204 4702 15260
rect 4702 15204 4758 15260
rect 4758 15204 4762 15260
rect 4698 15200 4762 15204
rect 4778 15260 4842 15264
rect 4778 15204 4782 15260
rect 4782 15204 4838 15260
rect 4838 15204 4842 15260
rect 4778 15200 4842 15204
rect 4858 15260 4922 15264
rect 4858 15204 4862 15260
rect 4862 15204 4918 15260
rect 4918 15204 4922 15260
rect 4858 15200 4922 15204
rect 11952 15260 12016 15264
rect 11952 15204 11956 15260
rect 11956 15204 12012 15260
rect 12012 15204 12016 15260
rect 11952 15200 12016 15204
rect 12032 15260 12096 15264
rect 12032 15204 12036 15260
rect 12036 15204 12092 15260
rect 12092 15204 12096 15260
rect 12032 15200 12096 15204
rect 12112 15260 12176 15264
rect 12112 15204 12116 15260
rect 12116 15204 12172 15260
rect 12172 15204 12176 15260
rect 12112 15200 12176 15204
rect 12192 15260 12256 15264
rect 12192 15204 12196 15260
rect 12196 15204 12252 15260
rect 12252 15204 12256 15260
rect 12192 15200 12256 15204
rect 19285 15260 19349 15264
rect 19285 15204 19289 15260
rect 19289 15204 19345 15260
rect 19345 15204 19349 15260
rect 19285 15200 19349 15204
rect 19365 15260 19429 15264
rect 19365 15204 19369 15260
rect 19369 15204 19425 15260
rect 19425 15204 19429 15260
rect 19365 15200 19429 15204
rect 19445 15260 19509 15264
rect 19445 15204 19449 15260
rect 19449 15204 19505 15260
rect 19505 15204 19509 15260
rect 19445 15200 19509 15204
rect 19525 15260 19589 15264
rect 19525 15204 19529 15260
rect 19529 15204 19585 15260
rect 19585 15204 19589 15260
rect 19525 15200 19589 15204
rect 8285 14716 8349 14720
rect 8285 14660 8289 14716
rect 8289 14660 8345 14716
rect 8345 14660 8349 14716
rect 8285 14656 8349 14660
rect 8365 14716 8429 14720
rect 8365 14660 8369 14716
rect 8369 14660 8425 14716
rect 8425 14660 8429 14716
rect 8365 14656 8429 14660
rect 8445 14716 8509 14720
rect 8445 14660 8449 14716
rect 8449 14660 8505 14716
rect 8505 14660 8509 14716
rect 8445 14656 8509 14660
rect 8525 14716 8589 14720
rect 8525 14660 8529 14716
rect 8529 14660 8585 14716
rect 8585 14660 8589 14716
rect 8525 14656 8589 14660
rect 15618 14716 15682 14720
rect 15618 14660 15622 14716
rect 15622 14660 15678 14716
rect 15678 14660 15682 14716
rect 15618 14656 15682 14660
rect 15698 14716 15762 14720
rect 15698 14660 15702 14716
rect 15702 14660 15758 14716
rect 15758 14660 15762 14716
rect 15698 14656 15762 14660
rect 15778 14716 15842 14720
rect 15778 14660 15782 14716
rect 15782 14660 15838 14716
rect 15838 14660 15842 14716
rect 15778 14656 15842 14660
rect 15858 14716 15922 14720
rect 15858 14660 15862 14716
rect 15862 14660 15918 14716
rect 15918 14660 15922 14716
rect 15858 14656 15922 14660
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 4698 14172 4762 14176
rect 4698 14116 4702 14172
rect 4702 14116 4758 14172
rect 4758 14116 4762 14172
rect 4698 14112 4762 14116
rect 4778 14172 4842 14176
rect 4778 14116 4782 14172
rect 4782 14116 4838 14172
rect 4838 14116 4842 14172
rect 4778 14112 4842 14116
rect 4858 14172 4922 14176
rect 4858 14116 4862 14172
rect 4862 14116 4918 14172
rect 4918 14116 4922 14172
rect 4858 14112 4922 14116
rect 11952 14172 12016 14176
rect 11952 14116 11956 14172
rect 11956 14116 12012 14172
rect 12012 14116 12016 14172
rect 11952 14112 12016 14116
rect 12032 14172 12096 14176
rect 12032 14116 12036 14172
rect 12036 14116 12092 14172
rect 12092 14116 12096 14172
rect 12032 14112 12096 14116
rect 12112 14172 12176 14176
rect 12112 14116 12116 14172
rect 12116 14116 12172 14172
rect 12172 14116 12176 14172
rect 12112 14112 12176 14116
rect 12192 14172 12256 14176
rect 12192 14116 12196 14172
rect 12196 14116 12252 14172
rect 12252 14116 12256 14172
rect 12192 14112 12256 14116
rect 19285 14172 19349 14176
rect 19285 14116 19289 14172
rect 19289 14116 19345 14172
rect 19345 14116 19349 14172
rect 19285 14112 19349 14116
rect 19365 14172 19429 14176
rect 19365 14116 19369 14172
rect 19369 14116 19425 14172
rect 19425 14116 19429 14172
rect 19365 14112 19429 14116
rect 19445 14172 19509 14176
rect 19445 14116 19449 14172
rect 19449 14116 19505 14172
rect 19505 14116 19509 14172
rect 19445 14112 19509 14116
rect 19525 14172 19589 14176
rect 19525 14116 19529 14172
rect 19529 14116 19585 14172
rect 19585 14116 19589 14172
rect 19525 14112 19589 14116
rect 7972 13772 8036 13836
rect 21588 13636 21652 13700
rect 8285 13628 8349 13632
rect 8285 13572 8289 13628
rect 8289 13572 8345 13628
rect 8345 13572 8349 13628
rect 8285 13568 8349 13572
rect 8365 13628 8429 13632
rect 8365 13572 8369 13628
rect 8369 13572 8425 13628
rect 8425 13572 8429 13628
rect 8365 13568 8429 13572
rect 8445 13628 8509 13632
rect 8445 13572 8449 13628
rect 8449 13572 8505 13628
rect 8505 13572 8509 13628
rect 8445 13568 8509 13572
rect 8525 13628 8589 13632
rect 8525 13572 8529 13628
rect 8529 13572 8585 13628
rect 8585 13572 8589 13628
rect 8525 13568 8589 13572
rect 15618 13628 15682 13632
rect 15618 13572 15622 13628
rect 15622 13572 15678 13628
rect 15678 13572 15682 13628
rect 15618 13568 15682 13572
rect 15698 13628 15762 13632
rect 15698 13572 15702 13628
rect 15702 13572 15758 13628
rect 15758 13572 15762 13628
rect 15698 13568 15762 13572
rect 15778 13628 15842 13632
rect 15778 13572 15782 13628
rect 15782 13572 15838 13628
rect 15838 13572 15842 13628
rect 15778 13568 15842 13572
rect 15858 13628 15922 13632
rect 15858 13572 15862 13628
rect 15862 13572 15918 13628
rect 15918 13572 15922 13628
rect 15858 13568 15922 13572
rect 21588 13364 21652 13428
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 4698 13084 4762 13088
rect 4698 13028 4702 13084
rect 4702 13028 4758 13084
rect 4758 13028 4762 13084
rect 4698 13024 4762 13028
rect 4778 13084 4842 13088
rect 4778 13028 4782 13084
rect 4782 13028 4838 13084
rect 4838 13028 4842 13084
rect 4778 13024 4842 13028
rect 4858 13084 4922 13088
rect 4858 13028 4862 13084
rect 4862 13028 4918 13084
rect 4918 13028 4922 13084
rect 4858 13024 4922 13028
rect 11952 13084 12016 13088
rect 11952 13028 11956 13084
rect 11956 13028 12012 13084
rect 12012 13028 12016 13084
rect 11952 13024 12016 13028
rect 12032 13084 12096 13088
rect 12032 13028 12036 13084
rect 12036 13028 12092 13084
rect 12092 13028 12096 13084
rect 12032 13024 12096 13028
rect 12112 13084 12176 13088
rect 12112 13028 12116 13084
rect 12116 13028 12172 13084
rect 12172 13028 12176 13084
rect 12112 13024 12176 13028
rect 12192 13084 12256 13088
rect 12192 13028 12196 13084
rect 12196 13028 12252 13084
rect 12252 13028 12256 13084
rect 12192 13024 12256 13028
rect 19285 13084 19349 13088
rect 19285 13028 19289 13084
rect 19289 13028 19345 13084
rect 19345 13028 19349 13084
rect 19285 13024 19349 13028
rect 19365 13084 19429 13088
rect 19365 13028 19369 13084
rect 19369 13028 19425 13084
rect 19425 13028 19429 13084
rect 19365 13024 19429 13028
rect 19445 13084 19509 13088
rect 19445 13028 19449 13084
rect 19449 13028 19505 13084
rect 19505 13028 19509 13084
rect 19445 13024 19509 13028
rect 19525 13084 19589 13088
rect 19525 13028 19529 13084
rect 19529 13028 19585 13084
rect 19585 13028 19589 13084
rect 19525 13024 19589 13028
rect 8285 12540 8349 12544
rect 8285 12484 8289 12540
rect 8289 12484 8345 12540
rect 8345 12484 8349 12540
rect 8285 12480 8349 12484
rect 8365 12540 8429 12544
rect 8365 12484 8369 12540
rect 8369 12484 8425 12540
rect 8425 12484 8429 12540
rect 8365 12480 8429 12484
rect 8445 12540 8509 12544
rect 8445 12484 8449 12540
rect 8449 12484 8505 12540
rect 8505 12484 8509 12540
rect 8445 12480 8509 12484
rect 8525 12540 8589 12544
rect 8525 12484 8529 12540
rect 8529 12484 8585 12540
rect 8585 12484 8589 12540
rect 8525 12480 8589 12484
rect 15618 12540 15682 12544
rect 15618 12484 15622 12540
rect 15622 12484 15678 12540
rect 15678 12484 15682 12540
rect 15618 12480 15682 12484
rect 15698 12540 15762 12544
rect 15698 12484 15702 12540
rect 15702 12484 15758 12540
rect 15758 12484 15762 12540
rect 15698 12480 15762 12484
rect 15778 12540 15842 12544
rect 15778 12484 15782 12540
rect 15782 12484 15838 12540
rect 15838 12484 15842 12540
rect 15778 12480 15842 12484
rect 15858 12540 15922 12544
rect 15858 12484 15862 12540
rect 15862 12484 15918 12540
rect 15918 12484 15922 12540
rect 15858 12480 15922 12484
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 4698 11996 4762 12000
rect 4698 11940 4702 11996
rect 4702 11940 4758 11996
rect 4758 11940 4762 11996
rect 4698 11936 4762 11940
rect 4778 11996 4842 12000
rect 4778 11940 4782 11996
rect 4782 11940 4838 11996
rect 4838 11940 4842 11996
rect 4778 11936 4842 11940
rect 4858 11996 4922 12000
rect 4858 11940 4862 11996
rect 4862 11940 4918 11996
rect 4918 11940 4922 11996
rect 4858 11936 4922 11940
rect 11952 11996 12016 12000
rect 11952 11940 11956 11996
rect 11956 11940 12012 11996
rect 12012 11940 12016 11996
rect 11952 11936 12016 11940
rect 12032 11996 12096 12000
rect 12032 11940 12036 11996
rect 12036 11940 12092 11996
rect 12092 11940 12096 11996
rect 12032 11936 12096 11940
rect 12112 11996 12176 12000
rect 12112 11940 12116 11996
rect 12116 11940 12172 11996
rect 12172 11940 12176 11996
rect 12112 11936 12176 11940
rect 12192 11996 12256 12000
rect 12192 11940 12196 11996
rect 12196 11940 12252 11996
rect 12252 11940 12256 11996
rect 12192 11936 12256 11940
rect 19285 11996 19349 12000
rect 19285 11940 19289 11996
rect 19289 11940 19345 11996
rect 19345 11940 19349 11996
rect 19285 11936 19349 11940
rect 19365 11996 19429 12000
rect 19365 11940 19369 11996
rect 19369 11940 19425 11996
rect 19425 11940 19429 11996
rect 19365 11936 19429 11940
rect 19445 11996 19509 12000
rect 19445 11940 19449 11996
rect 19449 11940 19505 11996
rect 19505 11940 19509 11996
rect 19445 11936 19509 11940
rect 19525 11996 19589 12000
rect 19525 11940 19529 11996
rect 19529 11940 19585 11996
rect 19585 11940 19589 11996
rect 19525 11936 19589 11940
rect 8285 11452 8349 11456
rect 8285 11396 8289 11452
rect 8289 11396 8345 11452
rect 8345 11396 8349 11452
rect 8285 11392 8349 11396
rect 8365 11452 8429 11456
rect 8365 11396 8369 11452
rect 8369 11396 8425 11452
rect 8425 11396 8429 11452
rect 8365 11392 8429 11396
rect 8445 11452 8509 11456
rect 8445 11396 8449 11452
rect 8449 11396 8505 11452
rect 8505 11396 8509 11452
rect 8445 11392 8509 11396
rect 8525 11452 8589 11456
rect 8525 11396 8529 11452
rect 8529 11396 8585 11452
rect 8585 11396 8589 11452
rect 8525 11392 8589 11396
rect 15618 11452 15682 11456
rect 15618 11396 15622 11452
rect 15622 11396 15678 11452
rect 15678 11396 15682 11452
rect 15618 11392 15682 11396
rect 15698 11452 15762 11456
rect 15698 11396 15702 11452
rect 15702 11396 15758 11452
rect 15758 11396 15762 11452
rect 15698 11392 15762 11396
rect 15778 11452 15842 11456
rect 15778 11396 15782 11452
rect 15782 11396 15838 11452
rect 15838 11396 15842 11452
rect 15778 11392 15842 11396
rect 15858 11452 15922 11456
rect 15858 11396 15862 11452
rect 15862 11396 15918 11452
rect 15918 11396 15922 11452
rect 15858 11392 15922 11396
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 4698 10908 4762 10912
rect 4698 10852 4702 10908
rect 4702 10852 4758 10908
rect 4758 10852 4762 10908
rect 4698 10848 4762 10852
rect 4778 10908 4842 10912
rect 4778 10852 4782 10908
rect 4782 10852 4838 10908
rect 4838 10852 4842 10908
rect 4778 10848 4842 10852
rect 4858 10908 4922 10912
rect 4858 10852 4862 10908
rect 4862 10852 4918 10908
rect 4918 10852 4922 10908
rect 4858 10848 4922 10852
rect 11952 10908 12016 10912
rect 11952 10852 11956 10908
rect 11956 10852 12012 10908
rect 12012 10852 12016 10908
rect 11952 10848 12016 10852
rect 12032 10908 12096 10912
rect 12032 10852 12036 10908
rect 12036 10852 12092 10908
rect 12092 10852 12096 10908
rect 12032 10848 12096 10852
rect 12112 10908 12176 10912
rect 12112 10852 12116 10908
rect 12116 10852 12172 10908
rect 12172 10852 12176 10908
rect 12112 10848 12176 10852
rect 12192 10908 12256 10912
rect 12192 10852 12196 10908
rect 12196 10852 12252 10908
rect 12252 10852 12256 10908
rect 12192 10848 12256 10852
rect 19285 10908 19349 10912
rect 19285 10852 19289 10908
rect 19289 10852 19345 10908
rect 19345 10852 19349 10908
rect 19285 10848 19349 10852
rect 19365 10908 19429 10912
rect 19365 10852 19369 10908
rect 19369 10852 19425 10908
rect 19425 10852 19429 10908
rect 19365 10848 19429 10852
rect 19445 10908 19509 10912
rect 19445 10852 19449 10908
rect 19449 10852 19505 10908
rect 19505 10852 19509 10908
rect 19445 10848 19509 10852
rect 19525 10908 19589 10912
rect 19525 10852 19529 10908
rect 19529 10852 19585 10908
rect 19585 10852 19589 10908
rect 19525 10848 19589 10852
rect 8285 10364 8349 10368
rect 8285 10308 8289 10364
rect 8289 10308 8345 10364
rect 8345 10308 8349 10364
rect 8285 10304 8349 10308
rect 8365 10364 8429 10368
rect 8365 10308 8369 10364
rect 8369 10308 8425 10364
rect 8425 10308 8429 10364
rect 8365 10304 8429 10308
rect 8445 10364 8509 10368
rect 8445 10308 8449 10364
rect 8449 10308 8505 10364
rect 8505 10308 8509 10364
rect 8445 10304 8509 10308
rect 8525 10364 8589 10368
rect 8525 10308 8529 10364
rect 8529 10308 8585 10364
rect 8585 10308 8589 10364
rect 8525 10304 8589 10308
rect 15618 10364 15682 10368
rect 15618 10308 15622 10364
rect 15622 10308 15678 10364
rect 15678 10308 15682 10364
rect 15618 10304 15682 10308
rect 15698 10364 15762 10368
rect 15698 10308 15702 10364
rect 15702 10308 15758 10364
rect 15758 10308 15762 10364
rect 15698 10304 15762 10308
rect 15778 10364 15842 10368
rect 15778 10308 15782 10364
rect 15782 10308 15838 10364
rect 15838 10308 15842 10364
rect 15778 10304 15842 10308
rect 15858 10364 15922 10368
rect 15858 10308 15862 10364
rect 15862 10308 15918 10364
rect 15918 10308 15922 10364
rect 15858 10304 15922 10308
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 4698 9820 4762 9824
rect 4698 9764 4702 9820
rect 4702 9764 4758 9820
rect 4758 9764 4762 9820
rect 4698 9760 4762 9764
rect 4778 9820 4842 9824
rect 4778 9764 4782 9820
rect 4782 9764 4838 9820
rect 4838 9764 4842 9820
rect 4778 9760 4842 9764
rect 4858 9820 4922 9824
rect 4858 9764 4862 9820
rect 4862 9764 4918 9820
rect 4918 9764 4922 9820
rect 4858 9760 4922 9764
rect 11952 9820 12016 9824
rect 11952 9764 11956 9820
rect 11956 9764 12012 9820
rect 12012 9764 12016 9820
rect 11952 9760 12016 9764
rect 12032 9820 12096 9824
rect 12032 9764 12036 9820
rect 12036 9764 12092 9820
rect 12092 9764 12096 9820
rect 12032 9760 12096 9764
rect 12112 9820 12176 9824
rect 12112 9764 12116 9820
rect 12116 9764 12172 9820
rect 12172 9764 12176 9820
rect 12112 9760 12176 9764
rect 12192 9820 12256 9824
rect 12192 9764 12196 9820
rect 12196 9764 12252 9820
rect 12252 9764 12256 9820
rect 12192 9760 12256 9764
rect 19285 9820 19349 9824
rect 19285 9764 19289 9820
rect 19289 9764 19345 9820
rect 19345 9764 19349 9820
rect 19285 9760 19349 9764
rect 19365 9820 19429 9824
rect 19365 9764 19369 9820
rect 19369 9764 19425 9820
rect 19425 9764 19429 9820
rect 19365 9760 19429 9764
rect 19445 9820 19509 9824
rect 19445 9764 19449 9820
rect 19449 9764 19505 9820
rect 19505 9764 19509 9820
rect 19445 9760 19509 9764
rect 19525 9820 19589 9824
rect 19525 9764 19529 9820
rect 19529 9764 19585 9820
rect 19585 9764 19589 9820
rect 19525 9760 19589 9764
rect 8285 9276 8349 9280
rect 8285 9220 8289 9276
rect 8289 9220 8345 9276
rect 8345 9220 8349 9276
rect 8285 9216 8349 9220
rect 8365 9276 8429 9280
rect 8365 9220 8369 9276
rect 8369 9220 8425 9276
rect 8425 9220 8429 9276
rect 8365 9216 8429 9220
rect 8445 9276 8509 9280
rect 8445 9220 8449 9276
rect 8449 9220 8505 9276
rect 8505 9220 8509 9276
rect 8445 9216 8509 9220
rect 8525 9276 8589 9280
rect 8525 9220 8529 9276
rect 8529 9220 8585 9276
rect 8585 9220 8589 9276
rect 8525 9216 8589 9220
rect 15618 9276 15682 9280
rect 15618 9220 15622 9276
rect 15622 9220 15678 9276
rect 15678 9220 15682 9276
rect 15618 9216 15682 9220
rect 15698 9276 15762 9280
rect 15698 9220 15702 9276
rect 15702 9220 15758 9276
rect 15758 9220 15762 9276
rect 15698 9216 15762 9220
rect 15778 9276 15842 9280
rect 15778 9220 15782 9276
rect 15782 9220 15838 9276
rect 15838 9220 15842 9276
rect 15778 9216 15842 9220
rect 15858 9276 15922 9280
rect 15858 9220 15862 9276
rect 15862 9220 15918 9276
rect 15918 9220 15922 9276
rect 15858 9216 15922 9220
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 4698 8732 4762 8736
rect 4698 8676 4702 8732
rect 4702 8676 4758 8732
rect 4758 8676 4762 8732
rect 4698 8672 4762 8676
rect 4778 8732 4842 8736
rect 4778 8676 4782 8732
rect 4782 8676 4838 8732
rect 4838 8676 4842 8732
rect 4778 8672 4842 8676
rect 4858 8732 4922 8736
rect 4858 8676 4862 8732
rect 4862 8676 4918 8732
rect 4918 8676 4922 8732
rect 4858 8672 4922 8676
rect 11952 8732 12016 8736
rect 11952 8676 11956 8732
rect 11956 8676 12012 8732
rect 12012 8676 12016 8732
rect 11952 8672 12016 8676
rect 12032 8732 12096 8736
rect 12032 8676 12036 8732
rect 12036 8676 12092 8732
rect 12092 8676 12096 8732
rect 12032 8672 12096 8676
rect 12112 8732 12176 8736
rect 12112 8676 12116 8732
rect 12116 8676 12172 8732
rect 12172 8676 12176 8732
rect 12112 8672 12176 8676
rect 12192 8732 12256 8736
rect 12192 8676 12196 8732
rect 12196 8676 12252 8732
rect 12252 8676 12256 8732
rect 12192 8672 12256 8676
rect 19285 8732 19349 8736
rect 19285 8676 19289 8732
rect 19289 8676 19345 8732
rect 19345 8676 19349 8732
rect 19285 8672 19349 8676
rect 19365 8732 19429 8736
rect 19365 8676 19369 8732
rect 19369 8676 19425 8732
rect 19425 8676 19429 8732
rect 19365 8672 19429 8676
rect 19445 8732 19509 8736
rect 19445 8676 19449 8732
rect 19449 8676 19505 8732
rect 19505 8676 19509 8732
rect 19445 8672 19509 8676
rect 19525 8732 19589 8736
rect 19525 8676 19529 8732
rect 19529 8676 19585 8732
rect 19585 8676 19589 8732
rect 19525 8672 19589 8676
rect 7972 8468 8036 8532
rect 9260 8468 9324 8532
rect 8285 8188 8349 8192
rect 8285 8132 8289 8188
rect 8289 8132 8345 8188
rect 8345 8132 8349 8188
rect 8285 8128 8349 8132
rect 8365 8188 8429 8192
rect 8365 8132 8369 8188
rect 8369 8132 8425 8188
rect 8425 8132 8429 8188
rect 8365 8128 8429 8132
rect 8445 8188 8509 8192
rect 8445 8132 8449 8188
rect 8449 8132 8505 8188
rect 8505 8132 8509 8188
rect 8445 8128 8509 8132
rect 8525 8188 8589 8192
rect 8525 8132 8529 8188
rect 8529 8132 8585 8188
rect 8585 8132 8589 8188
rect 8525 8128 8589 8132
rect 15618 8188 15682 8192
rect 15618 8132 15622 8188
rect 15622 8132 15678 8188
rect 15678 8132 15682 8188
rect 15618 8128 15682 8132
rect 15698 8188 15762 8192
rect 15698 8132 15702 8188
rect 15702 8132 15758 8188
rect 15758 8132 15762 8188
rect 15698 8128 15762 8132
rect 15778 8188 15842 8192
rect 15778 8132 15782 8188
rect 15782 8132 15838 8188
rect 15838 8132 15842 8188
rect 15778 8128 15842 8132
rect 15858 8188 15922 8192
rect 15858 8132 15862 8188
rect 15862 8132 15918 8188
rect 15918 8132 15922 8188
rect 15858 8128 15922 8132
rect 60 7924 124 7988
rect 60 7652 124 7716
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 4698 7644 4762 7648
rect 4698 7588 4702 7644
rect 4702 7588 4758 7644
rect 4758 7588 4762 7644
rect 4698 7584 4762 7588
rect 4778 7644 4842 7648
rect 4778 7588 4782 7644
rect 4782 7588 4838 7644
rect 4838 7588 4842 7644
rect 4778 7584 4842 7588
rect 4858 7644 4922 7648
rect 4858 7588 4862 7644
rect 4862 7588 4918 7644
rect 4918 7588 4922 7644
rect 4858 7584 4922 7588
rect 11952 7644 12016 7648
rect 11952 7588 11956 7644
rect 11956 7588 12012 7644
rect 12012 7588 12016 7644
rect 11952 7584 12016 7588
rect 12032 7644 12096 7648
rect 12032 7588 12036 7644
rect 12036 7588 12092 7644
rect 12092 7588 12096 7644
rect 12032 7584 12096 7588
rect 12112 7644 12176 7648
rect 12112 7588 12116 7644
rect 12116 7588 12172 7644
rect 12172 7588 12176 7644
rect 12112 7584 12176 7588
rect 12192 7644 12256 7648
rect 12192 7588 12196 7644
rect 12196 7588 12252 7644
rect 12252 7588 12256 7644
rect 12192 7584 12256 7588
rect 19285 7644 19349 7648
rect 19285 7588 19289 7644
rect 19289 7588 19345 7644
rect 19345 7588 19349 7644
rect 19285 7584 19349 7588
rect 19365 7644 19429 7648
rect 19365 7588 19369 7644
rect 19369 7588 19425 7644
rect 19425 7588 19429 7644
rect 19365 7584 19429 7588
rect 19445 7644 19509 7648
rect 19445 7588 19449 7644
rect 19449 7588 19505 7644
rect 19505 7588 19509 7644
rect 19445 7584 19509 7588
rect 19525 7644 19589 7648
rect 19525 7588 19529 7644
rect 19529 7588 19585 7644
rect 19585 7588 19589 7644
rect 19525 7584 19589 7588
rect 8285 7100 8349 7104
rect 8285 7044 8289 7100
rect 8289 7044 8345 7100
rect 8345 7044 8349 7100
rect 8285 7040 8349 7044
rect 8365 7100 8429 7104
rect 8365 7044 8369 7100
rect 8369 7044 8425 7100
rect 8425 7044 8429 7100
rect 8365 7040 8429 7044
rect 8445 7100 8509 7104
rect 8445 7044 8449 7100
rect 8449 7044 8505 7100
rect 8505 7044 8509 7100
rect 8445 7040 8509 7044
rect 8525 7100 8589 7104
rect 8525 7044 8529 7100
rect 8529 7044 8585 7100
rect 8585 7044 8589 7100
rect 8525 7040 8589 7044
rect 15618 7100 15682 7104
rect 15618 7044 15622 7100
rect 15622 7044 15678 7100
rect 15678 7044 15682 7100
rect 15618 7040 15682 7044
rect 15698 7100 15762 7104
rect 15698 7044 15702 7100
rect 15702 7044 15758 7100
rect 15758 7044 15762 7100
rect 15698 7040 15762 7044
rect 15778 7100 15842 7104
rect 15778 7044 15782 7100
rect 15782 7044 15838 7100
rect 15838 7044 15842 7100
rect 15778 7040 15842 7044
rect 15858 7100 15922 7104
rect 15858 7044 15862 7100
rect 15862 7044 15918 7100
rect 15918 7044 15922 7100
rect 15858 7040 15922 7044
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 4698 6556 4762 6560
rect 4698 6500 4702 6556
rect 4702 6500 4758 6556
rect 4758 6500 4762 6556
rect 4698 6496 4762 6500
rect 4778 6556 4842 6560
rect 4778 6500 4782 6556
rect 4782 6500 4838 6556
rect 4838 6500 4842 6556
rect 4778 6496 4842 6500
rect 4858 6556 4922 6560
rect 4858 6500 4862 6556
rect 4862 6500 4918 6556
rect 4918 6500 4922 6556
rect 4858 6496 4922 6500
rect 11952 6556 12016 6560
rect 11952 6500 11956 6556
rect 11956 6500 12012 6556
rect 12012 6500 12016 6556
rect 11952 6496 12016 6500
rect 12032 6556 12096 6560
rect 12032 6500 12036 6556
rect 12036 6500 12092 6556
rect 12092 6500 12096 6556
rect 12032 6496 12096 6500
rect 12112 6556 12176 6560
rect 12112 6500 12116 6556
rect 12116 6500 12172 6556
rect 12172 6500 12176 6556
rect 12112 6496 12176 6500
rect 12192 6556 12256 6560
rect 12192 6500 12196 6556
rect 12196 6500 12252 6556
rect 12252 6500 12256 6556
rect 12192 6496 12256 6500
rect 19285 6556 19349 6560
rect 19285 6500 19289 6556
rect 19289 6500 19345 6556
rect 19345 6500 19349 6556
rect 19285 6496 19349 6500
rect 19365 6556 19429 6560
rect 19365 6500 19369 6556
rect 19369 6500 19425 6556
rect 19425 6500 19429 6556
rect 19365 6496 19429 6500
rect 19445 6556 19509 6560
rect 19445 6500 19449 6556
rect 19449 6500 19505 6556
rect 19505 6500 19509 6556
rect 19445 6496 19509 6500
rect 19525 6556 19589 6560
rect 19525 6500 19529 6556
rect 19529 6500 19585 6556
rect 19585 6500 19589 6556
rect 19525 6496 19589 6500
rect 8285 6012 8349 6016
rect 8285 5956 8289 6012
rect 8289 5956 8345 6012
rect 8345 5956 8349 6012
rect 8285 5952 8349 5956
rect 8365 6012 8429 6016
rect 8365 5956 8369 6012
rect 8369 5956 8425 6012
rect 8425 5956 8429 6012
rect 8365 5952 8429 5956
rect 8445 6012 8509 6016
rect 8445 5956 8449 6012
rect 8449 5956 8505 6012
rect 8505 5956 8509 6012
rect 8445 5952 8509 5956
rect 8525 6012 8589 6016
rect 8525 5956 8529 6012
rect 8529 5956 8585 6012
rect 8585 5956 8589 6012
rect 8525 5952 8589 5956
rect 15618 6012 15682 6016
rect 15618 5956 15622 6012
rect 15622 5956 15678 6012
rect 15678 5956 15682 6012
rect 15618 5952 15682 5956
rect 15698 6012 15762 6016
rect 15698 5956 15702 6012
rect 15702 5956 15758 6012
rect 15758 5956 15762 6012
rect 15698 5952 15762 5956
rect 15778 6012 15842 6016
rect 15778 5956 15782 6012
rect 15782 5956 15838 6012
rect 15838 5956 15842 6012
rect 15778 5952 15842 5956
rect 15858 6012 15922 6016
rect 15858 5956 15862 6012
rect 15862 5956 15918 6012
rect 15918 5956 15922 6012
rect 15858 5952 15922 5956
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 4698 5468 4762 5472
rect 4698 5412 4702 5468
rect 4702 5412 4758 5468
rect 4758 5412 4762 5468
rect 4698 5408 4762 5412
rect 4778 5468 4842 5472
rect 4778 5412 4782 5468
rect 4782 5412 4838 5468
rect 4838 5412 4842 5468
rect 4778 5408 4842 5412
rect 4858 5468 4922 5472
rect 4858 5412 4862 5468
rect 4862 5412 4918 5468
rect 4918 5412 4922 5468
rect 4858 5408 4922 5412
rect 11952 5468 12016 5472
rect 11952 5412 11956 5468
rect 11956 5412 12012 5468
rect 12012 5412 12016 5468
rect 11952 5408 12016 5412
rect 12032 5468 12096 5472
rect 12032 5412 12036 5468
rect 12036 5412 12092 5468
rect 12092 5412 12096 5468
rect 12032 5408 12096 5412
rect 12112 5468 12176 5472
rect 12112 5412 12116 5468
rect 12116 5412 12172 5468
rect 12172 5412 12176 5468
rect 12112 5408 12176 5412
rect 12192 5468 12256 5472
rect 12192 5412 12196 5468
rect 12196 5412 12252 5468
rect 12252 5412 12256 5468
rect 12192 5408 12256 5412
rect 19285 5468 19349 5472
rect 19285 5412 19289 5468
rect 19289 5412 19345 5468
rect 19345 5412 19349 5468
rect 19285 5408 19349 5412
rect 19365 5468 19429 5472
rect 19365 5412 19369 5468
rect 19369 5412 19425 5468
rect 19425 5412 19429 5468
rect 19365 5408 19429 5412
rect 19445 5468 19509 5472
rect 19445 5412 19449 5468
rect 19449 5412 19505 5468
rect 19505 5412 19509 5468
rect 19445 5408 19509 5412
rect 19525 5468 19589 5472
rect 19525 5412 19529 5468
rect 19529 5412 19585 5468
rect 19585 5412 19589 5468
rect 19525 5408 19589 5412
rect 8285 4924 8349 4928
rect 8285 4868 8289 4924
rect 8289 4868 8345 4924
rect 8345 4868 8349 4924
rect 8285 4864 8349 4868
rect 8365 4924 8429 4928
rect 8365 4868 8369 4924
rect 8369 4868 8425 4924
rect 8425 4868 8429 4924
rect 8365 4864 8429 4868
rect 8445 4924 8509 4928
rect 8445 4868 8449 4924
rect 8449 4868 8505 4924
rect 8505 4868 8509 4924
rect 8445 4864 8509 4868
rect 8525 4924 8589 4928
rect 8525 4868 8529 4924
rect 8529 4868 8585 4924
rect 8585 4868 8589 4924
rect 8525 4864 8589 4868
rect 15618 4924 15682 4928
rect 15618 4868 15622 4924
rect 15622 4868 15678 4924
rect 15678 4868 15682 4924
rect 15618 4864 15682 4868
rect 15698 4924 15762 4928
rect 15698 4868 15702 4924
rect 15702 4868 15758 4924
rect 15758 4868 15762 4924
rect 15698 4864 15762 4868
rect 15778 4924 15842 4928
rect 15778 4868 15782 4924
rect 15782 4868 15838 4924
rect 15838 4868 15842 4924
rect 15778 4864 15842 4868
rect 15858 4924 15922 4928
rect 15858 4868 15862 4924
rect 15862 4868 15918 4924
rect 15918 4868 15922 4924
rect 15858 4864 15922 4868
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 4698 4380 4762 4384
rect 4698 4324 4702 4380
rect 4702 4324 4758 4380
rect 4758 4324 4762 4380
rect 4698 4320 4762 4324
rect 4778 4380 4842 4384
rect 4778 4324 4782 4380
rect 4782 4324 4838 4380
rect 4838 4324 4842 4380
rect 4778 4320 4842 4324
rect 4858 4380 4922 4384
rect 4858 4324 4862 4380
rect 4862 4324 4918 4380
rect 4918 4324 4922 4380
rect 4858 4320 4922 4324
rect 11952 4380 12016 4384
rect 11952 4324 11956 4380
rect 11956 4324 12012 4380
rect 12012 4324 12016 4380
rect 11952 4320 12016 4324
rect 12032 4380 12096 4384
rect 12032 4324 12036 4380
rect 12036 4324 12092 4380
rect 12092 4324 12096 4380
rect 12032 4320 12096 4324
rect 12112 4380 12176 4384
rect 12112 4324 12116 4380
rect 12116 4324 12172 4380
rect 12172 4324 12176 4380
rect 12112 4320 12176 4324
rect 12192 4380 12256 4384
rect 12192 4324 12196 4380
rect 12196 4324 12252 4380
rect 12252 4324 12256 4380
rect 12192 4320 12256 4324
rect 19285 4380 19349 4384
rect 19285 4324 19289 4380
rect 19289 4324 19345 4380
rect 19345 4324 19349 4380
rect 19285 4320 19349 4324
rect 19365 4380 19429 4384
rect 19365 4324 19369 4380
rect 19369 4324 19425 4380
rect 19425 4324 19429 4380
rect 19365 4320 19429 4324
rect 19445 4380 19509 4384
rect 19445 4324 19449 4380
rect 19449 4324 19505 4380
rect 19505 4324 19509 4380
rect 19445 4320 19509 4324
rect 19525 4380 19589 4384
rect 19525 4324 19529 4380
rect 19529 4324 19585 4380
rect 19585 4324 19589 4380
rect 19525 4320 19589 4324
rect 9260 3980 9324 4044
rect 8285 3836 8349 3840
rect 8285 3780 8289 3836
rect 8289 3780 8345 3836
rect 8345 3780 8349 3836
rect 8285 3776 8349 3780
rect 8365 3836 8429 3840
rect 8365 3780 8369 3836
rect 8369 3780 8425 3836
rect 8425 3780 8429 3836
rect 8365 3776 8429 3780
rect 8445 3836 8509 3840
rect 8445 3780 8449 3836
rect 8449 3780 8505 3836
rect 8505 3780 8509 3836
rect 8445 3776 8509 3780
rect 8525 3836 8589 3840
rect 8525 3780 8529 3836
rect 8529 3780 8585 3836
rect 8585 3780 8589 3836
rect 8525 3776 8589 3780
rect 15618 3836 15682 3840
rect 15618 3780 15622 3836
rect 15622 3780 15678 3836
rect 15678 3780 15682 3836
rect 15618 3776 15682 3780
rect 15698 3836 15762 3840
rect 15698 3780 15702 3836
rect 15702 3780 15758 3836
rect 15758 3780 15762 3836
rect 15698 3776 15762 3780
rect 15778 3836 15842 3840
rect 15778 3780 15782 3836
rect 15782 3780 15838 3836
rect 15838 3780 15842 3836
rect 15778 3776 15842 3780
rect 15858 3836 15922 3840
rect 15858 3780 15862 3836
rect 15862 3780 15918 3836
rect 15918 3780 15922 3836
rect 15858 3776 15922 3780
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 4698 3292 4762 3296
rect 4698 3236 4702 3292
rect 4702 3236 4758 3292
rect 4758 3236 4762 3292
rect 4698 3232 4762 3236
rect 4778 3292 4842 3296
rect 4778 3236 4782 3292
rect 4782 3236 4838 3292
rect 4838 3236 4842 3292
rect 4778 3232 4842 3236
rect 4858 3292 4922 3296
rect 4858 3236 4862 3292
rect 4862 3236 4918 3292
rect 4918 3236 4922 3292
rect 4858 3232 4922 3236
rect 11952 3292 12016 3296
rect 11952 3236 11956 3292
rect 11956 3236 12012 3292
rect 12012 3236 12016 3292
rect 11952 3232 12016 3236
rect 12032 3292 12096 3296
rect 12032 3236 12036 3292
rect 12036 3236 12092 3292
rect 12092 3236 12096 3292
rect 12032 3232 12096 3236
rect 12112 3292 12176 3296
rect 12112 3236 12116 3292
rect 12116 3236 12172 3292
rect 12172 3236 12176 3292
rect 12112 3232 12176 3236
rect 12192 3292 12256 3296
rect 12192 3236 12196 3292
rect 12196 3236 12252 3292
rect 12252 3236 12256 3292
rect 12192 3232 12256 3236
rect 19285 3292 19349 3296
rect 19285 3236 19289 3292
rect 19289 3236 19345 3292
rect 19345 3236 19349 3292
rect 19285 3232 19349 3236
rect 19365 3292 19429 3296
rect 19365 3236 19369 3292
rect 19369 3236 19425 3292
rect 19425 3236 19429 3292
rect 19365 3232 19429 3236
rect 19445 3292 19509 3296
rect 19445 3236 19449 3292
rect 19449 3236 19505 3292
rect 19505 3236 19509 3292
rect 19445 3232 19509 3236
rect 19525 3292 19589 3296
rect 19525 3236 19529 3292
rect 19529 3236 19585 3292
rect 19585 3236 19589 3292
rect 19525 3232 19589 3236
rect 8285 2748 8349 2752
rect 8285 2692 8289 2748
rect 8289 2692 8345 2748
rect 8345 2692 8349 2748
rect 8285 2688 8349 2692
rect 8365 2748 8429 2752
rect 8365 2692 8369 2748
rect 8369 2692 8425 2748
rect 8425 2692 8429 2748
rect 8365 2688 8429 2692
rect 8445 2748 8509 2752
rect 8445 2692 8449 2748
rect 8449 2692 8505 2748
rect 8505 2692 8509 2748
rect 8445 2688 8509 2692
rect 8525 2748 8589 2752
rect 8525 2692 8529 2748
rect 8529 2692 8585 2748
rect 8585 2692 8589 2748
rect 8525 2688 8589 2692
rect 15618 2748 15682 2752
rect 15618 2692 15622 2748
rect 15622 2692 15678 2748
rect 15678 2692 15682 2748
rect 15618 2688 15682 2692
rect 15698 2748 15762 2752
rect 15698 2692 15702 2748
rect 15702 2692 15758 2748
rect 15758 2692 15762 2748
rect 15698 2688 15762 2692
rect 15778 2748 15842 2752
rect 15778 2692 15782 2748
rect 15782 2692 15838 2748
rect 15838 2692 15842 2748
rect 15778 2688 15842 2692
rect 15858 2748 15922 2752
rect 15858 2692 15862 2748
rect 15862 2692 15918 2748
rect 15918 2692 15922 2748
rect 15858 2688 15922 2692
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 4698 2204 4762 2208
rect 4698 2148 4702 2204
rect 4702 2148 4758 2204
rect 4758 2148 4762 2204
rect 4698 2144 4762 2148
rect 4778 2204 4842 2208
rect 4778 2148 4782 2204
rect 4782 2148 4838 2204
rect 4838 2148 4842 2204
rect 4778 2144 4842 2148
rect 4858 2204 4922 2208
rect 4858 2148 4862 2204
rect 4862 2148 4918 2204
rect 4918 2148 4922 2204
rect 4858 2144 4922 2148
rect 11952 2204 12016 2208
rect 11952 2148 11956 2204
rect 11956 2148 12012 2204
rect 12012 2148 12016 2204
rect 11952 2144 12016 2148
rect 12032 2204 12096 2208
rect 12032 2148 12036 2204
rect 12036 2148 12092 2204
rect 12092 2148 12096 2204
rect 12032 2144 12096 2148
rect 12112 2204 12176 2208
rect 12112 2148 12116 2204
rect 12116 2148 12172 2204
rect 12172 2148 12176 2204
rect 12112 2144 12176 2148
rect 12192 2204 12256 2208
rect 12192 2148 12196 2204
rect 12196 2148 12252 2204
rect 12252 2148 12256 2204
rect 12192 2144 12256 2148
rect 19285 2204 19349 2208
rect 19285 2148 19289 2204
rect 19289 2148 19345 2204
rect 19345 2148 19349 2204
rect 19285 2144 19349 2148
rect 19365 2204 19429 2208
rect 19365 2148 19369 2204
rect 19369 2148 19425 2204
rect 19425 2148 19429 2204
rect 19365 2144 19429 2148
rect 19445 2204 19509 2208
rect 19445 2148 19449 2204
rect 19449 2148 19505 2204
rect 19505 2148 19509 2204
rect 19445 2144 19509 2148
rect 19525 2204 19589 2208
rect 19525 2148 19529 2204
rect 19529 2148 19585 2204
rect 19585 2148 19589 2204
rect 19525 2144 19589 2148
<< metal4 >>
rect 4610 19616 4931 19632
rect 4610 19552 4618 19616
rect 4682 19552 4698 19616
rect 4762 19552 4778 19616
rect 4842 19552 4858 19616
rect 4922 19552 4931 19616
rect 4610 18528 4931 19552
rect 4610 18464 4618 18528
rect 4682 18464 4698 18528
rect 4762 18464 4778 18528
rect 4842 18464 4858 18528
rect 4922 18464 4931 18528
rect 4610 17440 4931 18464
rect 4610 17376 4618 17440
rect 4682 17376 4698 17440
rect 4762 17376 4778 17440
rect 4842 17376 4858 17440
rect 4922 17376 4931 17440
rect 4610 16352 4931 17376
rect 4610 16288 4618 16352
rect 4682 16288 4698 16352
rect 4762 16288 4778 16352
rect 4842 16288 4858 16352
rect 4922 16288 4931 16352
rect 4610 15264 4931 16288
rect 4610 15200 4618 15264
rect 4682 15200 4698 15264
rect 4762 15200 4778 15264
rect 4842 15200 4858 15264
rect 4922 15200 4931 15264
rect 4610 14176 4931 15200
rect 4610 14112 4618 14176
rect 4682 14112 4698 14176
rect 4762 14112 4778 14176
rect 4842 14112 4858 14176
rect 4922 14112 4931 14176
rect 4610 13088 4931 14112
rect 8277 19072 8597 19632
rect 8277 19008 8285 19072
rect 8349 19008 8365 19072
rect 8429 19008 8445 19072
rect 8509 19008 8525 19072
rect 8589 19008 8597 19072
rect 8277 17984 8597 19008
rect 8277 17920 8285 17984
rect 8349 17920 8365 17984
rect 8429 17920 8445 17984
rect 8509 17920 8525 17984
rect 8589 17920 8597 17984
rect 8277 16896 8597 17920
rect 8277 16832 8285 16896
rect 8349 16832 8365 16896
rect 8429 16832 8445 16896
rect 8509 16832 8525 16896
rect 8589 16832 8597 16896
rect 8277 15808 8597 16832
rect 8277 15744 8285 15808
rect 8349 15744 8365 15808
rect 8429 15744 8445 15808
rect 8509 15744 8525 15808
rect 8589 15744 8597 15808
rect 8277 14720 8597 15744
rect 8277 14656 8285 14720
rect 8349 14656 8365 14720
rect 8429 14656 8445 14720
rect 8509 14656 8525 14720
rect 8589 14656 8597 14720
rect 7971 13836 8037 13837
rect 7971 13772 7972 13836
rect 8036 13772 8037 13836
rect 7971 13771 8037 13772
rect 4610 13024 4618 13088
rect 4682 13024 4698 13088
rect 4762 13024 4778 13088
rect 4842 13024 4858 13088
rect 4922 13024 4931 13088
rect 4610 12000 4931 13024
rect 4610 11936 4618 12000
rect 4682 11936 4698 12000
rect 4762 11936 4778 12000
rect 4842 11936 4858 12000
rect 4922 11936 4931 12000
rect 4610 10912 4931 11936
rect 4610 10848 4618 10912
rect 4682 10848 4698 10912
rect 4762 10848 4778 10912
rect 4842 10848 4858 10912
rect 4922 10848 4931 10912
rect 4610 9824 4931 10848
rect 4610 9760 4618 9824
rect 4682 9760 4698 9824
rect 4762 9760 4778 9824
rect 4842 9760 4858 9824
rect 4922 9760 4931 9824
rect 4610 8736 4931 9760
rect 4610 8672 4618 8736
rect 4682 8672 4698 8736
rect 4762 8672 4778 8736
rect 4842 8672 4858 8736
rect 4922 8672 4931 8736
rect 59 7988 125 7989
rect 59 7924 60 7988
rect 124 7924 125 7988
rect 59 7923 125 7924
rect 62 7717 122 7923
rect 59 7716 125 7717
rect 59 7652 60 7716
rect 124 7652 125 7716
rect 59 7651 125 7652
rect 4610 7648 4931 8672
rect 7974 8533 8034 13771
rect 8277 13632 8597 14656
rect 8277 13568 8285 13632
rect 8349 13568 8365 13632
rect 8429 13568 8445 13632
rect 8509 13568 8525 13632
rect 8589 13568 8597 13632
rect 8277 12544 8597 13568
rect 8277 12480 8285 12544
rect 8349 12480 8365 12544
rect 8429 12480 8445 12544
rect 8509 12480 8525 12544
rect 8589 12480 8597 12544
rect 8277 11456 8597 12480
rect 8277 11392 8285 11456
rect 8349 11392 8365 11456
rect 8429 11392 8445 11456
rect 8509 11392 8525 11456
rect 8589 11392 8597 11456
rect 8277 10368 8597 11392
rect 8277 10304 8285 10368
rect 8349 10304 8365 10368
rect 8429 10304 8445 10368
rect 8509 10304 8525 10368
rect 8589 10304 8597 10368
rect 8277 9280 8597 10304
rect 8277 9216 8285 9280
rect 8349 9216 8365 9280
rect 8429 9216 8445 9280
rect 8509 9216 8525 9280
rect 8589 9216 8597 9280
rect 7971 8532 8037 8533
rect 7971 8468 7972 8532
rect 8036 8468 8037 8532
rect 7971 8467 8037 8468
rect 4610 7584 4618 7648
rect 4682 7584 4698 7648
rect 4762 7584 4778 7648
rect 4842 7584 4858 7648
rect 4922 7584 4931 7648
rect 4610 6560 4931 7584
rect 4610 6496 4618 6560
rect 4682 6496 4698 6560
rect 4762 6496 4778 6560
rect 4842 6496 4858 6560
rect 4922 6496 4931 6560
rect 4610 5472 4931 6496
rect 4610 5408 4618 5472
rect 4682 5408 4698 5472
rect 4762 5408 4778 5472
rect 4842 5408 4858 5472
rect 4922 5408 4931 5472
rect 4610 4384 4931 5408
rect 4610 4320 4618 4384
rect 4682 4320 4698 4384
rect 4762 4320 4778 4384
rect 4842 4320 4858 4384
rect 4922 4320 4931 4384
rect 4610 3296 4931 4320
rect 4610 3232 4618 3296
rect 4682 3232 4698 3296
rect 4762 3232 4778 3296
rect 4842 3232 4858 3296
rect 4922 3232 4931 3296
rect 4610 2208 4931 3232
rect 4610 2144 4618 2208
rect 4682 2144 4698 2208
rect 4762 2144 4778 2208
rect 4842 2144 4858 2208
rect 4922 2144 4931 2208
rect 4610 2128 4931 2144
rect 8277 8192 8597 9216
rect 11944 19616 12264 19632
rect 11944 19552 11952 19616
rect 12016 19552 12032 19616
rect 12096 19552 12112 19616
rect 12176 19552 12192 19616
rect 12256 19552 12264 19616
rect 11944 18528 12264 19552
rect 11944 18464 11952 18528
rect 12016 18464 12032 18528
rect 12096 18464 12112 18528
rect 12176 18464 12192 18528
rect 12256 18464 12264 18528
rect 11944 17440 12264 18464
rect 11944 17376 11952 17440
rect 12016 17376 12032 17440
rect 12096 17376 12112 17440
rect 12176 17376 12192 17440
rect 12256 17376 12264 17440
rect 11944 16352 12264 17376
rect 11944 16288 11952 16352
rect 12016 16288 12032 16352
rect 12096 16288 12112 16352
rect 12176 16288 12192 16352
rect 12256 16288 12264 16352
rect 11944 15264 12264 16288
rect 11944 15200 11952 15264
rect 12016 15200 12032 15264
rect 12096 15200 12112 15264
rect 12176 15200 12192 15264
rect 12256 15200 12264 15264
rect 11944 14176 12264 15200
rect 11944 14112 11952 14176
rect 12016 14112 12032 14176
rect 12096 14112 12112 14176
rect 12176 14112 12192 14176
rect 12256 14112 12264 14176
rect 11944 13088 12264 14112
rect 11944 13024 11952 13088
rect 12016 13024 12032 13088
rect 12096 13024 12112 13088
rect 12176 13024 12192 13088
rect 12256 13024 12264 13088
rect 11944 12000 12264 13024
rect 11944 11936 11952 12000
rect 12016 11936 12032 12000
rect 12096 11936 12112 12000
rect 12176 11936 12192 12000
rect 12256 11936 12264 12000
rect 11944 10912 12264 11936
rect 11944 10848 11952 10912
rect 12016 10848 12032 10912
rect 12096 10848 12112 10912
rect 12176 10848 12192 10912
rect 12256 10848 12264 10912
rect 11944 9824 12264 10848
rect 11944 9760 11952 9824
rect 12016 9760 12032 9824
rect 12096 9760 12112 9824
rect 12176 9760 12192 9824
rect 12256 9760 12264 9824
rect 11944 8736 12264 9760
rect 11944 8672 11952 8736
rect 12016 8672 12032 8736
rect 12096 8672 12112 8736
rect 12176 8672 12192 8736
rect 12256 8672 12264 8736
rect 9259 8532 9325 8533
rect 9259 8468 9260 8532
rect 9324 8468 9325 8532
rect 9259 8467 9325 8468
rect 8277 8128 8285 8192
rect 8349 8128 8365 8192
rect 8429 8128 8445 8192
rect 8509 8128 8525 8192
rect 8589 8128 8597 8192
rect 8277 7104 8597 8128
rect 8277 7040 8285 7104
rect 8349 7040 8365 7104
rect 8429 7040 8445 7104
rect 8509 7040 8525 7104
rect 8589 7040 8597 7104
rect 8277 6016 8597 7040
rect 8277 5952 8285 6016
rect 8349 5952 8365 6016
rect 8429 5952 8445 6016
rect 8509 5952 8525 6016
rect 8589 5952 8597 6016
rect 8277 4928 8597 5952
rect 8277 4864 8285 4928
rect 8349 4864 8365 4928
rect 8429 4864 8445 4928
rect 8509 4864 8525 4928
rect 8589 4864 8597 4928
rect 8277 3840 8597 4864
rect 9262 4045 9322 8467
rect 11944 7648 12264 8672
rect 11944 7584 11952 7648
rect 12016 7584 12032 7648
rect 12096 7584 12112 7648
rect 12176 7584 12192 7648
rect 12256 7584 12264 7648
rect 11944 6560 12264 7584
rect 11944 6496 11952 6560
rect 12016 6496 12032 6560
rect 12096 6496 12112 6560
rect 12176 6496 12192 6560
rect 12256 6496 12264 6560
rect 11944 5472 12264 6496
rect 11944 5408 11952 5472
rect 12016 5408 12032 5472
rect 12096 5408 12112 5472
rect 12176 5408 12192 5472
rect 12256 5408 12264 5472
rect 11944 4384 12264 5408
rect 11944 4320 11952 4384
rect 12016 4320 12032 4384
rect 12096 4320 12112 4384
rect 12176 4320 12192 4384
rect 12256 4320 12264 4384
rect 9259 4044 9325 4045
rect 9259 3980 9260 4044
rect 9324 3980 9325 4044
rect 9259 3979 9325 3980
rect 8277 3776 8285 3840
rect 8349 3776 8365 3840
rect 8429 3776 8445 3840
rect 8509 3776 8525 3840
rect 8589 3776 8597 3840
rect 8277 2752 8597 3776
rect 8277 2688 8285 2752
rect 8349 2688 8365 2752
rect 8429 2688 8445 2752
rect 8509 2688 8525 2752
rect 8589 2688 8597 2752
rect 8277 2128 8597 2688
rect 11944 3296 12264 4320
rect 11944 3232 11952 3296
rect 12016 3232 12032 3296
rect 12096 3232 12112 3296
rect 12176 3232 12192 3296
rect 12256 3232 12264 3296
rect 11944 2208 12264 3232
rect 11944 2144 11952 2208
rect 12016 2144 12032 2208
rect 12096 2144 12112 2208
rect 12176 2144 12192 2208
rect 12256 2144 12264 2208
rect 11944 2128 12264 2144
rect 15610 19072 15930 19632
rect 15610 19008 15618 19072
rect 15682 19008 15698 19072
rect 15762 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15930 19072
rect 15610 17984 15930 19008
rect 15610 17920 15618 17984
rect 15682 17920 15698 17984
rect 15762 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15930 17984
rect 15610 16896 15930 17920
rect 15610 16832 15618 16896
rect 15682 16832 15698 16896
rect 15762 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15930 16896
rect 15610 15808 15930 16832
rect 15610 15744 15618 15808
rect 15682 15744 15698 15808
rect 15762 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15930 15808
rect 15610 14720 15930 15744
rect 15610 14656 15618 14720
rect 15682 14656 15698 14720
rect 15762 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15930 14720
rect 15610 13632 15930 14656
rect 15610 13568 15618 13632
rect 15682 13568 15698 13632
rect 15762 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15930 13632
rect 15610 12544 15930 13568
rect 15610 12480 15618 12544
rect 15682 12480 15698 12544
rect 15762 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15930 12544
rect 15610 11456 15930 12480
rect 15610 11392 15618 11456
rect 15682 11392 15698 11456
rect 15762 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15930 11456
rect 15610 10368 15930 11392
rect 15610 10304 15618 10368
rect 15682 10304 15698 10368
rect 15762 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15930 10368
rect 15610 9280 15930 10304
rect 15610 9216 15618 9280
rect 15682 9216 15698 9280
rect 15762 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15930 9280
rect 15610 8192 15930 9216
rect 15610 8128 15618 8192
rect 15682 8128 15698 8192
rect 15762 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15930 8192
rect 15610 7104 15930 8128
rect 15610 7040 15618 7104
rect 15682 7040 15698 7104
rect 15762 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15930 7104
rect 15610 6016 15930 7040
rect 15610 5952 15618 6016
rect 15682 5952 15698 6016
rect 15762 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15930 6016
rect 15610 4928 15930 5952
rect 15610 4864 15618 4928
rect 15682 4864 15698 4928
rect 15762 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15930 4928
rect 15610 3840 15930 4864
rect 15610 3776 15618 3840
rect 15682 3776 15698 3840
rect 15762 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15930 3840
rect 15610 2752 15930 3776
rect 15610 2688 15618 2752
rect 15682 2688 15698 2752
rect 15762 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15930 2752
rect 15610 2128 15930 2688
rect 19277 19616 19597 19632
rect 19277 19552 19285 19616
rect 19349 19552 19365 19616
rect 19429 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19597 19616
rect 19277 18528 19597 19552
rect 19277 18464 19285 18528
rect 19349 18464 19365 18528
rect 19429 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19597 18528
rect 19277 17440 19597 18464
rect 19277 17376 19285 17440
rect 19349 17376 19365 17440
rect 19429 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19597 17440
rect 19277 16352 19597 17376
rect 19277 16288 19285 16352
rect 19349 16288 19365 16352
rect 19429 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19597 16352
rect 19277 15264 19597 16288
rect 19277 15200 19285 15264
rect 19349 15200 19365 15264
rect 19429 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19597 15264
rect 19277 14176 19597 15200
rect 19277 14112 19285 14176
rect 19349 14112 19365 14176
rect 19429 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19597 14176
rect 19277 13088 19597 14112
rect 21587 13700 21653 13701
rect 21587 13636 21588 13700
rect 21652 13636 21653 13700
rect 21587 13635 21653 13636
rect 21590 13429 21650 13635
rect 21587 13428 21653 13429
rect 21587 13364 21588 13428
rect 21652 13364 21653 13428
rect 21587 13363 21653 13364
rect 19277 13024 19285 13088
rect 19349 13024 19365 13088
rect 19429 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19597 13088
rect 19277 12000 19597 13024
rect 19277 11936 19285 12000
rect 19349 11936 19365 12000
rect 19429 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19597 12000
rect 19277 10912 19597 11936
rect 19277 10848 19285 10912
rect 19349 10848 19365 10912
rect 19429 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19597 10912
rect 19277 9824 19597 10848
rect 19277 9760 19285 9824
rect 19349 9760 19365 9824
rect 19429 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19597 9824
rect 19277 8736 19597 9760
rect 19277 8672 19285 8736
rect 19349 8672 19365 8736
rect 19429 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19597 8736
rect 19277 7648 19597 8672
rect 19277 7584 19285 7648
rect 19349 7584 19365 7648
rect 19429 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19597 7648
rect 19277 6560 19597 7584
rect 19277 6496 19285 6560
rect 19349 6496 19365 6560
rect 19429 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19597 6560
rect 19277 5472 19597 6496
rect 19277 5408 19285 5472
rect 19349 5408 19365 5472
rect 19429 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19597 5472
rect 19277 4384 19597 5408
rect 19277 4320 19285 4384
rect 19349 4320 19365 4384
rect 19429 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19597 4384
rect 19277 3296 19597 4320
rect 19277 3232 19285 3296
rect 19349 3232 19365 3296
rect 19429 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19597 3296
rect 19277 2208 19597 3232
rect 19277 2144 19285 2208
rect 19349 2144 19365 2208
rect 19429 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19597 2208
rect 19277 2128 19597 2144
use scs8hd_decap_3  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 314 592
use scs8hd_conb_1  _70_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_13 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_9
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_11
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_28
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_32
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_64 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_35
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__D
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use scs8hd_nor4_4  _63_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_39
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__62__B
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__D
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__B
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_or2_4  _37_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 682 592
use scs8hd_fill_2  FILLER_1_69
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__D
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_nor4_4  _64_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1602 592
use scs8hd_nor4_4  _44_
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__44__C
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__B
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_80
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_73
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__77__A
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_99
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_105
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__C
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_0_109
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__D
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__B
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__C
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__B
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_nor4_4  _39_
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13524 0 -1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__C
timestamp 1586364061
transform 1 0 12788 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_129 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_150
timestamp 1586364061
transform 1 0 14904 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__D
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_159
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_154 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15088 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_1_168
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_163
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_172
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_176
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_204
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_204
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 20884 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 20884 0 -1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 1050 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__63__C
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__C
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_20
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_24
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_nor4_4  _62_
timestamp 1586364061
transform 1 0 4968 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__63__B
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__62__D
timestamp 1586364061
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_38
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _65_
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__65__B
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 6716 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_59
timestamp 1586364061
transform 1 0 6532 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_63
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__B
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _40_
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 1602 592
use scs8hd_buf_2  _77_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__B
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_98
timestamp 1586364061
transform 1 0 10120 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_123
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__B
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_128
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_140
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__47__D
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__D
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_148
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_152
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_203 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__62__C
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__60__C
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_32
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _29_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__29__A
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__60__D
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_49
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__B
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__60__B
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_68
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _43_
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_3_89
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_93
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _72_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__72__A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__C
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_108
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _47_
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__47__C
timestamp 1586364061
transform 1 0 13708 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_127
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_131
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_177
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 20884 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__30__A
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__C
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__D
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_22
timestamp 1586364061
transform 1 0 3128 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__B
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_47
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_51
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _60_
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 1602 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__C
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__D
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_72
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_76
timestamp 1586364061
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_or2_4  _52_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__D
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_100
timestamp 1586364061
transform 1 0 10304 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11132 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_108
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_120
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_124
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _46_
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__46__B
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15548 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__48__C
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__D
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17296 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_172
timestamp 1586364061
transform 1 0 16928 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _35_
timestamp 1586364061
transform 1 0 18860 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_185
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_189
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _30_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_12
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_17
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _33_
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__38__C
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__61__C
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_30
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_or4_4  _53_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__61__D
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__B
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6992 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__61__B
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_55
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _42_
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__42__C
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__B
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_79
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__78__A
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__D
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_100
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_104
timestamp 1586364061
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_buf_2  _78_
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__41__B
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_116
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use scs8hd_nor4_4  _48_
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__48__B
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__89__A
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_133
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_158
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _71_
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 20884 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_8
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _85_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__85__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 314 592
use scs8hd_inv_8  _34_
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_22
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_18
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_24
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_20
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__28__A
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__D
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_or4_4  _38_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_8  _28_
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__54__B
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__25__A
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_46
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 314 592
use scs8hd_nor4_4  _61_
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 1602 592
use scs8hd_inv_8  _25_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_or4_4  _45_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__C
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_66
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_70
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_79
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_74
timestamp 1586364061
transform 1 0 7912 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__55__B
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__55__C
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_89
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__56__C
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_93
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__56__B
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__B
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__C
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 866 592
use scs8hd_nor4_4  _59_
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 1602 592
use scs8hd_nor4_4  _41_
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 1602 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__57__C
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__C
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__D
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_120
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_130
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_126
timestamp 1586364061
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_131
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__B
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_137
timestamp 1586364061
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 13524 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 13892 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__C
timestamp 1586364061
transform 1 0 13708 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _89_
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 406 592
use scs8hd_nor4_4  _51_
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__D
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__D
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_160
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__C
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17388 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__49__B
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_169
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_173
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__84__A
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _36_
timestamp 1586364061
transform 1 0 18952 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 20884 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 20884 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_203
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_198
timestamp 1586364061
transform 1 0 19320 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_13
timestamp 1586364061
transform 1 0 2300 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_17
timestamp 1586364061
transform 1 0 2668 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_21
timestamp 1586364061
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_25
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_29
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use scs8hd_nor4_4  _54_
timestamp 1586364061
transform 1 0 4968 0 -1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__45__B
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_38
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _55_
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__45__C
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_59
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__45__D
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _56_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _57_
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__D
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_110
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_114
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__B
timestamp 1586364061
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_135
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _49_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__50__C
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17020 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_171
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_175
timestamp 1586364061
transform 1 0 17204 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _84_
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_188
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_192
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 20884 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_200 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _26_
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__26__A
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__54__D
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_36
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_40
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _58_
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__C
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_66
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__56__D
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_90
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_105
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__D
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_109
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_116
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_120
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _50_
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__B
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_126
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_155
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use scs8hd_buf_2  _81_
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 406 592
use scs8hd_buf_2  _87_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__87__A
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_188
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_192
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 20884 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__81__A
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_200
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_204
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4324 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use scs8hd_conb_1  _69_
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_40
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__B
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_59
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__58__D
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_104
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_108
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_142
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__50__D
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_146 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14536 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_169
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_182
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 774 592
use scs8hd_conb_1  _68_
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_204
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_11_31
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 590 592
use scs8hd_inv_8  _27_
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__27__A
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_52
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_56
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__55__D
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_77
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_84
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_116
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_120
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_149
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_153
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_157
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_162
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__86__A
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 20884 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_204
timestamp 1586364061
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1472 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_19
timestamp 1586364061
transform 1 0 2852 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_inv_8  _32_
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_78
timestamp 1586364061
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_82
timestamp 1586364061
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_86
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_90
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_100
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_104
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_108
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_120
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_137
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_142
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_146
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_158
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_175
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_2  _86_
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17940 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_42
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_46
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_67
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_72
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_89
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _80_
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_96
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_100
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_104
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_8  _24_
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__24__A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__80__A
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_111
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_115
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_119
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_114
timestamp 1586364061
transform 1 0 11592 0 -1 10336
box -38 -48 590 592
use scs8hd_conb_1  _66_
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_145
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_160
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _83_
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__83__A
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_164
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_172
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_176
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_187
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_191
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 20884 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_198
timestamp 1586364061
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_202
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use scs8hd_inv_8  _31_
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__31__A
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_88
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_95
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_99
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_103
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_126
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_130
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_154
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_166
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__76__A
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_182
timestamp 1586364061
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_15_192
timestamp 1586364061
transform 1 0 18768 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 20884 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_15_209
timestamp 1586364061
transform 1 0 20332 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 1142 592
use scs8hd_conb_1  _67_
timestamp 1586364061
transform 1 0 8188 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_76
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_108
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_132
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _76_
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_4  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_194
timestamp 1586364061
transform 1 0 18952 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 20884 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _74_
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__74__A
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_192
timestamp 1586364061
transform 1 0 18768 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_194
timestamp 1586364061
transform 1 0 18952 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 20884 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_19_209
timestamp 1586364061
transform 1 0 20332 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 20884 0 1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_210
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__88__A
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_19
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_31
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_43
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_23_55
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 590 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 20884 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 406 592
use scs8hd_buf_2  _88_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 20884 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 20884 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 20884 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_2  _82_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__82__A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 130 592
use scs8hd_buf_2  _79_
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__79__A
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_40
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_44
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _75_
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_56
timestamp 1586364061
transform 1 0 6256 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_60
timestamp 1586364061
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_68
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__75__A
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_73
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_77
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_89
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_29_113
timestamp 1586364061
transform 1 0 11500 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 20884 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_210
timestamp 1586364061
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_31_32
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_63
timestamp 1586364061
transform 1 0 6900 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_31_87
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_106
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12512 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_125
timestamp 1586364061
transform 1 0 12604 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_137
timestamp 1586364061
transform 1 0 13708 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_149
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_168
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 18216 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_180
timestamp 1586364061
transform 1 0 17664 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_187
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 20884 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_199
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_31_211
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 130 592
<< labels >>
rlabel metal3 s 21520 824 22000 944 6 address[0]
port 0 nsew default input
rlabel metal2 s 2502 0 2558 480 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 1096 480 1216 6 address[2]
port 2 nsew default input
rlabel metal2 s 3606 0 3662 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 4618 0 4674 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 5630 0 5686 480 6 address[5]
port 5 nsew default input
rlabel metal3 s 0 3272 480 3392 6 bottom_grid_pin_0_
port 6 nsew default tristate
rlabel metal2 s 6734 0 6790 480 6 bottom_grid_pin_4_
port 7 nsew default tristate
rlabel metal3 s 21520 2592 22000 2712 6 bottom_grid_pin_8_
port 8 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal3 s 21520 4496 22000 4616 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal2 s 8850 0 8906 480 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 21520 6264 22000 6384 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal3 s 0 5448 480 5568 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal2 s 9862 0 9918 480 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 21520 8168 22000 8288 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal2 s 1582 21520 1638 22000 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal3 s 21520 9936 22000 10056 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal2 s 4710 21520 4766 22000 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal2 s 10874 0 10930 480 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal2 s 11978 0 12034 480 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal3 s 21520 11840 22000 11960 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal2 s 7838 21520 7894 22000 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal3 s 21520 13608 22000 13728 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal2 s 12990 0 13046 480 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal2 s 14002 0 14058 480 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal2 s 10966 21520 11022 22000 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal3 s 21520 15512 22000 15632 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal3 s 21520 17280 22000 17400 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal3 s 0 12112 480 12232 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal2 s 15106 0 15162 480 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 21520 19184 22000 19304 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal2 s 14094 21520 14150 22000 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal2 s 16118 0 16174 480 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal2 s 17222 0 17278 480 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 21520 20952 22000 21072 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal2 s 17222 21520 17278 22000 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal2 s 19246 0 19302 480 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 1490 0 1546 480 6 data_in
port 45 nsew default input
rlabel metal2 s 478 0 534 480 6 enable
port 46 nsew default input
rlabel metal2 s 21362 0 21418 480 6 top_grid_pin_14_
port 47 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 top_grid_pin_2_
port 48 nsew default tristate
rlabel metal2 s 20350 21520 20406 22000 6 top_grid_pin_6_
port 49 nsew default tristate
rlabel metal4 s 4611 2128 4931 19632 6 vpwr
port 50 nsew default input
rlabel metal4 s 8277 2128 8597 19632 6 vgnd
port 51 nsew default input
<< end >>
