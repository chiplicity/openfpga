magic
tech EFS8A
magscale 1 2
timestamp 1603801028
<< locali >>
rect 15669 22423 15703 22525
rect 11621 20315 11655 20417
rect 12081 5015 12115 5253
<< viali >>
rect 9965 25381 9999 25415
rect 12700 25313 12734 25347
rect 9873 25245 9907 25279
rect 10149 25245 10183 25279
rect 10793 25109 10827 25143
rect 12771 25109 12805 25143
rect 12725 24905 12759 24939
rect 5733 24769 5767 24803
rect 8585 24769 8619 24803
rect 9781 24769 9815 24803
rect 15945 24769 15979 24803
rect 5340 24701 5374 24735
rect 8100 24701 8134 24735
rect 13277 24701 13311 24735
rect 13829 24701 13863 24735
rect 15460 24701 15494 24735
rect 9137 24633 9171 24667
rect 9229 24633 9263 24667
rect 10701 24633 10735 24667
rect 10793 24633 10827 24667
rect 11345 24633 11379 24667
rect 5411 24565 5445 24599
rect 6837 24565 6871 24599
rect 8171 24565 8205 24599
rect 8953 24565 8987 24599
rect 10057 24565 10091 24599
rect 10517 24565 10551 24599
rect 13461 24565 13495 24599
rect 15531 24565 15565 24599
rect 4491 24361 4525 24395
rect 9137 24361 9171 24395
rect 18245 24361 18279 24395
rect 6561 24293 6595 24327
rect 8125 24293 8159 24327
rect 8217 24293 8251 24327
rect 10885 24293 10919 24327
rect 11437 24293 11471 24327
rect 13001 24293 13035 24327
rect 1476 24225 1510 24259
rect 4420 24225 4454 24259
rect 5432 24225 5466 24259
rect 8769 24225 8803 24259
rect 15368 24225 15402 24259
rect 16313 24225 16347 24259
rect 18061 24225 18095 24259
rect 6469 24157 6503 24191
rect 6745 24157 6779 24191
rect 9689 24157 9723 24191
rect 10793 24157 10827 24191
rect 12909 24157 12943 24191
rect 13553 24157 13587 24191
rect 1547 24089 1581 24123
rect 10149 24089 10183 24123
rect 16497 24089 16531 24123
rect 5273 24021 5307 24055
rect 5503 24021 5537 24055
rect 7573 24021 7607 24055
rect 10609 24021 10643 24055
rect 14105 24021 14139 24055
rect 15439 24021 15473 24055
rect 2237 23817 2271 23851
rect 4997 23817 5031 23851
rect 6285 23817 6319 23851
rect 8861 23817 8895 23851
rect 9183 23817 9217 23851
rect 9965 23817 9999 23851
rect 11529 23817 11563 23851
rect 12173 23817 12207 23851
rect 15945 23817 15979 23851
rect 16681 23817 16715 23851
rect 17049 23817 17083 23851
rect 19257 23817 19291 23851
rect 21281 23817 21315 23851
rect 22385 23817 22419 23851
rect 6561 23749 6595 23783
rect 8493 23749 8527 23783
rect 1547 23681 1581 23715
rect 5273 23681 5307 23715
rect 7849 23681 7883 23715
rect 10609 23681 10643 23715
rect 12541 23681 12575 23715
rect 12817 23681 12851 23715
rect 14381 23681 14415 23715
rect 1444 23613 1478 23647
rect 1869 23613 1903 23647
rect 2488 23613 2522 23647
rect 2881 23613 2915 23647
rect 4204 23613 4238 23647
rect 4629 23613 4663 23647
rect 9080 23613 9114 23647
rect 9505 23613 9539 23647
rect 15393 23613 15427 23647
rect 15761 23613 15795 23647
rect 16865 23613 16899 23647
rect 17417 23613 17451 23647
rect 18096 23613 18130 23647
rect 18199 23613 18233 23647
rect 19073 23613 19107 23647
rect 19625 23613 19659 23647
rect 21097 23613 21131 23647
rect 22201 23613 22235 23647
rect 22753 23613 22787 23647
rect 5365 23545 5399 23579
rect 5917 23545 5951 23579
rect 7573 23545 7607 23579
rect 7665 23545 7699 23579
rect 10701 23545 10735 23579
rect 11253 23545 11287 23579
rect 12633 23545 12667 23579
rect 14105 23545 14139 23579
rect 14197 23545 14231 23579
rect 18889 23545 18923 23579
rect 2559 23477 2593 23511
rect 4307 23477 4341 23511
rect 7297 23477 7331 23511
rect 10425 23477 10459 23511
rect 13461 23477 13495 23511
rect 13921 23477 13955 23511
rect 16405 23477 16439 23511
rect 18521 23477 18555 23511
rect 21649 23477 21683 23511
rect 5273 23273 5307 23307
rect 6561 23273 6595 23307
rect 10287 23273 10321 23307
rect 12541 23273 12575 23307
rect 12817 23273 12851 23307
rect 16451 23273 16485 23307
rect 5641 23205 5675 23239
rect 5733 23205 5767 23239
rect 7297 23205 7331 23239
rect 7849 23205 7883 23239
rect 11345 23205 11379 23239
rect 13829 23205 13863 23239
rect 10216 23137 10250 23171
rect 15336 23137 15370 23171
rect 16348 23137 16382 23171
rect 17360 23137 17394 23171
rect 6285 23069 6319 23103
rect 7205 23069 7239 23103
rect 11253 23069 11287 23103
rect 11529 23069 11563 23103
rect 13737 23069 13771 23103
rect 14197 23069 14231 23103
rect 15439 22933 15473 22967
rect 17463 22933 17497 22967
rect 5917 22729 5951 22763
rect 7113 22729 7147 22763
rect 10609 22729 10643 22763
rect 11345 22729 11379 22763
rect 12587 22729 12621 22763
rect 13369 22729 13403 22763
rect 16543 22729 16577 22763
rect 17325 22729 17359 22763
rect 11621 22661 11655 22695
rect 7665 22593 7699 22627
rect 7941 22593 7975 22627
rect 13921 22593 13955 22627
rect 15301 22593 15335 22627
rect 9689 22525 9723 22559
rect 10977 22525 11011 22559
rect 12516 22525 12550 22559
rect 12909 22525 12943 22559
rect 15460 22525 15494 22559
rect 15669 22525 15703 22559
rect 16440 22525 16474 22559
rect 7757 22457 7791 22491
rect 9597 22457 9631 22491
rect 10010 22457 10044 22491
rect 14013 22457 14047 22491
rect 14565 22457 14599 22491
rect 16221 22457 16255 22491
rect 16865 22457 16899 22491
rect 5641 22389 5675 22423
rect 6653 22389 6687 22423
rect 9137 22389 9171 22423
rect 13737 22389 13771 22423
rect 15531 22389 15565 22423
rect 15669 22389 15703 22423
rect 15945 22389 15979 22423
rect 5089 22185 5123 22219
rect 7573 22185 7607 22219
rect 11253 22185 11287 22219
rect 13921 22185 13955 22219
rect 14197 22185 14231 22219
rect 15393 22185 15427 22219
rect 6698 22117 6732 22151
rect 7941 22117 7975 22151
rect 10654 22117 10688 22151
rect 12862 22117 12896 22151
rect 5089 22049 5123 22083
rect 5365 22049 5399 22083
rect 8160 22049 8194 22083
rect 8585 22049 8619 22083
rect 13461 22049 13495 22083
rect 15577 22049 15611 22083
rect 15761 22049 15795 22083
rect 16871 22049 16905 22083
rect 6377 21981 6411 22015
rect 8263 21981 8297 22015
rect 10333 21981 10367 22015
rect 12541 21981 12575 22015
rect 17049 21913 17083 21947
rect 5917 21845 5951 21879
rect 7297 21845 7331 21879
rect 14565 21845 14599 21879
rect 16313 21845 16347 21879
rect 6193 21641 6227 21675
rect 6561 21641 6595 21675
rect 11897 21641 11931 21675
rect 13737 21641 13771 21675
rect 8677 21505 8711 21539
rect 9321 21505 9355 21539
rect 12725 21505 12759 21539
rect 14749 21505 14783 21539
rect 16129 21505 16163 21539
rect 5457 21437 5491 21471
rect 5641 21437 5675 21471
rect 5917 21437 5951 21471
rect 6837 21437 6871 21471
rect 10793 21437 10827 21471
rect 11253 21437 11287 21471
rect 7199 21369 7233 21403
rect 8769 21369 8803 21403
rect 10057 21369 10091 21403
rect 11529 21369 11563 21403
rect 12817 21369 12851 21403
rect 13369 21369 13403 21403
rect 14289 21369 14323 21403
rect 14381 21369 14415 21403
rect 15853 21369 15887 21403
rect 15945 21369 15979 21403
rect 4537 21301 4571 21335
rect 4905 21301 4939 21335
rect 7757 21301 7791 21335
rect 8217 21301 8251 21335
rect 10333 21301 10367 21335
rect 12265 21301 12299 21335
rect 14013 21301 14047 21335
rect 15301 21301 15335 21335
rect 16957 21301 16991 21335
rect 7021 21097 7055 21131
rect 8677 21097 8711 21131
rect 12725 21097 12759 21131
rect 13737 21097 13771 21131
rect 15025 21097 15059 21131
rect 16313 21097 16347 21131
rect 6377 21029 6411 21063
rect 6653 21029 6687 21063
rect 7389 21029 7423 21063
rect 7941 21029 7975 21063
rect 11253 21029 11287 21063
rect 13138 21029 13172 21063
rect 15393 21029 15427 21063
rect 15485 21029 15519 21063
rect 16037 21029 16071 21063
rect 4905 20961 4939 20995
rect 5641 20961 5675 20995
rect 6193 20961 6227 20995
rect 9756 20961 9790 20995
rect 7297 20893 7331 20927
rect 10793 20893 10827 20927
rect 11161 20893 11195 20927
rect 11621 20893 11655 20927
rect 12817 20893 12851 20927
rect 10333 20825 10367 20859
rect 5273 20757 5307 20791
rect 9827 20757 9861 20791
rect 14473 20757 14507 20791
rect 6193 20553 6227 20587
rect 6653 20553 6687 20587
rect 7297 20553 7331 20587
rect 10057 20553 10091 20587
rect 11069 20553 11103 20587
rect 13829 20553 13863 20587
rect 15761 20553 15795 20587
rect 8217 20485 8251 20519
rect 12173 20485 12207 20519
rect 15485 20485 15519 20519
rect 5917 20417 5951 20451
rect 9137 20417 9171 20451
rect 10793 20417 10827 20451
rect 11483 20417 11517 20451
rect 11621 20417 11655 20451
rect 14749 20417 14783 20451
rect 15945 20417 15979 20451
rect 5089 20349 5123 20383
rect 5365 20349 5399 20383
rect 5733 20349 5767 20383
rect 10425 20349 10459 20383
rect 11396 20349 11430 20383
rect 12633 20349 12667 20383
rect 13553 20349 13587 20383
rect 7665 20281 7699 20315
rect 7757 20281 7791 20315
rect 9458 20281 9492 20315
rect 11621 20281 11655 20315
rect 12954 20281 12988 20315
rect 14473 20281 14507 20315
rect 14565 20281 14599 20315
rect 8585 20213 8619 20247
rect 8953 20213 8987 20247
rect 11897 20213 11931 20247
rect 14197 20213 14231 20247
rect 5641 20009 5675 20043
rect 7113 20009 7147 20043
rect 7665 20009 7699 20043
rect 9137 20009 9171 20043
rect 11069 20009 11103 20043
rect 13277 20009 13311 20043
rect 6555 19941 6589 19975
rect 8125 19941 8159 19975
rect 10470 19941 10504 19975
rect 12081 19941 12115 19975
rect 12633 19941 12667 19975
rect 13829 19941 13863 19975
rect 5216 19873 5250 19907
rect 5319 19873 5353 19907
rect 15352 19873 15386 19907
rect 6193 19805 6227 19839
rect 8033 19805 8067 19839
rect 10149 19805 10183 19839
rect 11989 19805 12023 19839
rect 12909 19805 12943 19839
rect 13737 19805 13771 19839
rect 14381 19805 14415 19839
rect 8585 19737 8619 19771
rect 15439 19737 15473 19771
rect 6009 19669 6043 19703
rect 10057 19669 10091 19703
rect 11713 19669 11747 19703
rect 6285 19465 6319 19499
rect 6561 19465 6595 19499
rect 7757 19465 7791 19499
rect 8033 19465 8067 19499
rect 11897 19465 11931 19499
rect 13001 19465 13035 19499
rect 14105 19465 14139 19499
rect 14381 19397 14415 19431
rect 16037 19397 16071 19431
rect 5917 19329 5951 19363
rect 9597 19329 9631 19363
rect 4721 19261 4755 19295
rect 5457 19261 5491 19295
rect 5733 19261 5767 19295
rect 6837 19261 6871 19295
rect 8401 19261 8435 19295
rect 9045 19261 9079 19295
rect 9413 19261 9447 19295
rect 10701 19261 10735 19295
rect 11069 19261 11103 19295
rect 11529 19261 11563 19295
rect 12725 19261 12759 19295
rect 13185 19261 13219 19295
rect 14749 19261 14783 19295
rect 14933 19261 14967 19295
rect 15393 19261 15427 19295
rect 7158 19193 7192 19227
rect 11253 19193 11287 19227
rect 13506 19193 13540 19227
rect 5089 19125 5123 19159
rect 8861 19125 8895 19159
rect 10149 19125 10183 19159
rect 15209 19125 15243 19159
rect 10701 18921 10735 18955
rect 12449 18921 12483 18955
rect 13093 18921 13127 18955
rect 13921 18921 13955 18955
rect 14933 18921 14967 18955
rect 6653 18853 6687 18887
rect 7297 18853 7331 18887
rect 7665 18853 7699 18887
rect 10425 18853 10459 18887
rect 11437 18853 11471 18887
rect 5917 18785 5951 18819
rect 6469 18785 6503 18819
rect 9965 18785 9999 18819
rect 10241 18785 10275 18819
rect 13093 18785 13127 18819
rect 13369 18785 13403 18819
rect 15368 18785 15402 18819
rect 7573 18717 7607 18751
rect 8217 18717 8251 18751
rect 9045 18717 9079 18751
rect 11345 18717 11379 18751
rect 11621 18717 11655 18751
rect 5273 18581 5307 18615
rect 6929 18581 6963 18615
rect 14289 18581 14323 18615
rect 15439 18581 15473 18615
rect 5917 18377 5951 18411
rect 6561 18377 6595 18411
rect 7757 18377 7791 18411
rect 8033 18377 8067 18411
rect 10057 18377 10091 18411
rect 11161 18377 11195 18411
rect 11483 18377 11517 18411
rect 11897 18377 11931 18411
rect 13645 18377 13679 18411
rect 15393 18377 15427 18411
rect 5641 18241 5675 18275
rect 12449 18241 12483 18275
rect 14565 18241 14599 18275
rect 6837 18173 6871 18207
rect 9137 18173 9171 18207
rect 10425 18173 10459 18207
rect 11412 18173 11446 18207
rect 13369 18173 13403 18207
rect 14013 18173 14047 18207
rect 16129 18173 16163 18207
rect 16589 18173 16623 18207
rect 7158 18105 7192 18139
rect 8953 18105 8987 18139
rect 9458 18105 9492 18139
rect 12811 18105 12845 18139
rect 14289 18105 14323 18139
rect 14381 18105 14415 18139
rect 10793 18037 10827 18071
rect 12173 18037 12207 18071
rect 16681 18037 16715 18071
rect 7389 17833 7423 17867
rect 7665 17833 7699 17867
rect 8355 17833 8389 17867
rect 10609 17833 10643 17867
rect 11345 17833 11379 17867
rect 12817 17833 12851 17867
rect 13185 17833 13219 17867
rect 16221 17833 16255 17867
rect 6790 17765 6824 17799
rect 10051 17765 10085 17799
rect 12218 17765 12252 17799
rect 13829 17765 13863 17799
rect 14381 17765 14415 17799
rect 16681 17765 16715 17799
rect 5181 17697 5215 17731
rect 5365 17697 5399 17731
rect 8284 17697 8318 17731
rect 15368 17697 15402 17731
rect 5457 17629 5491 17663
rect 6469 17629 6503 17663
rect 9689 17629 9723 17663
rect 11897 17629 11931 17663
rect 13737 17629 13771 17663
rect 16589 17629 16623 17663
rect 18061 17629 18095 17663
rect 17141 17561 17175 17595
rect 9229 17493 9263 17527
rect 10977 17493 11011 17527
rect 15439 17493 15473 17527
rect 5273 17289 5307 17323
rect 6285 17289 6319 17323
rect 6653 17289 6687 17323
rect 7389 17289 7423 17323
rect 10149 17289 10183 17323
rect 10701 17289 10735 17323
rect 11897 17289 11931 17323
rect 13461 17289 13495 17323
rect 13691 17289 13725 17323
rect 14473 17289 14507 17323
rect 15393 17289 15427 17323
rect 4997 17221 5031 17255
rect 8217 17221 8251 17255
rect 8677 17221 8711 17255
rect 11437 17221 11471 17255
rect 10885 17153 10919 17187
rect 12587 17153 12621 17187
rect 16313 17153 16347 17187
rect 5768 17085 5802 17119
rect 5871 17085 5905 17119
rect 9045 17085 9079 17119
rect 9413 17085 9447 17119
rect 9597 17085 9631 17119
rect 12500 17085 12534 17119
rect 13604 17085 13638 17119
rect 14105 17085 14139 17119
rect 14632 17085 14666 17119
rect 17877 17085 17911 17119
rect 18153 17085 18187 17119
rect 7021 17017 7055 17051
rect 7665 17017 7699 17051
rect 7757 17017 7791 17051
rect 10977 17017 11011 17051
rect 16129 17017 16163 17051
rect 16405 17017 16439 17051
rect 16957 17017 16991 17051
rect 18061 17017 18095 17051
rect 9229 16949 9263 16983
rect 13001 16949 13035 16983
rect 14703 16949 14737 16983
rect 15761 16949 15795 16983
rect 17325 16949 17359 16983
rect 4353 16745 4387 16779
rect 6009 16745 6043 16779
rect 6469 16745 6503 16779
rect 9229 16745 9263 16779
rect 13599 16745 13633 16779
rect 13921 16745 13955 16779
rect 19855 16745 19889 16779
rect 5319 16677 5353 16711
rect 7573 16677 7607 16711
rect 8769 16677 8803 16711
rect 9873 16677 9907 16711
rect 11069 16677 11103 16711
rect 11713 16677 11747 16711
rect 11989 16677 12023 16711
rect 12081 16677 12115 16711
rect 15439 16677 15473 16711
rect 16681 16677 16715 16711
rect 16773 16677 16807 16711
rect 18245 16677 18279 16711
rect 18337 16677 18371 16711
rect 4169 16609 4203 16643
rect 5216 16609 5250 16643
rect 6193 16609 6227 16643
rect 6745 16609 6779 16643
rect 8033 16609 8067 16643
rect 8585 16609 8619 16643
rect 10333 16609 10367 16643
rect 10793 16609 10827 16643
rect 13496 16609 13530 16643
rect 15336 16609 15370 16643
rect 19752 16609 19786 16643
rect 12265 16541 12299 16575
rect 17325 16541 17359 16575
rect 17969 16541 18003 16575
rect 18521 16541 18555 16575
rect 12909 16405 12943 16439
rect 13369 16405 13403 16439
rect 15761 16405 15795 16439
rect 16221 16405 16255 16439
rect 5917 16201 5951 16235
rect 8493 16201 8527 16235
rect 10333 16201 10367 16235
rect 15163 16201 15197 16235
rect 15577 16201 15611 16235
rect 17049 16201 17083 16235
rect 17325 16201 17359 16235
rect 17877 16201 17911 16235
rect 9965 16133 9999 16167
rect 14473 16133 14507 16167
rect 15853 16133 15887 16167
rect 12541 16065 12575 16099
rect 18153 16065 18187 16099
rect 5273 15997 5307 16031
rect 5733 15997 5767 16031
rect 7297 15997 7331 16031
rect 7573 15997 7607 16031
rect 8953 15997 8987 16031
rect 9505 15997 9539 16031
rect 10517 15997 10551 16031
rect 11069 15997 11103 16031
rect 11529 15997 11563 16031
rect 14080 15997 14114 16031
rect 15092 15997 15126 16031
rect 16129 15997 16163 16031
rect 19717 15997 19751 16031
rect 7757 15929 7791 15963
rect 9689 15929 9723 15963
rect 12633 15929 12667 15963
rect 13185 15929 13219 15963
rect 16450 15929 16484 15963
rect 18245 15929 18279 15963
rect 18797 15929 18831 15963
rect 19625 15929 19659 15963
rect 4261 15861 4295 15895
rect 5641 15861 5675 15895
rect 6285 15861 6319 15895
rect 6653 15861 6687 15895
rect 8033 15861 8067 15895
rect 8769 15861 8803 15895
rect 10793 15861 10827 15895
rect 11989 15861 12023 15895
rect 13461 15861 13495 15895
rect 14151 15861 14185 15895
rect 19073 15861 19107 15895
rect 19441 15861 19475 15895
rect 6377 15657 6411 15691
rect 7113 15657 7147 15691
rect 9045 15657 9079 15691
rect 9873 15657 9907 15691
rect 10425 15657 10459 15691
rect 11713 15657 11747 15691
rect 13277 15657 13311 15691
rect 16497 15657 16531 15691
rect 16773 15657 16807 15691
rect 18337 15657 18371 15691
rect 18797 15657 18831 15691
rect 7843 15589 7877 15623
rect 10793 15589 10827 15623
rect 11345 15589 11379 15623
rect 12357 15589 12391 15623
rect 15939 15589 15973 15623
rect 17509 15589 17543 15623
rect 18981 15589 19015 15623
rect 19073 15589 19107 15623
rect 5917 15521 5951 15555
rect 6193 15521 6227 15555
rect 8401 15521 8435 15555
rect 13772 15521 13806 15555
rect 7481 15453 7515 15487
rect 10701 15453 10735 15487
rect 12081 15453 12115 15487
rect 12265 15453 12299 15487
rect 13875 15453 13909 15487
rect 15577 15453 15611 15487
rect 17417 15453 17451 15487
rect 6009 15385 6043 15419
rect 12817 15385 12851 15419
rect 17969 15385 18003 15419
rect 19533 15385 19567 15419
rect 15117 15317 15151 15351
rect 19993 15317 20027 15351
rect 7297 15113 7331 15147
rect 8953 15113 8987 15147
rect 10517 15113 10551 15147
rect 11253 15113 11287 15147
rect 13737 15113 13771 15147
rect 14841 15113 14875 15147
rect 15301 15113 15335 15147
rect 17509 15113 17543 15147
rect 18245 15113 18279 15147
rect 18981 15113 19015 15147
rect 21143 15113 21177 15147
rect 5917 15045 5951 15079
rect 9413 15045 9447 15079
rect 11529 15045 11563 15079
rect 13369 15045 13403 15079
rect 6193 14977 6227 15011
rect 7389 14977 7423 15011
rect 8585 14977 8619 15011
rect 9597 14977 9631 15011
rect 12173 14977 12207 15011
rect 12817 14977 12851 15011
rect 19533 14977 19567 15011
rect 19993 14977 20027 15011
rect 5733 14909 5767 14943
rect 11345 14909 11379 14943
rect 11805 14909 11839 14943
rect 14356 14909 14390 14943
rect 15485 14909 15519 14943
rect 15853 14909 15887 14943
rect 16221 14909 16255 14943
rect 16773 14909 16807 14943
rect 21040 14909 21074 14943
rect 21465 14909 21499 14943
rect 23708 14909 23742 14943
rect 24133 14909 24167 14943
rect 7751 14841 7785 14875
rect 9938 14841 9972 14875
rect 10885 14841 10919 14875
rect 12909 14841 12943 14875
rect 19349 14841 19383 14875
rect 19625 14841 19659 14875
rect 23811 14841 23845 14875
rect 5549 14773 5583 14807
rect 6653 14773 6687 14807
rect 8309 14773 8343 14807
rect 14427 14773 14461 14807
rect 15669 14773 15703 14807
rect 17233 14773 17267 14807
rect 18429 14773 18463 14807
rect 7481 14569 7515 14603
rect 10793 14569 10827 14603
rect 12725 14569 12759 14603
rect 15531 14569 15565 14603
rect 18981 14569 19015 14603
rect 7021 14501 7055 14535
rect 8033 14501 8067 14535
rect 9965 14501 9999 14535
rect 11707 14501 11741 14535
rect 13455 14501 13489 14535
rect 19349 14501 19383 14535
rect 19441 14501 19475 14535
rect 19993 14501 20027 14535
rect 21097 14501 21131 14535
rect 5273 14433 5307 14467
rect 6561 14433 6595 14467
rect 6837 14433 6871 14467
rect 13093 14433 13127 14467
rect 15428 14433 15462 14467
rect 16589 14433 16623 14467
rect 16865 14433 16899 14467
rect 17233 14433 17267 14467
rect 17601 14433 17635 14467
rect 7941 14365 7975 14399
rect 8861 14365 8895 14399
rect 9873 14365 9907 14399
rect 10517 14365 10551 14399
rect 11345 14365 11379 14399
rect 16313 14365 16347 14399
rect 17877 14365 17911 14399
rect 21005 14365 21039 14399
rect 21281 14365 21315 14399
rect 8493 14297 8527 14331
rect 5457 14229 5491 14263
rect 6009 14229 6043 14263
rect 9229 14229 9263 14263
rect 11161 14229 11195 14263
rect 12265 14229 12299 14263
rect 14013 14229 14047 14263
rect 14749 14229 14783 14263
rect 15117 14229 15151 14263
rect 15945 14229 15979 14263
rect 4169 14025 4203 14059
rect 6377 14025 6411 14059
rect 7113 14025 7147 14059
rect 8677 14025 8711 14059
rect 9045 14025 9079 14059
rect 10241 14025 10275 14059
rect 10609 14025 10643 14059
rect 15025 14025 15059 14059
rect 17785 14025 17819 14059
rect 18981 14025 19015 14059
rect 19257 14025 19291 14059
rect 19625 14025 19659 14059
rect 21189 14025 21223 14059
rect 9321 13957 9355 13991
rect 11437 13957 11471 13991
rect 14749 13957 14783 13991
rect 7757 13889 7791 13923
rect 8401 13889 8435 13923
rect 9689 13889 9723 13923
rect 10885 13889 10919 13923
rect 12265 13889 12299 13923
rect 13001 13889 13035 13923
rect 20269 13889 20303 13923
rect 4445 13821 4479 13855
rect 5365 13821 5399 13855
rect 7573 13821 7607 13855
rect 9229 13821 9263 13855
rect 9505 13821 9539 13855
rect 15485 13821 15519 13855
rect 15853 13821 15887 13855
rect 16037 13821 16071 13855
rect 16497 13821 16531 13855
rect 17325 13821 17359 13855
rect 18061 13821 18095 13855
rect 20085 13821 20119 13855
rect 20913 13821 20947 13855
rect 21557 13821 21591 13855
rect 4353 13753 4387 13787
rect 7849 13753 7883 13787
rect 10977 13753 11011 13787
rect 12725 13753 12759 13787
rect 12817 13753 12851 13787
rect 18382 13753 18416 13787
rect 20361 13753 20395 13787
rect 11805 13685 11839 13719
rect 13645 13685 13679 13719
rect 14381 13685 14415 13719
rect 15301 13685 15335 13719
rect 17049 13685 17083 13719
rect 9781 13481 9815 13515
rect 10333 13481 10367 13515
rect 12449 13481 12483 13515
rect 13553 13481 13587 13515
rect 14381 13481 14415 13515
rect 19901 13481 19935 13515
rect 20269 13481 20303 13515
rect 11155 13413 11189 13447
rect 12725 13413 12759 13447
rect 17785 13413 17819 13447
rect 18061 13413 18095 13447
rect 18934 13413 18968 13447
rect 20913 13413 20947 13447
rect 4813 13345 4847 13379
rect 5089 13345 5123 13379
rect 7297 13345 7331 13379
rect 8585 13345 8619 13379
rect 14197 13345 14231 13379
rect 16221 13345 16255 13379
rect 16589 13345 16623 13379
rect 16773 13345 16807 13379
rect 17141 13345 17175 13379
rect 17509 13345 17543 13379
rect 18613 13345 18647 13379
rect 19533 13345 19567 13379
rect 21005 13345 21039 13379
rect 4905 13277 4939 13311
rect 5457 13277 5491 13311
rect 10793 13277 10827 13311
rect 12633 13277 12667 13311
rect 12909 13277 12943 13311
rect 15025 13277 15059 13311
rect 6929 13209 6963 13243
rect 9229 13209 9263 13243
rect 13921 13209 13955 13243
rect 15485 13209 15519 13243
rect 7481 13141 7515 13175
rect 8125 13141 8159 13175
rect 8493 13141 8527 13175
rect 8769 13141 8803 13175
rect 11713 13141 11747 13175
rect 11989 13141 12023 13175
rect 14657 13141 14691 13175
rect 4261 12937 4295 12971
rect 5825 12937 5859 12971
rect 7113 12937 7147 12971
rect 8769 12937 8803 12971
rect 10149 12937 10183 12971
rect 11805 12937 11839 12971
rect 17417 12937 17451 12971
rect 18245 12937 18279 12971
rect 18705 12937 18739 12971
rect 18935 12937 18969 12971
rect 21005 12937 21039 12971
rect 12265 12869 12299 12903
rect 8309 12801 8343 12835
rect 9781 12801 9815 12835
rect 11069 12801 11103 12835
rect 12541 12801 12575 12835
rect 12817 12801 12851 12835
rect 13461 12801 13495 12835
rect 19257 12801 19291 12835
rect 19993 12801 20027 12835
rect 20637 12801 20671 12835
rect 2421 12733 2455 12767
rect 3433 12733 3467 12767
rect 4537 12733 4571 12767
rect 5457 12733 5491 12767
rect 7757 12733 7791 12767
rect 7849 12733 7883 12767
rect 8033 12733 8067 12767
rect 9321 12733 9355 12767
rect 10333 12733 10367 12767
rect 10793 12733 10827 12767
rect 14381 12733 14415 12767
rect 14841 12733 14875 12767
rect 15301 12733 15335 12767
rect 15577 12733 15611 12767
rect 17049 12733 17083 12767
rect 18864 12733 18898 12767
rect 21500 12733 21534 12767
rect 21925 12733 21959 12767
rect 22512 12733 22546 12767
rect 22937 12733 22971 12767
rect 2881 12665 2915 12699
rect 5181 12665 5215 12699
rect 7573 12665 7607 12699
rect 12633 12665 12667 12699
rect 15853 12665 15887 12699
rect 20085 12665 20119 12699
rect 2605 12597 2639 12631
rect 3617 12597 3651 12631
rect 3985 12597 4019 12631
rect 6193 12597 6227 12631
rect 9505 12597 9539 12631
rect 11345 12597 11379 12631
rect 13829 12597 13863 12631
rect 14197 12597 14231 12631
rect 16313 12597 16347 12631
rect 16681 12597 16715 12631
rect 19809 12597 19843 12631
rect 21603 12597 21637 12631
rect 22615 12597 22649 12631
rect 5273 12393 5307 12427
rect 12081 12393 12115 12427
rect 24777 12393 24811 12427
rect 7573 12325 7607 12359
rect 12817 12325 12851 12359
rect 19118 12325 19152 12359
rect 21097 12325 21131 12359
rect 2329 12257 2363 12291
rect 2421 12257 2455 12291
rect 2697 12257 2731 12291
rect 4721 12257 4755 12291
rect 4813 12257 4847 12291
rect 4905 12257 4939 12291
rect 5089 12257 5123 12291
rect 6377 12257 6411 12291
rect 7205 12257 7239 12291
rect 8217 12257 8251 12291
rect 9965 12257 9999 12291
rect 10425 12257 10459 12291
rect 11564 12257 11598 12291
rect 12909 12257 12943 12291
rect 13369 12257 13403 12291
rect 13737 12257 13771 12291
rect 14105 12257 14139 12291
rect 15301 12257 15335 12291
rect 15761 12257 15795 12291
rect 16313 12257 16347 12291
rect 16773 12257 16807 12291
rect 17141 12257 17175 12291
rect 17509 12257 17543 12291
rect 18797 12257 18831 12291
rect 22512 12257 22546 12291
rect 2881 12189 2915 12223
rect 10701 12189 10735 12223
rect 10977 12189 11011 12223
rect 11437 12189 11471 12223
rect 16129 12189 16163 12223
rect 21005 12189 21039 12223
rect 21281 12189 21315 12223
rect 21925 12189 21959 12223
rect 2513 12121 2547 12155
rect 8769 12121 8803 12155
rect 14289 12121 14323 12155
rect 17693 12121 17727 12155
rect 6561 12053 6595 12087
rect 11667 12053 11701 12087
rect 12449 12053 12483 12087
rect 14657 12053 14691 12087
rect 15485 12053 15519 12087
rect 19717 12053 19751 12087
rect 22615 12053 22649 12087
rect 1961 11849 1995 11883
rect 2605 11849 2639 11883
rect 4169 11849 4203 11883
rect 4445 11849 4479 11883
rect 6101 11849 6135 11883
rect 6377 11849 6411 11883
rect 8309 11849 8343 11883
rect 8585 11849 8619 11883
rect 10057 11849 10091 11883
rect 11805 11849 11839 11883
rect 12725 11849 12759 11883
rect 14197 11849 14231 11883
rect 18429 11849 18463 11883
rect 18705 11849 18739 11883
rect 20637 11849 20671 11883
rect 4721 11781 4755 11815
rect 7113 11781 7147 11815
rect 7297 11781 7331 11815
rect 8861 11781 8895 11815
rect 17509 11781 17543 11815
rect 5365 11713 5399 11747
rect 7941 11713 7975 11747
rect 15853 11713 15887 11747
rect 18889 11713 18923 11747
rect 20085 11713 20119 11747
rect 2053 11645 2087 11679
rect 3157 11645 3191 11679
rect 3801 11645 3835 11679
rect 4629 11645 4663 11679
rect 4905 11645 4939 11679
rect 7205 11645 7239 11679
rect 7481 11645 7515 11679
rect 8769 11645 8803 11679
rect 9045 11645 9079 11679
rect 11437 11645 11471 11679
rect 13461 11645 13495 11679
rect 13921 11645 13955 11679
rect 14657 11645 14691 11679
rect 14841 11645 14875 11679
rect 15393 11645 15427 11679
rect 15761 11645 15795 11679
rect 16681 11645 16715 11679
rect 17141 11645 17175 11679
rect 19809 11645 19843 11679
rect 5641 11577 5675 11611
rect 9505 11577 9539 11611
rect 13553 11577 13587 11611
rect 16313 11577 16347 11611
rect 19210 11577 19244 11611
rect 21465 11577 21499 11611
rect 21557 11577 21591 11611
rect 22109 11577 22143 11611
rect 2237 11509 2271 11543
rect 2881 11509 2915 11543
rect 10333 11509 10367 11543
rect 11069 11509 11103 11543
rect 12173 11509 12207 11543
rect 16865 11509 16899 11543
rect 20913 11509 20947 11543
rect 22477 11509 22511 11543
rect 2053 11305 2087 11339
rect 4721 11305 4755 11339
rect 6745 11305 6779 11339
rect 7941 11305 7975 11339
rect 9045 11305 9079 11339
rect 10149 11305 10183 11339
rect 12081 11305 12115 11339
rect 12449 11305 12483 11339
rect 14473 11305 14507 11339
rect 15761 11305 15795 11339
rect 16313 11305 16347 11339
rect 18797 11305 18831 11339
rect 21373 11305 21407 11339
rect 7389 11237 7423 11271
rect 19993 11237 20027 11271
rect 21925 11237 21959 11271
rect 22477 11237 22511 11271
rect 2421 11169 2455 11203
rect 2513 11169 2547 11203
rect 2697 11169 2731 11203
rect 4997 11169 5031 11203
rect 5273 11169 5307 11203
rect 6561 11169 6595 11203
rect 7021 11169 7055 11203
rect 8033 11169 8067 11203
rect 8493 11169 8527 11203
rect 10057 11169 10091 11203
rect 10333 11169 10367 11203
rect 10701 11169 10735 11203
rect 11069 11169 11103 11203
rect 12173 11169 12207 11203
rect 12909 11169 12943 11203
rect 13001 11169 13035 11203
rect 13553 11169 13587 11203
rect 15301 11169 15335 11203
rect 16497 11169 16531 11203
rect 16957 11169 16991 11203
rect 17325 11169 17359 11203
rect 17693 11169 17727 11203
rect 19533 11169 19567 11203
rect 24352 11169 24386 11203
rect 3157 11101 3191 11135
rect 5733 11101 5767 11135
rect 8769 11101 8803 11135
rect 21833 11101 21867 11135
rect 23305 11101 23339 11135
rect 5089 11033 5123 11067
rect 15485 11033 15519 11067
rect 17877 11033 17911 11067
rect 14013 10965 14047 10999
rect 14749 10965 14783 10999
rect 24455 10965 24489 10999
rect 2053 10761 2087 10795
rect 2329 10761 2363 10795
rect 2973 10761 3007 10795
rect 3341 10761 3375 10795
rect 8033 10761 8067 10795
rect 9505 10761 9539 10795
rect 11805 10761 11839 10795
rect 12265 10761 12299 10795
rect 12725 10761 12759 10795
rect 13185 10761 13219 10795
rect 18245 10761 18279 10795
rect 19809 10761 19843 10795
rect 20177 10761 20211 10795
rect 21465 10761 21499 10795
rect 21833 10761 21867 10795
rect 24777 10761 24811 10795
rect 3709 10693 3743 10727
rect 15301 10693 15335 10727
rect 8493 10625 8527 10659
rect 8769 10625 8803 10659
rect 10425 10625 10459 10659
rect 17417 10625 17451 10659
rect 20453 10625 20487 10659
rect 21097 10625 21131 10659
rect 21925 10625 21959 10659
rect 2513 10557 2547 10591
rect 3525 10557 3559 10591
rect 4905 10557 4939 10591
rect 5917 10557 5951 10591
rect 6561 10557 6595 10591
rect 6837 10557 6871 10591
rect 6929 10557 6963 10591
rect 7113 10557 7147 10591
rect 13369 10557 13403 10591
rect 13829 10557 13863 10591
rect 14197 10557 14231 10591
rect 14565 10557 14599 10591
rect 15669 10557 15703 10591
rect 16129 10557 16163 10591
rect 16681 10557 16715 10591
rect 16957 10557 16991 10591
rect 18705 10557 18739 10591
rect 18889 10557 18923 10591
rect 22017 10557 22051 10591
rect 24317 10557 24351 10591
rect 24593 10557 24627 10591
rect 25145 10557 25179 10591
rect 5273 10489 5307 10523
rect 8585 10489 8619 10523
rect 10333 10489 10367 10523
rect 10787 10489 10821 10523
rect 14841 10489 14875 10523
rect 17785 10489 17819 10523
rect 20545 10489 20579 10523
rect 2697 10421 2731 10455
rect 4077 10421 4111 10455
rect 4445 10421 4479 10455
rect 5549 10421 5583 10455
rect 7297 10421 7331 10455
rect 9873 10421 9907 10455
rect 11345 10421 11379 10455
rect 16865 10421 16899 10455
rect 19073 10421 19107 10455
rect 4905 10217 4939 10251
rect 7941 10217 7975 10251
rect 10885 10217 10919 10251
rect 12633 10217 12667 10251
rect 13645 10217 13679 10251
rect 15025 10217 15059 10251
rect 15853 10217 15887 10251
rect 20453 10217 20487 10251
rect 22017 10217 22051 10251
rect 5733 10149 5767 10183
rect 8125 10149 8159 10183
rect 8217 10149 8251 10183
rect 10517 10149 10551 10183
rect 11345 10149 11379 10183
rect 11897 10149 11931 10183
rect 13087 10149 13121 10183
rect 13921 10149 13955 10183
rect 16221 10149 16255 10183
rect 19026 10149 19060 10183
rect 21097 10149 21131 10183
rect 2421 10081 2455 10115
rect 2697 10081 2731 10115
rect 3157 10081 3191 10115
rect 4997 10081 5031 10115
rect 5273 10081 5307 10115
rect 6561 10081 6595 10115
rect 9689 10081 9723 10115
rect 10149 10081 10183 10115
rect 12725 10081 12759 10115
rect 16405 10081 16439 10115
rect 16865 10081 16899 10115
rect 17233 10081 17267 10115
rect 17601 10081 17635 10115
rect 18705 10081 18739 10115
rect 23156 10081 23190 10115
rect 4537 10013 4571 10047
rect 8401 10013 8435 10047
rect 11253 10013 11287 10047
rect 15301 10013 15335 10047
rect 17877 10013 17911 10047
rect 21005 10013 21039 10047
rect 21649 10013 21683 10047
rect 2513 9945 2547 9979
rect 5089 9945 5123 9979
rect 6745 9945 6779 9979
rect 7021 9877 7055 9911
rect 7481 9877 7515 9911
rect 9045 9877 9079 9911
rect 9873 9877 9907 9911
rect 12173 9877 12207 9911
rect 19625 9877 19659 9911
rect 23259 9877 23293 9911
rect 2145 9673 2179 9707
rect 6653 9673 6687 9707
rect 9781 9673 9815 9707
rect 11897 9673 11931 9707
rect 15485 9673 15519 9707
rect 17325 9673 17359 9707
rect 18981 9673 19015 9707
rect 23121 9673 23155 9707
rect 2881 9605 2915 9639
rect 3985 9605 4019 9639
rect 9137 9605 9171 9639
rect 9505 9605 9539 9639
rect 10701 9605 10735 9639
rect 13829 9605 13863 9639
rect 14657 9605 14691 9639
rect 15853 9605 15887 9639
rect 17049 9605 17083 9639
rect 19625 9605 19659 9639
rect 20821 9605 20855 9639
rect 22385 9605 22419 9639
rect 24777 9605 24811 9639
rect 3341 9537 3375 9571
rect 5181 9537 5215 9571
rect 5549 9537 5583 9571
rect 12541 9537 12575 9571
rect 13001 9537 13035 9571
rect 14105 9537 14139 9571
rect 18061 9537 18095 9571
rect 19257 9537 19291 9571
rect 20177 9537 20211 9571
rect 21465 9537 21499 9571
rect 21741 9537 21775 9571
rect 3617 9469 3651 9503
rect 4537 9469 4571 9503
rect 5089 9469 5123 9503
rect 5365 9469 5399 9503
rect 6101 9469 6135 9503
rect 7573 9469 7607 9503
rect 9321 9469 9355 9503
rect 10149 9469 10183 9503
rect 24593 9469 24627 9503
rect 25145 9469 25179 9503
rect 7935 9401 7969 9435
rect 10885 9401 10919 9435
rect 10977 9401 11011 9435
rect 11529 9401 11563 9435
rect 12633 9401 12667 9435
rect 14197 9401 14231 9435
rect 15117 9401 15151 9435
rect 16037 9401 16071 9435
rect 16129 9401 16163 9435
rect 16681 9401 16715 9435
rect 17877 9401 17911 9435
rect 18423 9401 18457 9435
rect 19901 9401 19935 9435
rect 19993 9401 20027 9435
rect 21557 9401 21591 9435
rect 2513 9333 2547 9367
rect 4905 9333 4939 9367
rect 7021 9333 7055 9367
rect 7481 9333 7515 9367
rect 8493 9333 8527 9367
rect 8769 9333 8803 9367
rect 12265 9333 12299 9367
rect 13553 9333 13587 9367
rect 21281 9333 21315 9367
rect 5549 9129 5583 9163
rect 6285 9129 6319 9163
rect 7205 9129 7239 9163
rect 8493 9129 8527 9163
rect 11345 9129 11379 9163
rect 13277 9129 13311 9163
rect 14013 9129 14047 9163
rect 14381 9129 14415 9163
rect 15117 9129 15151 9163
rect 16221 9129 16255 9163
rect 16589 9129 16623 9163
rect 18061 9129 18095 9163
rect 18613 9129 18647 9163
rect 23719 9129 23753 9163
rect 5273 9061 5307 9095
rect 5917 9061 5951 9095
rect 7935 9061 7969 9095
rect 8861 9061 8895 9095
rect 10746 9061 10780 9095
rect 12449 9061 12483 9095
rect 13001 9061 13035 9095
rect 15663 9061 15697 9095
rect 18889 9061 18923 9095
rect 18981 9061 19015 9095
rect 19533 9061 19567 9095
rect 21097 9061 21131 9095
rect 4629 8993 4663 9027
rect 6101 8993 6135 9027
rect 10333 8993 10367 9027
rect 13829 8993 13863 9027
rect 15301 8993 15335 9027
rect 17141 8993 17175 9027
rect 23616 8993 23650 9027
rect 7573 8925 7607 8959
rect 10425 8925 10459 8959
rect 12357 8925 12391 8959
rect 17049 8925 17083 8959
rect 21005 8925 21039 8959
rect 21281 8925 21315 8959
rect 21925 8925 21959 8959
rect 11621 8857 11655 8891
rect 12173 8857 12207 8891
rect 19809 8789 19843 8823
rect 4077 8585 4111 8619
rect 4445 8585 4479 8619
rect 8677 8585 8711 8619
rect 13369 8585 13403 8619
rect 13737 8585 13771 8619
rect 15393 8585 15427 8619
rect 17141 8585 17175 8619
rect 18613 8585 18647 8619
rect 19257 8585 19291 8619
rect 19717 8585 19751 8619
rect 21649 8585 21683 8619
rect 23857 8585 23891 8619
rect 5089 8517 5123 8551
rect 6009 8517 6043 8551
rect 10241 8517 10275 8551
rect 16681 8517 16715 8551
rect 20913 8517 20947 8551
rect 5733 8449 5767 8483
rect 6377 8449 6411 8483
rect 9873 8449 9907 8483
rect 11621 8449 11655 8483
rect 13829 8449 13863 8483
rect 15945 8449 15979 8483
rect 18797 8449 18831 8483
rect 19901 8449 19935 8483
rect 20545 8449 20579 8483
rect 4813 8381 4847 8415
rect 4997 8381 5031 8415
rect 5227 8381 5261 8415
rect 7389 8381 7423 8415
rect 7573 8381 7607 8415
rect 8861 8381 8895 8415
rect 9321 8381 9355 8415
rect 10425 8381 10459 8415
rect 11345 8381 11379 8415
rect 12173 8381 12207 8415
rect 12449 8381 12483 8415
rect 12909 8381 12943 8415
rect 14749 8381 14783 8415
rect 21465 8381 21499 8415
rect 24409 8381 24443 8415
rect 24961 8381 24995 8415
rect 7849 8313 7883 8347
rect 9597 8313 9631 8347
rect 10746 8313 10780 8347
rect 14191 8313 14225 8347
rect 16129 8313 16163 8347
rect 16221 8313 16255 8347
rect 19993 8313 20027 8347
rect 8125 8245 8159 8279
rect 12633 8245 12667 8279
rect 24593 8245 24627 8279
rect 6009 8041 6043 8075
rect 7573 8041 7607 8075
rect 7849 8041 7883 8075
rect 10057 8041 10091 8075
rect 10885 8041 10919 8075
rect 12909 8041 12943 8075
rect 14657 8041 14691 8075
rect 15025 8041 15059 8075
rect 19487 8041 19521 8075
rect 21373 8041 21407 8075
rect 21741 8041 21775 8075
rect 24777 8041 24811 8075
rect 11253 7973 11287 8007
rect 11437 7973 11471 8007
rect 11529 7973 11563 8007
rect 13829 7973 13863 8007
rect 15485 7973 15519 8007
rect 16037 7973 16071 8007
rect 17922 7973 17956 8007
rect 5181 7905 5215 7939
rect 5365 7905 5399 7939
rect 6469 7905 6503 7939
rect 7021 7905 7055 7939
rect 8217 7905 8251 7939
rect 8585 7905 8619 7939
rect 9781 7905 9815 7939
rect 10241 7905 10275 7939
rect 17601 7905 17635 7939
rect 19416 7905 19450 7939
rect 20980 7905 21014 7939
rect 24593 7905 24627 7939
rect 5457 7837 5491 7871
rect 7205 7837 7239 7871
rect 8769 7837 8803 7871
rect 11713 7837 11747 7871
rect 13737 7837 13771 7871
rect 15393 7837 15427 7871
rect 12449 7769 12483 7803
rect 14289 7769 14323 7803
rect 16313 7769 16347 7803
rect 18521 7769 18555 7803
rect 9229 7701 9263 7735
rect 18889 7701 18923 7735
rect 19901 7701 19935 7735
rect 21051 7701 21085 7735
rect 4721 7497 4755 7531
rect 6561 7497 6595 7531
rect 8677 7497 8711 7531
rect 8953 7497 8987 7531
rect 10149 7497 10183 7531
rect 11713 7497 11747 7531
rect 14519 7497 14553 7531
rect 16773 7497 16807 7531
rect 18245 7497 18279 7531
rect 20499 7497 20533 7531
rect 21189 7497 21223 7531
rect 24731 7497 24765 7531
rect 25421 7497 25455 7531
rect 10517 7429 10551 7463
rect 14105 7429 14139 7463
rect 4997 7361 5031 7395
rect 9229 7361 9263 7395
rect 9689 7361 9723 7395
rect 11253 7361 11287 7395
rect 12449 7361 12483 7395
rect 14933 7361 14967 7395
rect 15485 7361 15519 7395
rect 15945 7361 15979 7395
rect 16957 7361 16991 7395
rect 17693 7361 17727 7395
rect 18889 7361 18923 7395
rect 3709 7293 3743 7327
rect 4169 7293 4203 7327
rect 5457 7293 5491 7327
rect 5641 7293 5675 7327
rect 7389 7293 7423 7327
rect 10701 7293 10735 7327
rect 11161 7293 11195 7327
rect 13369 7293 13403 7327
rect 14448 7293 14482 7327
rect 20396 7293 20430 7327
rect 20821 7293 20855 7327
rect 24660 7293 24694 7327
rect 25053 7293 25087 7327
rect 3525 7225 3559 7259
rect 5917 7225 5951 7259
rect 7710 7225 7744 7259
rect 9321 7225 9355 7259
rect 12811 7225 12845 7259
rect 13645 7225 13679 7259
rect 15577 7225 15611 7259
rect 18705 7225 18739 7259
rect 18981 7225 19015 7259
rect 19533 7225 19567 7259
rect 3893 7157 3927 7191
rect 7205 7157 7239 7191
rect 8309 7157 8343 7191
rect 12173 7157 12207 7191
rect 15301 7157 15335 7191
rect 16405 7157 16439 7191
rect 19901 7157 19935 7191
rect 3709 6953 3743 6987
rect 6469 6953 6503 6987
rect 8125 6953 8159 6987
rect 9137 6953 9171 6987
rect 10793 6953 10827 6987
rect 11161 6953 11195 6987
rect 4997 6885 5031 6919
rect 7250 6885 7284 6919
rect 9873 6885 9907 6919
rect 11615 6885 11649 6919
rect 13185 6885 13219 6919
rect 15485 6885 15519 6919
rect 16037 6885 16071 6919
rect 17227 6885 17261 6919
rect 18797 6885 18831 6919
rect 5457 6817 5491 6851
rect 5825 6817 5859 6851
rect 6929 6817 6963 6851
rect 8493 6817 8527 6851
rect 11253 6817 11287 6851
rect 12541 6817 12575 6851
rect 16865 6817 16899 6851
rect 21005 6817 21039 6851
rect 6101 6749 6135 6783
rect 9781 6749 9815 6783
rect 10149 6749 10183 6783
rect 13093 6749 13127 6783
rect 13369 6749 13403 6783
rect 15393 6749 15427 6783
rect 18705 6749 18739 6783
rect 18981 6749 19015 6783
rect 20913 6749 20947 6783
rect 7849 6613 7883 6647
rect 12173 6613 12207 6647
rect 14289 6613 14323 6647
rect 15025 6613 15059 6647
rect 17785 6613 17819 6647
rect 18061 6613 18095 6647
rect 19625 6613 19659 6647
rect 5089 6409 5123 6443
rect 6193 6409 6227 6443
rect 6653 6409 6687 6443
rect 9045 6409 9079 6443
rect 9413 6409 9447 6443
rect 10425 6409 10459 6443
rect 11529 6409 11563 6443
rect 13645 6409 13679 6443
rect 15393 6409 15427 6443
rect 17417 6409 17451 6443
rect 21005 6409 21039 6443
rect 19073 6341 19107 6375
rect 19441 6341 19475 6375
rect 24777 6341 24811 6375
rect 7757 6273 7791 6307
rect 10609 6273 10643 6307
rect 12449 6273 12483 6307
rect 14289 6273 14323 6307
rect 14565 6273 14599 6307
rect 15669 6273 15703 6307
rect 17141 6273 17175 6307
rect 18797 6273 18831 6307
rect 19993 6273 20027 6307
rect 4721 6205 4755 6239
rect 5457 6205 5491 6239
rect 5641 6205 5675 6239
rect 5917 6205 5951 6239
rect 8677 6205 8711 6239
rect 9572 6205 9606 6239
rect 13369 6205 13403 6239
rect 14013 6205 14047 6239
rect 16313 6205 16347 6239
rect 16497 6205 16531 6239
rect 17785 6205 17819 6239
rect 24593 6205 24627 6239
rect 25145 6205 25179 6239
rect 8078 6137 8112 6171
rect 10930 6137 10964 6171
rect 11805 6137 11839 6171
rect 12173 6137 12207 6171
rect 12770 6137 12804 6171
rect 14381 6137 14415 6171
rect 18153 6137 18187 6171
rect 18245 6137 18279 6171
rect 19717 6137 19751 6171
rect 19809 6137 19843 6171
rect 7113 6069 7147 6103
rect 7573 6069 7607 6103
rect 9643 6069 9677 6103
rect 10057 6069 10091 6103
rect 5273 5865 5307 5899
rect 8309 5865 8343 5899
rect 8723 5865 8757 5899
rect 9137 5865 9171 5899
rect 11253 5865 11287 5899
rect 14013 5865 14047 5899
rect 14335 5865 14369 5899
rect 16865 5865 16899 5899
rect 7107 5797 7141 5831
rect 8033 5797 8067 5831
rect 9873 5797 9907 5831
rect 12633 5797 12667 5831
rect 12725 5797 12759 5831
rect 15301 5797 15335 5831
rect 17785 5797 17819 5831
rect 19349 5797 19383 5831
rect 6745 5729 6779 5763
rect 7665 5729 7699 5763
rect 8652 5729 8686 5763
rect 14264 5729 14298 5763
rect 15485 5729 15519 5763
rect 9781 5661 9815 5695
rect 10057 5661 10091 5695
rect 11437 5661 11471 5695
rect 13645 5661 13679 5695
rect 17693 5661 17727 5695
rect 18337 5661 18371 5695
rect 19257 5661 19291 5695
rect 19533 5661 19567 5695
rect 10885 5593 10919 5627
rect 13185 5593 13219 5627
rect 18613 5525 18647 5559
rect 6193 5321 6227 5355
rect 7113 5321 7147 5355
rect 8677 5321 8711 5355
rect 9965 5321 9999 5355
rect 11805 5321 11839 5355
rect 13829 5321 13863 5355
rect 15025 5321 15059 5355
rect 15485 5321 15519 5355
rect 17095 5321 17129 5355
rect 19257 5321 19291 5355
rect 19533 5321 19567 5355
rect 24731 5321 24765 5355
rect 9597 5253 9631 5287
rect 12081 5253 12115 5287
rect 13093 5253 13127 5287
rect 9045 5185 9079 5219
rect 10701 5185 10735 5219
rect 10885 5185 10919 5219
rect 6653 5049 6687 5083
rect 7481 5049 7515 5083
rect 7573 5049 7607 5083
rect 8125 5049 8159 5083
rect 9137 5049 9171 5083
rect 10977 5049 11011 5083
rect 11529 5049 11563 5083
rect 12541 5185 12575 5219
rect 13461 5185 13495 5219
rect 14105 5185 14139 5219
rect 14381 5185 14415 5219
rect 17417 5185 17451 5219
rect 17785 5185 17819 5219
rect 18061 5185 18095 5219
rect 15612 5117 15646 5151
rect 16037 5117 16071 5151
rect 17024 5117 17058 5151
rect 24660 5117 24694 5151
rect 12633 5049 12667 5083
rect 14197 5049 14231 5083
rect 12081 4981 12115 5015
rect 12173 4981 12207 5015
rect 15715 4981 15749 5015
rect 16773 4981 16807 5015
rect 25145 4981 25179 5015
rect 6377 4777 6411 4811
rect 9045 4777 9079 4811
rect 10149 4777 10183 4811
rect 13277 4777 13311 4811
rect 17831 4777 17865 4811
rect 24777 4777 24811 4811
rect 7573 4709 7607 4743
rect 8125 4709 8159 4743
rect 10885 4709 10919 4743
rect 11437 4709 11471 4743
rect 12449 4709 12483 4743
rect 13001 4709 13035 4743
rect 9756 4641 9790 4675
rect 13880 4641 13914 4675
rect 15761 4641 15795 4675
rect 17728 4641 17762 4675
rect 24593 4641 24627 4675
rect 7481 4573 7515 4607
rect 10793 4573 10827 4607
rect 12357 4573 12391 4607
rect 13967 4573 14001 4607
rect 9827 4437 9861 4471
rect 15945 4437 15979 4471
rect 9873 4233 9907 4267
rect 10701 4233 10735 4267
rect 11897 4233 11931 4267
rect 13921 4233 13955 4267
rect 15761 4233 15795 4267
rect 17693 4233 17727 4267
rect 24593 4233 24627 4267
rect 9505 4165 9539 4199
rect 6653 4097 6687 4131
rect 8033 4097 8067 4131
rect 8309 4097 8343 4131
rect 8677 4097 8711 4131
rect 8953 4097 8987 4131
rect 11529 4097 11563 4131
rect 13185 4097 13219 4131
rect 12173 4029 12207 4063
rect 14448 4029 14482 4063
rect 20269 4029 20303 4063
rect 20821 4029 20855 4063
rect 7389 3961 7423 3995
rect 7481 3961 7515 3995
rect 9045 3961 9079 3995
rect 10885 3961 10919 3995
rect 10977 3961 11011 3995
rect 12541 3961 12575 3995
rect 12633 3961 12667 3995
rect 7205 3893 7239 3927
rect 10241 3893 10275 3927
rect 14519 3893 14553 3927
rect 14933 3893 14967 3927
rect 20453 3893 20487 3927
rect 2375 3689 2409 3723
rect 5503 3689 5537 3723
rect 6515 3689 6549 3723
rect 7297 3689 7331 3723
rect 8953 3689 8987 3723
rect 11161 3689 11195 3723
rect 11851 3689 11885 3723
rect 12449 3689 12483 3723
rect 7573 3621 7607 3655
rect 8125 3621 8159 3655
rect 9781 3621 9815 3655
rect 9873 3621 9907 3655
rect 12817 3621 12851 3655
rect 2304 3553 2338 3587
rect 5432 3553 5466 3587
rect 6412 3553 6446 3587
rect 10885 3553 10919 3587
rect 11780 3553 11814 3587
rect 21649 3553 21683 3587
rect 7481 3485 7515 3519
rect 10057 3485 10091 3519
rect 21833 3417 21867 3451
rect 6975 3145 7009 3179
rect 8033 3145 8067 3179
rect 9505 3145 9539 3179
rect 10517 3145 10551 3179
rect 11805 3145 11839 3179
rect 21741 3145 21775 3179
rect 22109 3145 22143 3179
rect 7757 3077 7791 3111
rect 10149 3077 10183 3111
rect 18245 3077 18279 3111
rect 6904 2941 6938 2975
rect 7297 2941 7331 2975
rect 9724 2941 9758 2975
rect 13588 2941 13622 2975
rect 14013 2941 14047 2975
rect 18061 2941 18095 2975
rect 18613 2941 18647 2975
rect 21189 2941 21223 2975
rect 24317 2941 24351 2975
rect 24869 2941 24903 2975
rect 9827 2873 9861 2907
rect 13691 2873 13725 2907
rect 2329 2805 2363 2839
rect 5457 2805 5491 2839
rect 6377 2805 6411 2839
rect 21373 2805 21407 2839
rect 24501 2805 24535 2839
rect 1547 2601 1581 2635
rect 4583 2601 4617 2635
rect 7159 2601 7193 2635
rect 10011 2601 10045 2635
rect 11023 2601 11057 2635
rect 16727 2601 16761 2635
rect 18981 2601 19015 2635
rect 20085 2601 20119 2635
rect 21925 2601 21959 2635
rect 1444 2465 1478 2499
rect 1869 2465 1903 2499
rect 4512 2465 4546 2499
rect 7088 2465 7122 2499
rect 9908 2465 9942 2499
rect 10333 2465 10367 2499
rect 10952 2465 10986 2499
rect 16656 2465 16690 2499
rect 18337 2465 18371 2499
rect 19441 2465 19475 2499
rect 21741 2465 21775 2499
rect 22293 2465 22327 2499
rect 22845 2465 22879 2499
rect 23397 2465 23431 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 4905 2397 4939 2431
rect 18521 2329 18555 2363
rect 19625 2329 19659 2363
rect 23029 2329 23063 2363
rect 7573 2261 7607 2295
rect 11437 2261 11471 2295
rect 17049 2261 17083 2295
rect 24777 2261 24811 2295
<< metal1 >>
rect 4062 26256 4068 26308
rect 4120 26296 4126 26308
rect 6178 26296 6184 26308
rect 4120 26268 6184 26296
rect 4120 26256 4126 26268
rect 6178 26256 6184 26268
rect 6236 26256 6242 26308
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 9953 25415 10011 25421
rect 9953 25381 9965 25415
rect 9999 25412 10011 25415
rect 10870 25412 10876 25424
rect 9999 25384 10876 25412
rect 9999 25381 10011 25384
rect 9953 25375 10011 25381
rect 10870 25372 10876 25384
rect 10928 25372 10934 25424
rect 12710 25353 12716 25356
rect 12688 25347 12716 25353
rect 12688 25313 12700 25347
rect 12688 25307 12716 25313
rect 12710 25304 12716 25307
rect 12768 25304 12774 25356
rect 9674 25236 9680 25288
rect 9732 25276 9738 25288
rect 9861 25279 9919 25285
rect 9861 25276 9873 25279
rect 9732 25248 9873 25276
rect 9732 25236 9738 25248
rect 9861 25245 9873 25248
rect 9907 25245 9919 25279
rect 10134 25276 10140 25288
rect 10095 25248 10140 25276
rect 9861 25239 9919 25245
rect 10134 25236 10140 25248
rect 10192 25236 10198 25288
rect 10686 25100 10692 25152
rect 10744 25140 10750 25152
rect 10781 25143 10839 25149
rect 10781 25140 10793 25143
rect 10744 25112 10793 25140
rect 10744 25100 10750 25112
rect 10781 25109 10793 25112
rect 10827 25109 10839 25143
rect 10781 25103 10839 25109
rect 12526 25100 12532 25152
rect 12584 25140 12590 25152
rect 12759 25143 12817 25149
rect 12759 25140 12771 25143
rect 12584 25112 12771 25140
rect 12584 25100 12590 25112
rect 12759 25109 12771 25112
rect 12805 25109 12817 25143
rect 12759 25103 12817 25109
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 12710 24936 12716 24948
rect 12671 24908 12716 24936
rect 12710 24896 12716 24908
rect 12768 24896 12774 24948
rect 5534 24760 5540 24812
rect 5592 24800 5598 24812
rect 5721 24803 5779 24809
rect 5721 24800 5733 24803
rect 5592 24772 5733 24800
rect 5592 24760 5598 24772
rect 5721 24769 5733 24772
rect 5767 24769 5779 24803
rect 8570 24800 8576 24812
rect 8531 24772 8576 24800
rect 5721 24763 5779 24769
rect 8570 24760 8576 24772
rect 8628 24760 8634 24812
rect 9769 24803 9827 24809
rect 9769 24769 9781 24803
rect 9815 24800 9827 24803
rect 10134 24800 10140 24812
rect 9815 24772 10140 24800
rect 9815 24769 9827 24772
rect 9769 24763 9827 24769
rect 5328 24735 5386 24741
rect 5328 24701 5340 24735
rect 5374 24732 5386 24735
rect 5552 24732 5580 24760
rect 5374 24704 5580 24732
rect 8088 24735 8146 24741
rect 5374 24701 5386 24704
rect 5328 24695 5386 24701
rect 8088 24701 8100 24735
rect 8134 24732 8146 24735
rect 8588 24732 8616 24760
rect 9968 24744 9996 24772
rect 10134 24760 10140 24772
rect 10192 24760 10198 24812
rect 15930 24800 15936 24812
rect 15891 24772 15936 24800
rect 15930 24760 15936 24772
rect 15988 24760 15994 24812
rect 8134 24704 8616 24732
rect 8134 24701 8146 24704
rect 8088 24695 8146 24701
rect 9950 24692 9956 24744
rect 10008 24692 10014 24744
rect 13262 24732 13268 24744
rect 13223 24704 13268 24732
rect 13262 24692 13268 24704
rect 13320 24732 13326 24744
rect 13817 24735 13875 24741
rect 13817 24732 13829 24735
rect 13320 24704 13829 24732
rect 13320 24692 13326 24704
rect 13817 24701 13829 24704
rect 13863 24701 13875 24735
rect 13817 24695 13875 24701
rect 15448 24735 15506 24741
rect 15448 24701 15460 24735
rect 15494 24732 15506 24735
rect 15948 24732 15976 24760
rect 15494 24704 15976 24732
rect 15494 24701 15506 24704
rect 15448 24695 15506 24701
rect 9122 24664 9128 24676
rect 9083 24636 9128 24664
rect 9122 24624 9128 24636
rect 9180 24624 9186 24676
rect 9214 24624 9220 24676
rect 9272 24664 9278 24676
rect 9272 24636 9317 24664
rect 9272 24624 9278 24636
rect 10134 24624 10140 24676
rect 10192 24664 10198 24676
rect 10686 24664 10692 24676
rect 10192 24636 10692 24664
rect 10192 24624 10198 24636
rect 10686 24624 10692 24636
rect 10744 24624 10750 24676
rect 10781 24667 10839 24673
rect 10781 24633 10793 24667
rect 10827 24664 10839 24667
rect 10870 24664 10876 24676
rect 10827 24636 10876 24664
rect 10827 24633 10839 24636
rect 10781 24627 10839 24633
rect 5442 24605 5448 24608
rect 5399 24599 5448 24605
rect 5399 24565 5411 24599
rect 5445 24565 5448 24599
rect 5399 24559 5448 24565
rect 5442 24556 5448 24559
rect 5500 24556 5506 24608
rect 6822 24596 6828 24608
rect 6783 24568 6828 24596
rect 6822 24556 6828 24568
rect 6880 24556 6886 24608
rect 7650 24556 7656 24608
rect 7708 24596 7714 24608
rect 8159 24599 8217 24605
rect 8159 24596 8171 24599
rect 7708 24568 8171 24596
rect 7708 24556 7714 24568
rect 8159 24565 8171 24568
rect 8205 24565 8217 24599
rect 8159 24559 8217 24565
rect 8941 24599 8999 24605
rect 8941 24565 8953 24599
rect 8987 24596 8999 24599
rect 9232 24596 9260 24624
rect 8987 24568 9260 24596
rect 10045 24599 10103 24605
rect 8987 24565 8999 24568
rect 8941 24559 8999 24565
rect 10045 24565 10057 24599
rect 10091 24596 10103 24599
rect 10505 24599 10563 24605
rect 10505 24596 10517 24599
rect 10091 24568 10517 24596
rect 10091 24565 10103 24568
rect 10045 24559 10103 24565
rect 10505 24565 10517 24568
rect 10551 24596 10563 24599
rect 10796 24596 10824 24627
rect 10870 24624 10876 24636
rect 10928 24624 10934 24676
rect 11333 24667 11391 24673
rect 11333 24633 11345 24667
rect 11379 24664 11391 24667
rect 11422 24664 11428 24676
rect 11379 24636 11428 24664
rect 11379 24633 11391 24636
rect 11333 24627 11391 24633
rect 11422 24624 11428 24636
rect 11480 24624 11486 24676
rect 13446 24596 13452 24608
rect 10551 24568 10824 24596
rect 13407 24568 13452 24596
rect 10551 24565 10563 24568
rect 10505 24559 10563 24565
rect 13446 24556 13452 24568
rect 13504 24556 13510 24608
rect 15519 24599 15577 24605
rect 15519 24565 15531 24599
rect 15565 24596 15577 24599
rect 16206 24596 16212 24608
rect 15565 24568 16212 24596
rect 15565 24565 15577 24568
rect 15519 24559 15577 24565
rect 16206 24556 16212 24568
rect 16264 24556 16270 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 4479 24395 4537 24401
rect 4479 24361 4491 24395
rect 4525 24392 4537 24395
rect 9122 24392 9128 24404
rect 4525 24364 8156 24392
rect 9083 24364 9128 24392
rect 4525 24361 4537 24364
rect 4479 24355 4537 24361
rect 8128 24336 8156 24364
rect 9122 24352 9128 24364
rect 9180 24352 9186 24404
rect 18230 24392 18236 24404
rect 18191 24364 18236 24392
rect 18230 24352 18236 24364
rect 18288 24352 18294 24404
rect 6546 24324 6552 24336
rect 6507 24296 6552 24324
rect 6546 24284 6552 24296
rect 6604 24284 6610 24336
rect 8110 24324 8116 24336
rect 8023 24296 8116 24324
rect 8110 24284 8116 24296
rect 8168 24284 8174 24336
rect 8205 24327 8263 24333
rect 8205 24293 8217 24327
rect 8251 24324 8263 24327
rect 8478 24324 8484 24336
rect 8251 24296 8484 24324
rect 8251 24293 8263 24296
rect 8205 24287 8263 24293
rect 8478 24284 8484 24296
rect 8536 24284 8542 24336
rect 9214 24284 9220 24336
rect 9272 24324 9278 24336
rect 10873 24327 10931 24333
rect 10873 24324 10885 24327
rect 9272 24296 10885 24324
rect 9272 24284 9278 24296
rect 10873 24293 10885 24296
rect 10919 24324 10931 24327
rect 10962 24324 10968 24336
rect 10919 24296 10968 24324
rect 10919 24293 10931 24296
rect 10873 24287 10931 24293
rect 10962 24284 10968 24296
rect 11020 24284 11026 24336
rect 11422 24324 11428 24336
rect 11383 24296 11428 24324
rect 11422 24284 11428 24296
rect 11480 24284 11486 24336
rect 12986 24324 12992 24336
rect 12947 24296 12992 24324
rect 12986 24284 12992 24296
rect 13044 24284 13050 24336
rect 1486 24265 1492 24268
rect 1464 24259 1492 24265
rect 1464 24225 1476 24259
rect 1464 24219 1492 24225
rect 1486 24216 1492 24219
rect 1544 24216 1550 24268
rect 4408 24259 4466 24265
rect 4408 24225 4420 24259
rect 4454 24256 4466 24259
rect 4614 24256 4620 24268
rect 4454 24228 4620 24256
rect 4454 24225 4466 24228
rect 4408 24219 4466 24225
rect 4614 24216 4620 24228
rect 4672 24216 4678 24268
rect 5420 24259 5478 24265
rect 5420 24225 5432 24259
rect 5466 24256 5478 24259
rect 8757 24259 8815 24265
rect 5466 24228 5672 24256
rect 5466 24225 5478 24228
rect 5420 24219 5478 24225
rect 1535 24123 1593 24129
rect 1535 24089 1547 24123
rect 1581 24120 1593 24123
rect 2682 24120 2688 24132
rect 1581 24092 2688 24120
rect 1581 24089 1593 24092
rect 1535 24083 1593 24089
rect 2682 24080 2688 24092
rect 2740 24080 2746 24132
rect 5644 24120 5672 24228
rect 8757 24225 8769 24259
rect 8803 24256 8815 24259
rect 9950 24256 9956 24268
rect 8803 24228 9956 24256
rect 8803 24225 8815 24228
rect 8757 24219 8815 24225
rect 9950 24216 9956 24228
rect 10008 24216 10014 24268
rect 15378 24265 15384 24268
rect 15356 24259 15384 24265
rect 15356 24225 15368 24259
rect 15356 24219 15384 24225
rect 15378 24216 15384 24219
rect 15436 24216 15442 24268
rect 16298 24256 16304 24268
rect 16259 24228 16304 24256
rect 16298 24216 16304 24228
rect 16356 24216 16362 24268
rect 18049 24259 18107 24265
rect 18049 24225 18061 24259
rect 18095 24256 18107 24259
rect 18414 24256 18420 24268
rect 18095 24228 18420 24256
rect 18095 24225 18107 24228
rect 18049 24219 18107 24225
rect 18414 24216 18420 24228
rect 18472 24216 18478 24268
rect 6454 24188 6460 24200
rect 6415 24160 6460 24188
rect 6454 24148 6460 24160
rect 6512 24148 6518 24200
rect 6730 24188 6736 24200
rect 6691 24160 6736 24188
rect 6730 24148 6736 24160
rect 6788 24148 6794 24200
rect 9677 24191 9735 24197
rect 9677 24157 9689 24191
rect 9723 24188 9735 24191
rect 10781 24191 10839 24197
rect 10781 24188 10793 24191
rect 9723 24160 10793 24188
rect 9723 24157 9735 24160
rect 9677 24151 9735 24157
rect 10781 24157 10793 24160
rect 10827 24188 10839 24191
rect 11514 24188 11520 24200
rect 10827 24160 11520 24188
rect 10827 24157 10839 24160
rect 10781 24151 10839 24157
rect 11514 24148 11520 24160
rect 11572 24148 11578 24200
rect 12710 24148 12716 24200
rect 12768 24188 12774 24200
rect 12897 24191 12955 24197
rect 12897 24188 12909 24191
rect 12768 24160 12909 24188
rect 12768 24148 12774 24160
rect 12897 24157 12909 24160
rect 12943 24157 12955 24191
rect 13538 24188 13544 24200
rect 13499 24160 13544 24188
rect 12897 24151 12955 24157
rect 13538 24148 13544 24160
rect 13596 24148 13602 24200
rect 6638 24120 6644 24132
rect 5644 24092 6644 24120
rect 6638 24080 6644 24092
rect 6696 24080 6702 24132
rect 9858 24080 9864 24132
rect 9916 24120 9922 24132
rect 10137 24123 10195 24129
rect 10137 24120 10149 24123
rect 9916 24092 10149 24120
rect 9916 24080 9922 24092
rect 10137 24089 10149 24092
rect 10183 24089 10195 24123
rect 16482 24120 16488 24132
rect 16443 24092 16488 24120
rect 10137 24083 10195 24089
rect 16482 24080 16488 24092
rect 16540 24080 16546 24132
rect 5258 24052 5264 24064
rect 5219 24024 5264 24052
rect 5258 24012 5264 24024
rect 5316 24012 5322 24064
rect 5534 24061 5540 24064
rect 5491 24055 5540 24061
rect 5491 24021 5503 24055
rect 5537 24021 5540 24055
rect 5491 24015 5540 24021
rect 5534 24012 5540 24015
rect 5592 24012 5598 24064
rect 7558 24052 7564 24064
rect 7519 24024 7564 24052
rect 7558 24012 7564 24024
rect 7616 24012 7622 24064
rect 10597 24055 10655 24061
rect 10597 24021 10609 24055
rect 10643 24052 10655 24055
rect 10686 24052 10692 24064
rect 10643 24024 10692 24052
rect 10643 24021 10655 24024
rect 10597 24015 10655 24021
rect 10686 24012 10692 24024
rect 10744 24012 10750 24064
rect 14090 24052 14096 24064
rect 14051 24024 14096 24052
rect 14090 24012 14096 24024
rect 14148 24012 14154 24064
rect 15286 24012 15292 24064
rect 15344 24052 15350 24064
rect 15427 24055 15485 24061
rect 15427 24052 15439 24055
rect 15344 24024 15439 24052
rect 15344 24012 15350 24024
rect 15427 24021 15439 24024
rect 15473 24021 15485 24055
rect 15427 24015 15485 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1486 23808 1492 23860
rect 1544 23848 1550 23860
rect 2225 23851 2283 23857
rect 2225 23848 2237 23851
rect 1544 23820 2237 23848
rect 1544 23808 1550 23820
rect 2225 23817 2237 23820
rect 2271 23817 2283 23851
rect 2225 23811 2283 23817
rect 4614 23808 4620 23860
rect 4672 23848 4678 23860
rect 4985 23851 5043 23857
rect 4985 23848 4997 23851
rect 4672 23820 4997 23848
rect 4672 23808 4678 23820
rect 4985 23817 4997 23820
rect 5031 23817 5043 23851
rect 4985 23811 5043 23817
rect 6273 23851 6331 23857
rect 6273 23817 6285 23851
rect 6319 23848 6331 23851
rect 6638 23848 6644 23860
rect 6319 23820 6644 23848
rect 6319 23817 6331 23820
rect 6273 23811 6331 23817
rect 6638 23808 6644 23820
rect 6696 23808 6702 23860
rect 8110 23808 8116 23860
rect 8168 23848 8174 23860
rect 8849 23851 8907 23857
rect 8849 23848 8861 23851
rect 8168 23820 8861 23848
rect 8168 23808 8174 23820
rect 8849 23817 8861 23820
rect 8895 23817 8907 23851
rect 8849 23811 8907 23817
rect 9122 23808 9128 23860
rect 9180 23857 9186 23860
rect 9180 23851 9229 23857
rect 9180 23817 9183 23851
rect 9217 23817 9229 23851
rect 9950 23848 9956 23860
rect 9911 23820 9956 23848
rect 9180 23811 9229 23817
rect 9180 23808 9186 23811
rect 9950 23808 9956 23820
rect 10008 23848 10014 23860
rect 11514 23848 11520 23860
rect 10008 23820 10640 23848
rect 11475 23820 11520 23848
rect 10008 23808 10014 23820
rect 6546 23780 6552 23792
rect 6507 23752 6552 23780
rect 6546 23740 6552 23752
rect 6604 23740 6610 23792
rect 8478 23780 8484 23792
rect 8439 23752 8484 23780
rect 8478 23740 8484 23752
rect 8536 23740 8542 23792
rect 1535 23715 1593 23721
rect 1535 23681 1547 23715
rect 1581 23712 1593 23715
rect 5258 23712 5264 23724
rect 1581 23684 5264 23712
rect 1581 23681 1593 23684
rect 1535 23675 1593 23681
rect 5258 23672 5264 23684
rect 5316 23672 5322 23724
rect 7834 23712 7840 23724
rect 7795 23684 7840 23712
rect 7834 23672 7840 23684
rect 7892 23672 7898 23724
rect 10612 23721 10640 23820
rect 11514 23808 11520 23820
rect 11572 23808 11578 23860
rect 12158 23848 12164 23860
rect 12119 23820 12164 23848
rect 12158 23808 12164 23820
rect 12216 23808 12222 23860
rect 15930 23848 15936 23860
rect 15891 23820 15936 23848
rect 15930 23808 15936 23820
rect 15988 23808 15994 23860
rect 16298 23808 16304 23860
rect 16356 23848 16362 23860
rect 16482 23848 16488 23860
rect 16356 23820 16488 23848
rect 16356 23808 16362 23820
rect 16482 23808 16488 23820
rect 16540 23848 16546 23860
rect 16669 23851 16727 23857
rect 16669 23848 16681 23851
rect 16540 23820 16681 23848
rect 16540 23808 16546 23820
rect 16669 23817 16681 23820
rect 16715 23817 16727 23851
rect 16669 23811 16727 23817
rect 17037 23851 17095 23857
rect 17037 23817 17049 23851
rect 17083 23848 17095 23851
rect 17126 23848 17132 23860
rect 17083 23820 17132 23848
rect 17083 23817 17095 23820
rect 17037 23811 17095 23817
rect 17126 23808 17132 23820
rect 17184 23808 17190 23860
rect 19242 23848 19248 23860
rect 19203 23820 19248 23848
rect 19242 23808 19248 23820
rect 19300 23808 19306 23860
rect 21266 23848 21272 23860
rect 21227 23820 21272 23848
rect 21266 23808 21272 23820
rect 21324 23808 21330 23860
rect 22370 23848 22376 23860
rect 22331 23820 22376 23848
rect 22370 23808 22376 23820
rect 22428 23808 22434 23860
rect 11238 23740 11244 23792
rect 11296 23780 11302 23792
rect 11296 23752 12848 23780
rect 11296 23740 11302 23752
rect 10597 23715 10655 23721
rect 10597 23681 10609 23715
rect 10643 23681 10655 23715
rect 12526 23712 12532 23724
rect 12487 23684 12532 23712
rect 10597 23675 10655 23681
rect 12526 23672 12532 23684
rect 12584 23672 12590 23724
rect 12820 23721 12848 23752
rect 12805 23715 12863 23721
rect 12805 23681 12817 23715
rect 12851 23681 12863 23715
rect 12805 23675 12863 23681
rect 13538 23672 13544 23724
rect 13596 23712 13602 23724
rect 14182 23712 14188 23724
rect 13596 23684 14188 23712
rect 13596 23672 13602 23684
rect 14182 23672 14188 23684
rect 14240 23712 14246 23724
rect 14369 23715 14427 23721
rect 14369 23712 14381 23715
rect 14240 23684 14381 23712
rect 14240 23672 14246 23684
rect 14369 23681 14381 23684
rect 14415 23681 14427 23715
rect 14369 23675 14427 23681
rect 17126 23672 17132 23724
rect 17184 23712 17190 23724
rect 17184 23684 19104 23712
rect 17184 23672 17190 23684
rect 474 23604 480 23656
rect 532 23644 538 23656
rect 2498 23653 2504 23656
rect 1432 23647 1490 23653
rect 1432 23644 1444 23647
rect 532 23616 1444 23644
rect 532 23604 538 23616
rect 1432 23613 1444 23616
rect 1478 23644 1490 23647
rect 1857 23647 1915 23653
rect 1857 23644 1869 23647
rect 1478 23616 1869 23644
rect 1478 23613 1490 23616
rect 1432 23607 1490 23613
rect 1857 23613 1869 23616
rect 1903 23613 1915 23647
rect 1857 23607 1915 23613
rect 2476 23647 2504 23653
rect 2476 23613 2488 23647
rect 2556 23644 2562 23656
rect 2869 23647 2927 23653
rect 2869 23644 2881 23647
rect 2556 23616 2881 23644
rect 2476 23607 2504 23613
rect 2498 23604 2504 23607
rect 2556 23604 2562 23616
rect 2869 23613 2881 23616
rect 2915 23613 2927 23647
rect 2869 23607 2927 23613
rect 3510 23604 3516 23656
rect 3568 23644 3574 23656
rect 4192 23647 4250 23653
rect 4192 23644 4204 23647
rect 3568 23616 4204 23644
rect 3568 23604 3574 23616
rect 4192 23613 4204 23616
rect 4238 23644 4250 23647
rect 4617 23647 4675 23653
rect 4617 23644 4629 23647
rect 4238 23616 4629 23644
rect 4238 23613 4250 23616
rect 4192 23607 4250 23613
rect 4617 23613 4629 23616
rect 4663 23613 4675 23647
rect 9068 23647 9126 23653
rect 9068 23644 9080 23647
rect 4617 23607 4675 23613
rect 8772 23616 9080 23644
rect 5350 23576 5356 23588
rect 5311 23548 5356 23576
rect 5350 23536 5356 23548
rect 5408 23536 5414 23588
rect 5902 23576 5908 23588
rect 5863 23548 5908 23576
rect 5902 23536 5908 23548
rect 5960 23536 5966 23588
rect 7558 23576 7564 23588
rect 7519 23548 7564 23576
rect 7558 23536 7564 23548
rect 7616 23536 7622 23588
rect 7653 23579 7711 23585
rect 7653 23545 7665 23579
rect 7699 23545 7711 23579
rect 7653 23539 7711 23545
rect 2547 23511 2605 23517
rect 2547 23477 2559 23511
rect 2593 23508 2605 23511
rect 2682 23508 2688 23520
rect 2593 23480 2688 23508
rect 2593 23477 2605 23480
rect 2547 23471 2605 23477
rect 2682 23468 2688 23480
rect 2740 23468 2746 23520
rect 4295 23511 4353 23517
rect 4295 23477 4307 23511
rect 4341 23508 4353 23511
rect 6454 23508 6460 23520
rect 4341 23480 6460 23508
rect 4341 23477 4353 23480
rect 4295 23471 4353 23477
rect 6454 23468 6460 23480
rect 6512 23468 6518 23520
rect 7098 23468 7104 23520
rect 7156 23508 7162 23520
rect 7285 23511 7343 23517
rect 7285 23508 7297 23511
rect 7156 23480 7297 23508
rect 7156 23468 7162 23480
rect 7285 23477 7297 23480
rect 7331 23508 7343 23511
rect 7668 23508 7696 23539
rect 7742 23536 7748 23588
rect 7800 23576 7806 23588
rect 8772 23576 8800 23616
rect 9068 23613 9080 23616
rect 9114 23644 9126 23647
rect 9493 23647 9551 23653
rect 9493 23644 9505 23647
rect 9114 23616 9505 23644
rect 9114 23613 9126 23616
rect 9068 23607 9126 23613
rect 9493 23613 9505 23616
rect 9539 23613 9551 23647
rect 15378 23644 15384 23656
rect 15339 23616 15384 23644
rect 9493 23607 9551 23613
rect 15378 23604 15384 23616
rect 15436 23604 15442 23656
rect 15749 23647 15807 23653
rect 15749 23613 15761 23647
rect 15795 23644 15807 23647
rect 16850 23644 16856 23656
rect 15795 23616 16436 23644
rect 16811 23616 16856 23644
rect 15795 23613 15807 23616
rect 15749 23607 15807 23613
rect 7800 23548 8800 23576
rect 7800 23536 7806 23548
rect 10686 23536 10692 23588
rect 10744 23576 10750 23588
rect 11241 23579 11299 23585
rect 10744 23548 10789 23576
rect 10744 23536 10750 23548
rect 11241 23545 11253 23579
rect 11287 23576 11299 23579
rect 11422 23576 11428 23588
rect 11287 23548 11428 23576
rect 11287 23545 11299 23548
rect 11241 23539 11299 23545
rect 11422 23536 11428 23548
rect 11480 23536 11486 23588
rect 12158 23536 12164 23588
rect 12216 23576 12222 23588
rect 12621 23579 12679 23585
rect 12621 23576 12633 23579
rect 12216 23548 12633 23576
rect 12216 23536 12222 23548
rect 12621 23545 12633 23548
rect 12667 23545 12679 23579
rect 14090 23576 14096 23588
rect 14051 23548 14096 23576
rect 12621 23539 12679 23545
rect 14090 23536 14096 23548
rect 14148 23536 14154 23588
rect 14185 23579 14243 23585
rect 14185 23545 14197 23579
rect 14231 23576 14243 23579
rect 15102 23576 15108 23588
rect 14231 23548 15108 23576
rect 14231 23545 14243 23548
rect 14185 23539 14243 23545
rect 7331 23480 7696 23508
rect 10413 23511 10471 23517
rect 7331 23477 7343 23480
rect 7285 23471 7343 23477
rect 10413 23477 10425 23511
rect 10459 23508 10471 23511
rect 10962 23508 10968 23520
rect 10459 23480 10968 23508
rect 10459 23477 10471 23480
rect 10413 23471 10471 23477
rect 10962 23468 10968 23480
rect 11020 23468 11026 23520
rect 12986 23468 12992 23520
rect 13044 23508 13050 23520
rect 13449 23511 13507 23517
rect 13449 23508 13461 23511
rect 13044 23480 13461 23508
rect 13044 23468 13050 23480
rect 13449 23477 13461 23480
rect 13495 23477 13507 23511
rect 13449 23471 13507 23477
rect 13909 23511 13967 23517
rect 13909 23477 13921 23511
rect 13955 23508 13967 23511
rect 14200 23508 14228 23539
rect 15102 23536 15108 23548
rect 15160 23536 15166 23588
rect 16408 23520 16436 23616
rect 16850 23604 16856 23616
rect 16908 23644 16914 23656
rect 17405 23647 17463 23653
rect 17405 23644 17417 23647
rect 16908 23616 17417 23644
rect 16908 23604 16914 23616
rect 17405 23613 17417 23616
rect 17451 23613 17463 23647
rect 17405 23607 17463 23613
rect 18046 23604 18052 23656
rect 18104 23653 18110 23656
rect 18104 23647 18142 23653
rect 18130 23613 18142 23647
rect 18104 23607 18142 23613
rect 18187 23647 18245 23653
rect 18187 23613 18199 23647
rect 18233 23644 18245 23647
rect 18506 23644 18512 23656
rect 18233 23616 18512 23644
rect 18233 23613 18245 23616
rect 18187 23607 18245 23613
rect 18104 23604 18110 23607
rect 18506 23604 18512 23616
rect 18564 23604 18570 23656
rect 19076 23653 19104 23684
rect 19426 23672 19432 23724
rect 19484 23712 19490 23724
rect 19484 23684 21128 23712
rect 19484 23672 19490 23684
rect 21100 23653 21128 23684
rect 19061 23647 19119 23653
rect 19061 23613 19073 23647
rect 19107 23644 19119 23647
rect 19613 23647 19671 23653
rect 19613 23644 19625 23647
rect 19107 23616 19625 23644
rect 19107 23613 19119 23616
rect 19061 23607 19119 23613
rect 19613 23613 19625 23616
rect 19659 23613 19671 23647
rect 19613 23607 19671 23613
rect 21085 23647 21143 23653
rect 21085 23613 21097 23647
rect 21131 23644 21143 23647
rect 22186 23644 22192 23656
rect 21131 23616 21680 23644
rect 22147 23616 22192 23644
rect 21131 23613 21143 23616
rect 21085 23607 21143 23613
rect 18064 23576 18092 23604
rect 18877 23579 18935 23585
rect 18877 23576 18889 23579
rect 18064 23548 18889 23576
rect 18877 23545 18889 23548
rect 18923 23545 18935 23579
rect 18877 23539 18935 23545
rect 21652 23520 21680 23616
rect 22186 23604 22192 23616
rect 22244 23644 22250 23656
rect 22741 23647 22799 23653
rect 22741 23644 22753 23647
rect 22244 23616 22753 23644
rect 22244 23604 22250 23616
rect 22741 23613 22753 23616
rect 22787 23613 22799 23647
rect 22741 23607 22799 23613
rect 16390 23508 16396 23520
rect 13955 23480 14228 23508
rect 16351 23480 16396 23508
rect 13955 23477 13967 23480
rect 13909 23471 13967 23477
rect 16390 23468 16396 23480
rect 16448 23468 16454 23520
rect 18414 23468 18420 23520
rect 18472 23508 18478 23520
rect 18509 23511 18567 23517
rect 18509 23508 18521 23511
rect 18472 23480 18521 23508
rect 18472 23468 18478 23480
rect 18509 23477 18521 23480
rect 18555 23477 18567 23511
rect 21634 23508 21640 23520
rect 21595 23480 21640 23508
rect 18509 23471 18567 23477
rect 21634 23468 21640 23480
rect 21692 23468 21698 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 5261 23307 5319 23313
rect 5261 23273 5273 23307
rect 5307 23304 5319 23307
rect 5350 23304 5356 23316
rect 5307 23276 5356 23304
rect 5307 23273 5319 23276
rect 5261 23267 5319 23273
rect 5350 23264 5356 23276
rect 5408 23264 5414 23316
rect 5534 23264 5540 23316
rect 5592 23264 5598 23316
rect 6454 23264 6460 23316
rect 6512 23304 6518 23316
rect 6549 23307 6607 23313
rect 6549 23304 6561 23307
rect 6512 23276 6561 23304
rect 6512 23264 6518 23276
rect 6549 23273 6561 23276
rect 6595 23273 6607 23307
rect 6549 23267 6607 23273
rect 10134 23264 10140 23316
rect 10192 23304 10198 23316
rect 10275 23307 10333 23313
rect 10275 23304 10287 23307
rect 10192 23276 10287 23304
rect 10192 23264 10198 23276
rect 10275 23273 10287 23276
rect 10321 23273 10333 23307
rect 12526 23304 12532 23316
rect 12487 23276 12532 23304
rect 10275 23267 10333 23273
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 12710 23264 12716 23316
rect 12768 23304 12774 23316
rect 12805 23307 12863 23313
rect 12805 23304 12817 23307
rect 12768 23276 12817 23304
rect 12768 23264 12774 23276
rect 12805 23273 12817 23276
rect 12851 23273 12863 23307
rect 12805 23267 12863 23273
rect 16390 23264 16396 23316
rect 16448 23313 16454 23316
rect 16448 23307 16497 23313
rect 16448 23273 16451 23307
rect 16485 23273 16497 23307
rect 16448 23267 16497 23273
rect 16448 23264 16454 23267
rect 5552 23236 5580 23264
rect 5629 23239 5687 23245
rect 5629 23236 5641 23239
rect 5552 23208 5641 23236
rect 5629 23205 5641 23208
rect 5675 23205 5687 23239
rect 5629 23199 5687 23205
rect 5721 23239 5779 23245
rect 5721 23205 5733 23239
rect 5767 23236 5779 23239
rect 5994 23236 6000 23248
rect 5767 23208 6000 23236
rect 5767 23205 5779 23208
rect 5721 23199 5779 23205
rect 5994 23196 6000 23208
rect 6052 23196 6058 23248
rect 7282 23196 7288 23248
rect 7340 23236 7346 23248
rect 7834 23236 7840 23248
rect 7340 23208 7385 23236
rect 7795 23208 7840 23236
rect 7340 23196 7346 23208
rect 7834 23196 7840 23208
rect 7892 23196 7898 23248
rect 11330 23236 11336 23248
rect 11291 23208 11336 23236
rect 11330 23196 11336 23208
rect 11388 23196 11394 23248
rect 13814 23236 13820 23248
rect 13775 23208 13820 23236
rect 13814 23196 13820 23208
rect 13872 23196 13878 23248
rect 10204 23171 10262 23177
rect 10204 23137 10216 23171
rect 10250 23168 10262 23171
rect 10962 23168 10968 23180
rect 10250 23140 10968 23168
rect 10250 23137 10262 23140
rect 10204 23131 10262 23137
rect 10962 23128 10968 23140
rect 11020 23128 11026 23180
rect 15286 23128 15292 23180
rect 15344 23177 15350 23180
rect 15344 23171 15382 23177
rect 15370 23137 15382 23171
rect 15344 23131 15382 23137
rect 15344 23128 15350 23131
rect 16298 23128 16304 23180
rect 16356 23177 16362 23180
rect 16356 23171 16394 23177
rect 16382 23137 16394 23171
rect 16356 23131 16394 23137
rect 16356 23128 16362 23131
rect 17034 23128 17040 23180
rect 17092 23168 17098 23180
rect 17348 23171 17406 23177
rect 17348 23168 17360 23171
rect 17092 23140 17360 23168
rect 17092 23128 17098 23140
rect 17348 23137 17360 23140
rect 17394 23137 17406 23171
rect 17348 23131 17406 23137
rect 5902 23060 5908 23112
rect 5960 23100 5966 23112
rect 6273 23103 6331 23109
rect 6273 23100 6285 23103
rect 5960 23072 6285 23100
rect 5960 23060 5966 23072
rect 6273 23069 6285 23072
rect 6319 23100 6331 23103
rect 6822 23100 6828 23112
rect 6319 23072 6828 23100
rect 6319 23069 6331 23072
rect 6273 23063 6331 23069
rect 6822 23060 6828 23072
rect 6880 23060 6886 23112
rect 6914 23060 6920 23112
rect 6972 23100 6978 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 6972 23072 7205 23100
rect 6972 23060 6978 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 11238 23100 11244 23112
rect 11199 23072 11244 23100
rect 7193 23063 7251 23069
rect 11238 23060 11244 23072
rect 11296 23060 11302 23112
rect 11422 23060 11428 23112
rect 11480 23100 11486 23112
rect 11517 23103 11575 23109
rect 11517 23100 11529 23103
rect 11480 23072 11529 23100
rect 11480 23060 11486 23072
rect 11517 23069 11529 23072
rect 11563 23100 11575 23103
rect 12618 23100 12624 23112
rect 11563 23072 12624 23100
rect 11563 23069 11575 23072
rect 11517 23063 11575 23069
rect 12618 23060 12624 23072
rect 12676 23060 12682 23112
rect 13722 23100 13728 23112
rect 13683 23072 13728 23100
rect 13722 23060 13728 23072
rect 13780 23060 13786 23112
rect 14182 23100 14188 23112
rect 14143 23072 14188 23100
rect 14182 23060 14188 23072
rect 14240 23060 14246 23112
rect 15378 22924 15384 22976
rect 15436 22973 15442 22976
rect 15436 22967 15485 22973
rect 15436 22933 15439 22967
rect 15473 22933 15485 22967
rect 15436 22927 15485 22933
rect 17451 22967 17509 22973
rect 17451 22933 17463 22967
rect 17497 22964 17509 22967
rect 17862 22964 17868 22976
rect 17497 22936 17868 22964
rect 17497 22933 17509 22936
rect 17451 22927 17509 22933
rect 15436 22924 15442 22927
rect 17862 22924 17868 22936
rect 17920 22924 17926 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 5534 22720 5540 22772
rect 5592 22760 5598 22772
rect 5905 22763 5963 22769
rect 5905 22760 5917 22763
rect 5592 22732 5917 22760
rect 5592 22720 5598 22732
rect 5905 22729 5917 22732
rect 5951 22729 5963 22763
rect 5905 22723 5963 22729
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 7101 22763 7159 22769
rect 7101 22760 7113 22763
rect 6972 22732 7113 22760
rect 6972 22720 6978 22732
rect 7101 22729 7113 22732
rect 7147 22729 7159 22763
rect 7101 22723 7159 22729
rect 10597 22763 10655 22769
rect 10597 22729 10609 22763
rect 10643 22760 10655 22763
rect 10686 22760 10692 22772
rect 10643 22732 10692 22760
rect 10643 22729 10655 22732
rect 10597 22723 10655 22729
rect 10686 22720 10692 22732
rect 10744 22720 10750 22772
rect 11330 22760 11336 22772
rect 11291 22732 11336 22760
rect 11330 22720 11336 22732
rect 11388 22720 11394 22772
rect 12575 22763 12633 22769
rect 12575 22729 12587 22763
rect 12621 22760 12633 22763
rect 13262 22760 13268 22772
rect 12621 22732 13268 22760
rect 12621 22729 12633 22732
rect 12575 22723 12633 22729
rect 13262 22720 13268 22732
rect 13320 22720 13326 22772
rect 13357 22763 13415 22769
rect 13357 22729 13369 22763
rect 13403 22760 13415 22763
rect 13722 22760 13728 22772
rect 13403 22732 13728 22760
rect 13403 22729 13415 22732
rect 13357 22723 13415 22729
rect 13722 22720 13728 22732
rect 13780 22720 13786 22772
rect 16482 22720 16488 22772
rect 16540 22769 16546 22772
rect 16540 22763 16589 22769
rect 16540 22729 16543 22763
rect 16577 22729 16589 22763
rect 16540 22723 16589 22729
rect 16540 22720 16546 22723
rect 17034 22720 17040 22772
rect 17092 22760 17098 22772
rect 17313 22763 17371 22769
rect 17313 22760 17325 22763
rect 17092 22732 17325 22760
rect 17092 22720 17098 22732
rect 17313 22729 17325 22732
rect 17359 22729 17371 22763
rect 17313 22723 17371 22729
rect 11238 22652 11244 22704
rect 11296 22692 11302 22704
rect 11609 22695 11667 22701
rect 11609 22692 11621 22695
rect 11296 22664 11621 22692
rect 11296 22652 11302 22664
rect 11609 22661 11621 22664
rect 11655 22661 11667 22695
rect 11609 22655 11667 22661
rect 7650 22624 7656 22636
rect 7611 22596 7656 22624
rect 7650 22584 7656 22596
rect 7708 22584 7714 22636
rect 7834 22584 7840 22636
rect 7892 22624 7898 22636
rect 7929 22627 7987 22633
rect 7929 22624 7941 22627
rect 7892 22596 7941 22624
rect 7892 22584 7898 22596
rect 7929 22593 7941 22596
rect 7975 22593 7987 22627
rect 7929 22587 7987 22593
rect 13909 22627 13967 22633
rect 13909 22593 13921 22627
rect 13955 22624 13967 22627
rect 14182 22624 14188 22636
rect 13955 22596 14188 22624
rect 13955 22593 13967 22596
rect 13909 22587 13967 22593
rect 14182 22584 14188 22596
rect 14240 22584 14246 22636
rect 15286 22624 15292 22636
rect 15199 22596 15292 22624
rect 15286 22584 15292 22596
rect 15344 22624 15350 22636
rect 17218 22624 17224 22636
rect 15344 22596 17224 22624
rect 15344 22584 15350 22596
rect 17218 22584 17224 22596
rect 17276 22584 17282 22636
rect 9677 22559 9735 22565
rect 9677 22556 9689 22559
rect 9140 22528 9689 22556
rect 6546 22448 6552 22500
rect 6604 22488 6610 22500
rect 7466 22488 7472 22500
rect 6604 22460 7472 22488
rect 6604 22448 6610 22460
rect 7466 22448 7472 22460
rect 7524 22488 7530 22500
rect 7745 22491 7803 22497
rect 7745 22488 7757 22491
rect 7524 22460 7757 22488
rect 7524 22448 7530 22460
rect 7745 22457 7757 22460
rect 7791 22457 7803 22491
rect 7745 22451 7803 22457
rect 9140 22432 9168 22528
rect 9677 22525 9689 22528
rect 9723 22525 9735 22559
rect 10962 22556 10968 22568
rect 10923 22528 10968 22556
rect 9677 22519 9735 22525
rect 10962 22516 10968 22528
rect 11020 22516 11026 22568
rect 12504 22559 12562 22565
rect 12504 22525 12516 22559
rect 12550 22556 12562 22559
rect 12618 22556 12624 22568
rect 12550 22528 12624 22556
rect 12550 22525 12562 22528
rect 12504 22519 12562 22525
rect 12618 22516 12624 22528
rect 12676 22556 12682 22568
rect 12897 22559 12955 22565
rect 12897 22556 12909 22559
rect 12676 22528 12909 22556
rect 12676 22516 12682 22528
rect 12897 22525 12909 22528
rect 12943 22525 12955 22559
rect 12897 22519 12955 22525
rect 15448 22559 15506 22565
rect 15448 22525 15460 22559
rect 15494 22556 15506 22559
rect 15657 22559 15715 22565
rect 15657 22556 15669 22559
rect 15494 22528 15669 22556
rect 15494 22525 15506 22528
rect 15448 22519 15506 22525
rect 15657 22525 15669 22528
rect 15703 22525 15715 22559
rect 16428 22559 16486 22565
rect 16428 22556 16440 22559
rect 15657 22519 15715 22525
rect 16224 22528 16440 22556
rect 9585 22491 9643 22497
rect 9585 22457 9597 22491
rect 9631 22488 9643 22491
rect 9950 22488 9956 22500
rect 9631 22460 9956 22488
rect 9631 22457 9643 22460
rect 9585 22451 9643 22457
rect 9950 22448 9956 22460
rect 10008 22497 10014 22500
rect 10008 22491 10056 22497
rect 10008 22457 10010 22491
rect 10044 22457 10056 22491
rect 10008 22451 10056 22457
rect 10008 22448 10014 22451
rect 13998 22448 14004 22500
rect 14056 22488 14062 22500
rect 14553 22491 14611 22497
rect 14056 22460 14101 22488
rect 14056 22448 14062 22460
rect 14553 22457 14565 22491
rect 14599 22488 14611 22491
rect 14734 22488 14740 22500
rect 14599 22460 14740 22488
rect 14599 22457 14611 22460
rect 14553 22451 14611 22457
rect 14734 22448 14740 22460
rect 14792 22488 14798 22500
rect 16224 22497 16252 22528
rect 16428 22525 16440 22528
rect 16474 22525 16486 22559
rect 16428 22519 16486 22525
rect 16209 22491 16267 22497
rect 16209 22488 16221 22491
rect 14792 22460 16221 22488
rect 14792 22448 14798 22460
rect 16209 22457 16221 22460
rect 16255 22457 16267 22491
rect 16209 22451 16267 22457
rect 16298 22448 16304 22500
rect 16356 22488 16362 22500
rect 16853 22491 16911 22497
rect 16853 22488 16865 22491
rect 16356 22460 16865 22488
rect 16356 22448 16362 22460
rect 16853 22457 16865 22460
rect 16899 22457 16911 22491
rect 16853 22451 16911 22457
rect 5629 22423 5687 22429
rect 5629 22389 5641 22423
rect 5675 22420 5687 22423
rect 5994 22420 6000 22432
rect 5675 22392 6000 22420
rect 5675 22389 5687 22392
rect 5629 22383 5687 22389
rect 5994 22380 6000 22392
rect 6052 22420 6058 22432
rect 6641 22423 6699 22429
rect 6641 22420 6653 22423
rect 6052 22392 6653 22420
rect 6052 22380 6058 22392
rect 6641 22389 6653 22392
rect 6687 22420 6699 22423
rect 7282 22420 7288 22432
rect 6687 22392 7288 22420
rect 6687 22389 6699 22392
rect 6641 22383 6699 22389
rect 7282 22380 7288 22392
rect 7340 22380 7346 22432
rect 9122 22420 9128 22432
rect 9083 22392 9128 22420
rect 9122 22380 9128 22392
rect 9180 22380 9186 22432
rect 13725 22423 13783 22429
rect 13725 22389 13737 22423
rect 13771 22420 13783 22423
rect 13814 22420 13820 22432
rect 13771 22392 13820 22420
rect 13771 22389 13783 22392
rect 13725 22383 13783 22389
rect 13814 22380 13820 22392
rect 13872 22420 13878 22432
rect 14642 22420 14648 22432
rect 13872 22392 14648 22420
rect 13872 22380 13878 22392
rect 14642 22380 14648 22392
rect 14700 22380 14706 22432
rect 15378 22380 15384 22432
rect 15436 22420 15442 22432
rect 15519 22423 15577 22429
rect 15519 22420 15531 22423
rect 15436 22392 15531 22420
rect 15436 22380 15442 22392
rect 15519 22389 15531 22392
rect 15565 22389 15577 22423
rect 15519 22383 15577 22389
rect 15657 22423 15715 22429
rect 15657 22389 15669 22423
rect 15703 22420 15715 22423
rect 15933 22423 15991 22429
rect 15933 22420 15945 22423
rect 15703 22392 15945 22420
rect 15703 22389 15715 22392
rect 15657 22383 15715 22389
rect 15933 22389 15945 22392
rect 15979 22420 15991 22423
rect 17126 22420 17132 22432
rect 15979 22392 17132 22420
rect 15979 22389 15991 22392
rect 15933 22383 15991 22389
rect 17126 22380 17132 22392
rect 17184 22380 17190 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 5074 22216 5080 22228
rect 5035 22188 5080 22216
rect 5074 22176 5080 22188
rect 5132 22176 5138 22228
rect 7466 22176 7472 22228
rect 7524 22216 7530 22228
rect 7561 22219 7619 22225
rect 7561 22216 7573 22219
rect 7524 22188 7573 22216
rect 7524 22176 7530 22188
rect 7561 22185 7573 22188
rect 7607 22185 7619 22219
rect 7561 22179 7619 22185
rect 7834 22176 7840 22228
rect 7892 22216 7898 22228
rect 11241 22219 11299 22225
rect 7892 22188 8248 22216
rect 7892 22176 7898 22188
rect 6178 22108 6184 22160
rect 6236 22148 6242 22160
rect 6686 22151 6744 22157
rect 6686 22148 6698 22151
rect 6236 22120 6698 22148
rect 6236 22108 6242 22120
rect 6686 22117 6698 22120
rect 6732 22117 6744 22151
rect 6686 22111 6744 22117
rect 7650 22108 7656 22160
rect 7708 22148 7714 22160
rect 7929 22151 7987 22157
rect 7929 22148 7941 22151
rect 7708 22120 7941 22148
rect 7708 22108 7714 22120
rect 7929 22117 7941 22120
rect 7975 22117 7987 22151
rect 8220 22148 8248 22188
rect 11241 22185 11253 22219
rect 11287 22216 11299 22219
rect 11330 22216 11336 22228
rect 11287 22188 11336 22216
rect 11287 22185 11299 22188
rect 11241 22179 11299 22185
rect 11330 22176 11336 22188
rect 11388 22176 11394 22228
rect 13909 22219 13967 22225
rect 13909 22185 13921 22219
rect 13955 22216 13967 22219
rect 13998 22216 14004 22228
rect 13955 22188 14004 22216
rect 13955 22185 13967 22188
rect 13909 22179 13967 22185
rect 8220 22120 8340 22148
rect 7929 22111 7987 22117
rect 5074 22080 5080 22092
rect 5035 22052 5080 22080
rect 5074 22040 5080 22052
rect 5132 22040 5138 22092
rect 5353 22083 5411 22089
rect 5353 22049 5365 22083
rect 5399 22080 5411 22083
rect 5442 22080 5448 22092
rect 5399 22052 5448 22080
rect 5399 22049 5411 22052
rect 5353 22043 5411 22049
rect 5442 22040 5448 22052
rect 5500 22040 5506 22092
rect 8110 22040 8116 22092
rect 8168 22089 8174 22092
rect 8168 22083 8206 22089
rect 8194 22049 8206 22083
rect 8312 22080 8340 22120
rect 9950 22108 9956 22160
rect 10008 22148 10014 22160
rect 10642 22151 10700 22157
rect 10642 22148 10654 22151
rect 10008 22120 10654 22148
rect 10008 22108 10014 22120
rect 10642 22117 10654 22120
rect 10688 22117 10700 22151
rect 12850 22151 12908 22157
rect 12850 22148 12862 22151
rect 10642 22111 10700 22117
rect 12452 22120 12862 22148
rect 8573 22083 8631 22089
rect 8573 22080 8585 22083
rect 8312 22052 8585 22080
rect 8168 22043 8206 22049
rect 8573 22049 8585 22052
rect 8619 22080 8631 22083
rect 8662 22080 8668 22092
rect 8619 22052 8668 22080
rect 8619 22049 8631 22052
rect 8573 22043 8631 22049
rect 8168 22040 8174 22043
rect 8662 22040 8668 22052
rect 8720 22040 8726 22092
rect 12250 22040 12256 22092
rect 12308 22080 12314 22092
rect 12452 22080 12480 22120
rect 12850 22117 12862 22120
rect 12896 22117 12908 22151
rect 12850 22111 12908 22117
rect 12308 22052 12480 22080
rect 13449 22083 13507 22089
rect 12308 22040 12314 22052
rect 13449 22049 13461 22083
rect 13495 22080 13507 22083
rect 13924 22080 13952 22179
rect 13998 22176 14004 22188
rect 14056 22176 14062 22228
rect 14182 22216 14188 22228
rect 14143 22188 14188 22216
rect 14182 22176 14188 22188
rect 14240 22176 14246 22228
rect 15381 22219 15439 22225
rect 15381 22216 15393 22219
rect 15166 22188 15393 22216
rect 15166 22080 15194 22188
rect 15381 22185 15393 22188
rect 15427 22185 15439 22219
rect 15381 22179 15439 22185
rect 17218 22148 17224 22160
rect 16868 22120 17224 22148
rect 15562 22080 15568 22092
rect 13495 22052 13952 22080
rect 14016 22052 15194 22080
rect 15523 22052 15568 22080
rect 13495 22049 13507 22052
rect 13449 22043 13507 22049
rect 6362 22012 6368 22024
rect 6323 21984 6368 22012
rect 6362 21972 6368 21984
rect 6420 21972 6426 22024
rect 7558 21972 7564 22024
rect 7616 22012 7622 22024
rect 8251 22015 8309 22021
rect 8251 22012 8263 22015
rect 7616 21984 8263 22012
rect 7616 21972 7622 21984
rect 8251 21981 8263 21984
rect 8297 21981 8309 22015
rect 8251 21975 8309 21981
rect 10134 21972 10140 22024
rect 10192 22012 10198 22024
rect 10321 22015 10379 22021
rect 10321 22012 10333 22015
rect 10192 21984 10333 22012
rect 10192 21972 10198 21984
rect 10321 21981 10333 21984
rect 10367 21981 10379 22015
rect 10321 21975 10379 21981
rect 11882 21972 11888 22024
rect 11940 22012 11946 22024
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 11940 21984 12541 22012
rect 11940 21972 11946 21984
rect 12529 21981 12541 21984
rect 12575 22012 12587 22015
rect 14016 22012 14044 22052
rect 15562 22040 15568 22052
rect 15620 22040 15626 22092
rect 15746 22080 15752 22092
rect 15707 22052 15752 22080
rect 15746 22040 15752 22052
rect 15804 22040 15810 22092
rect 16868 22089 16896 22120
rect 17218 22108 17224 22120
rect 17276 22108 17282 22160
rect 16859 22083 16917 22089
rect 16859 22049 16871 22083
rect 16905 22049 16917 22083
rect 16859 22043 16917 22049
rect 12575 21984 14044 22012
rect 12575 21981 12587 21984
rect 12529 21975 12587 21981
rect 17034 21944 17040 21956
rect 16995 21916 17040 21944
rect 17034 21904 17040 21916
rect 17092 21904 17098 21956
rect 5905 21879 5963 21885
rect 5905 21845 5917 21879
rect 5951 21876 5963 21879
rect 5994 21876 6000 21888
rect 5951 21848 6000 21876
rect 5951 21845 5963 21848
rect 5905 21839 5963 21845
rect 5994 21836 6000 21848
rect 6052 21836 6058 21888
rect 7282 21876 7288 21888
rect 7243 21848 7288 21876
rect 7282 21836 7288 21848
rect 7340 21836 7346 21888
rect 14274 21836 14280 21888
rect 14332 21876 14338 21888
rect 14553 21879 14611 21885
rect 14553 21876 14565 21879
rect 14332 21848 14565 21876
rect 14332 21836 14338 21848
rect 14553 21845 14565 21848
rect 14599 21845 14611 21879
rect 14553 21839 14611 21845
rect 14642 21836 14648 21888
rect 14700 21876 14706 21888
rect 16298 21876 16304 21888
rect 14700 21848 16304 21876
rect 14700 21836 14706 21848
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 6178 21672 6184 21684
rect 6139 21644 6184 21672
rect 6178 21632 6184 21644
rect 6236 21672 6242 21684
rect 6549 21675 6607 21681
rect 6549 21672 6561 21675
rect 6236 21644 6561 21672
rect 6236 21632 6242 21644
rect 6549 21641 6561 21644
rect 6595 21641 6607 21675
rect 11882 21672 11888 21684
rect 11843 21644 11888 21672
rect 6549 21635 6607 21641
rect 6564 21548 6592 21635
rect 11882 21632 11888 21644
rect 11940 21632 11946 21684
rect 13722 21672 13728 21684
rect 13683 21644 13728 21672
rect 13722 21632 13728 21644
rect 13780 21632 13786 21684
rect 5994 21536 6000 21548
rect 5460 21508 6000 21536
rect 5460 21477 5488 21508
rect 5994 21496 6000 21508
rect 6052 21496 6058 21548
rect 6546 21536 6552 21548
rect 6459 21508 6552 21536
rect 6546 21496 6552 21508
rect 6604 21536 6610 21548
rect 8662 21536 8668 21548
rect 6604 21508 7236 21536
rect 8623 21508 8668 21536
rect 6604 21496 6610 21508
rect 5445 21471 5503 21477
rect 5445 21437 5457 21471
rect 5491 21437 5503 21471
rect 5626 21468 5632 21480
rect 5587 21440 5632 21468
rect 5445 21431 5503 21437
rect 5626 21428 5632 21440
rect 5684 21428 5690 21480
rect 5905 21471 5963 21477
rect 5905 21437 5917 21471
rect 5951 21468 5963 21471
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 5951 21440 6837 21468
rect 5951 21437 5963 21440
rect 5905 21431 5963 21437
rect 6825 21437 6837 21440
rect 6871 21468 6883 21471
rect 7006 21468 7012 21480
rect 6871 21440 7012 21468
rect 6871 21437 6883 21440
rect 6825 21431 6883 21437
rect 7006 21428 7012 21440
rect 7064 21428 7070 21480
rect 7208 21409 7236 21508
rect 8662 21496 8668 21508
rect 8720 21496 8726 21548
rect 9306 21536 9312 21548
rect 9267 21508 9312 21536
rect 9306 21496 9312 21508
rect 9364 21496 9370 21548
rect 12713 21539 12771 21545
rect 12713 21505 12725 21539
rect 12759 21536 12771 21539
rect 13740 21536 13768 21632
rect 14274 21564 14280 21616
rect 14332 21604 14338 21616
rect 16022 21604 16028 21616
rect 14332 21576 16028 21604
rect 14332 21564 14338 21576
rect 16022 21564 16028 21576
rect 16080 21604 16086 21616
rect 16080 21576 16160 21604
rect 16080 21564 16086 21576
rect 14734 21536 14740 21548
rect 12759 21508 13768 21536
rect 14695 21508 14740 21536
rect 12759 21505 12771 21508
rect 12713 21499 12771 21505
rect 14734 21496 14740 21508
rect 14792 21496 14798 21548
rect 16132 21545 16160 21576
rect 16117 21539 16175 21545
rect 16117 21505 16129 21539
rect 16163 21505 16175 21539
rect 16117 21499 16175 21505
rect 10686 21428 10692 21480
rect 10744 21468 10750 21480
rect 10781 21471 10839 21477
rect 10781 21468 10793 21471
rect 10744 21440 10793 21468
rect 10744 21428 10750 21440
rect 10781 21437 10793 21440
rect 10827 21437 10839 21471
rect 10781 21431 10839 21437
rect 11241 21471 11299 21477
rect 11241 21437 11253 21471
rect 11287 21468 11299 21471
rect 11287 21440 11321 21468
rect 11287 21437 11299 21440
rect 11241 21431 11299 21437
rect 7187 21403 7245 21409
rect 7187 21369 7199 21403
rect 7233 21369 7245 21403
rect 8662 21400 8668 21412
rect 7187 21363 7245 21369
rect 7760 21372 8668 21400
rect 4522 21332 4528 21344
rect 4483 21304 4528 21332
rect 4522 21292 4528 21304
rect 4580 21292 4586 21344
rect 4893 21335 4951 21341
rect 4893 21301 4905 21335
rect 4939 21332 4951 21335
rect 5074 21332 5080 21344
rect 4939 21304 5080 21332
rect 4939 21301 4951 21304
rect 4893 21295 4951 21301
rect 5074 21292 5080 21304
rect 5132 21332 5138 21344
rect 6178 21332 6184 21344
rect 5132 21304 6184 21332
rect 5132 21292 5138 21304
rect 6178 21292 6184 21304
rect 6236 21292 6242 21344
rect 7760 21341 7788 21372
rect 8662 21360 8668 21372
rect 8720 21400 8726 21412
rect 8757 21403 8815 21409
rect 8757 21400 8769 21403
rect 8720 21372 8769 21400
rect 8720 21360 8726 21372
rect 8757 21369 8769 21372
rect 8803 21369 8815 21403
rect 8757 21363 8815 21369
rect 10045 21403 10103 21409
rect 10045 21369 10057 21403
rect 10091 21400 10103 21403
rect 11256 21400 11284 21431
rect 11330 21400 11336 21412
rect 10091 21372 11336 21400
rect 10091 21369 10103 21372
rect 10045 21363 10103 21369
rect 11330 21360 11336 21372
rect 11388 21360 11394 21412
rect 11517 21403 11575 21409
rect 11517 21369 11529 21403
rect 11563 21400 11575 21403
rect 12434 21400 12440 21412
rect 11563 21372 12440 21400
rect 11563 21369 11575 21372
rect 11517 21363 11575 21369
rect 12434 21360 12440 21372
rect 12492 21360 12498 21412
rect 12805 21403 12863 21409
rect 12805 21369 12817 21403
rect 12851 21400 12863 21403
rect 12986 21400 12992 21412
rect 12851 21372 12992 21400
rect 12851 21369 12863 21372
rect 12805 21363 12863 21369
rect 12986 21360 12992 21372
rect 13044 21360 13050 21412
rect 13357 21403 13415 21409
rect 13357 21369 13369 21403
rect 13403 21400 13415 21403
rect 14274 21400 14280 21412
rect 13403 21372 14280 21400
rect 13403 21369 13415 21372
rect 13357 21363 13415 21369
rect 14274 21360 14280 21372
rect 14332 21360 14338 21412
rect 14369 21403 14427 21409
rect 14369 21369 14381 21403
rect 14415 21369 14427 21403
rect 15838 21400 15844 21412
rect 15799 21372 15844 21400
rect 14369 21363 14427 21369
rect 7745 21335 7803 21341
rect 7745 21301 7757 21335
rect 7791 21301 7803 21335
rect 8202 21332 8208 21344
rect 8163 21304 8208 21332
rect 7745 21295 7803 21301
rect 8202 21292 8208 21304
rect 8260 21292 8266 21344
rect 9950 21292 9956 21344
rect 10008 21332 10014 21344
rect 10321 21335 10379 21341
rect 10321 21332 10333 21335
rect 10008 21304 10333 21332
rect 10008 21292 10014 21304
rect 10321 21301 10333 21304
rect 10367 21301 10379 21335
rect 12250 21332 12256 21344
rect 12211 21304 12256 21332
rect 10321 21295 10379 21301
rect 12250 21292 12256 21304
rect 12308 21292 12314 21344
rect 13998 21332 14004 21344
rect 13959 21304 14004 21332
rect 13998 21292 14004 21304
rect 14056 21332 14062 21344
rect 14384 21332 14412 21363
rect 15838 21360 15844 21372
rect 15896 21360 15902 21412
rect 15933 21403 15991 21409
rect 15933 21369 15945 21403
rect 15979 21400 15991 21403
rect 16298 21400 16304 21412
rect 15979 21372 16304 21400
rect 15979 21369 15991 21372
rect 15933 21363 15991 21369
rect 16298 21360 16304 21372
rect 16356 21360 16362 21412
rect 15286 21332 15292 21344
rect 14056 21304 14412 21332
rect 15247 21304 15292 21332
rect 14056 21292 14062 21304
rect 15286 21292 15292 21304
rect 15344 21332 15350 21344
rect 15562 21332 15568 21344
rect 15344 21304 15568 21332
rect 15344 21292 15350 21304
rect 15562 21292 15568 21304
rect 15620 21292 15626 21344
rect 16945 21335 17003 21341
rect 16945 21301 16957 21335
rect 16991 21332 17003 21335
rect 17218 21332 17224 21344
rect 16991 21304 17224 21332
rect 16991 21301 17003 21304
rect 16945 21295 17003 21301
rect 17218 21292 17224 21304
rect 17276 21292 17282 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 7006 21128 7012 21140
rect 6967 21100 7012 21128
rect 7006 21088 7012 21100
rect 7064 21088 7070 21140
rect 8662 21128 8668 21140
rect 8623 21100 8668 21128
rect 8662 21088 8668 21100
rect 8720 21088 8726 21140
rect 11054 21088 11060 21140
rect 11112 21128 11118 21140
rect 12713 21131 12771 21137
rect 11112 21100 11284 21128
rect 11112 21088 11118 21100
rect 6362 21060 6368 21072
rect 6323 21032 6368 21060
rect 6362 21020 6368 21032
rect 6420 21060 6426 21072
rect 6641 21063 6699 21069
rect 6641 21060 6653 21063
rect 6420 21032 6653 21060
rect 6420 21020 6426 21032
rect 6641 21029 6653 21032
rect 6687 21029 6699 21063
rect 6641 21023 6699 21029
rect 7282 21020 7288 21072
rect 7340 21060 7346 21072
rect 7377 21063 7435 21069
rect 7377 21060 7389 21063
rect 7340 21032 7389 21060
rect 7340 21020 7346 21032
rect 7377 21029 7389 21032
rect 7423 21029 7435 21063
rect 7377 21023 7435 21029
rect 7929 21063 7987 21069
rect 7929 21029 7941 21063
rect 7975 21060 7987 21063
rect 8202 21060 8208 21072
rect 7975 21032 8208 21060
rect 7975 21029 7987 21032
rect 7929 21023 7987 21029
rect 8202 21020 8208 21032
rect 8260 21060 8266 21072
rect 9306 21060 9312 21072
rect 8260 21032 9312 21060
rect 8260 21020 8266 21032
rect 9306 21020 9312 21032
rect 9364 21020 9370 21072
rect 11256 21069 11284 21100
rect 12713 21097 12725 21131
rect 12759 21128 12771 21131
rect 12986 21128 12992 21140
rect 12759 21100 12992 21128
rect 12759 21097 12771 21100
rect 12713 21091 12771 21097
rect 12986 21088 12992 21100
rect 13044 21088 13050 21140
rect 13725 21131 13783 21137
rect 13725 21097 13737 21131
rect 13771 21128 13783 21131
rect 13998 21128 14004 21140
rect 13771 21100 14004 21128
rect 13771 21097 13783 21100
rect 13725 21091 13783 21097
rect 13998 21088 14004 21100
rect 14056 21088 14062 21140
rect 15010 21128 15016 21140
rect 14971 21100 15016 21128
rect 15010 21088 15016 21100
rect 15068 21088 15074 21140
rect 15838 21088 15844 21140
rect 15896 21128 15902 21140
rect 16301 21131 16359 21137
rect 16301 21128 16313 21131
rect 15896 21100 16313 21128
rect 15896 21088 15902 21100
rect 16301 21097 16313 21100
rect 16347 21097 16359 21131
rect 16301 21091 16359 21097
rect 11241 21063 11299 21069
rect 11241 21029 11253 21063
rect 11287 21029 11299 21063
rect 11241 21023 11299 21029
rect 12250 21020 12256 21072
rect 12308 21060 12314 21072
rect 13126 21063 13184 21069
rect 13126 21060 13138 21063
rect 12308 21032 13138 21060
rect 12308 21020 12314 21032
rect 13126 21029 13138 21032
rect 13172 21029 13184 21063
rect 15378 21060 15384 21072
rect 15339 21032 15384 21060
rect 13126 21023 13184 21029
rect 15378 21020 15384 21032
rect 15436 21020 15442 21072
rect 15470 21020 15476 21072
rect 15528 21060 15534 21072
rect 16022 21060 16028 21072
rect 15528 21032 15573 21060
rect 15983 21032 16028 21060
rect 15528 21020 15534 21032
rect 16022 21020 16028 21032
rect 16080 21020 16086 21072
rect 4893 20995 4951 21001
rect 4893 20961 4905 20995
rect 4939 20992 4951 20995
rect 5626 20992 5632 21004
rect 4939 20964 5632 20992
rect 4939 20961 4951 20964
rect 4893 20955 4951 20961
rect 5626 20952 5632 20964
rect 5684 20952 5690 21004
rect 6178 20992 6184 21004
rect 6139 20964 6184 20992
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 9744 20995 9802 21001
rect 9744 20961 9756 20995
rect 9790 20992 9802 20995
rect 10410 20992 10416 21004
rect 9790 20964 10416 20992
rect 9790 20961 9802 20964
rect 9744 20955 9802 20961
rect 10410 20952 10416 20964
rect 10468 20952 10474 21004
rect 6914 20884 6920 20936
rect 6972 20924 6978 20936
rect 7285 20927 7343 20933
rect 7285 20924 7297 20927
rect 6972 20896 7297 20924
rect 6972 20884 6978 20896
rect 7285 20893 7297 20896
rect 7331 20893 7343 20927
rect 7285 20887 7343 20893
rect 9858 20884 9864 20936
rect 9916 20924 9922 20936
rect 10686 20924 10692 20936
rect 9916 20896 10692 20924
rect 9916 20884 9922 20896
rect 10686 20884 10692 20896
rect 10744 20924 10750 20936
rect 10781 20927 10839 20933
rect 10781 20924 10793 20927
rect 10744 20896 10793 20924
rect 10744 20884 10750 20896
rect 10781 20893 10793 20896
rect 10827 20893 10839 20927
rect 11146 20924 11152 20936
rect 11107 20896 11152 20924
rect 10781 20887 10839 20893
rect 11146 20884 11152 20896
rect 11204 20884 11210 20936
rect 11606 20924 11612 20936
rect 11567 20896 11612 20924
rect 11606 20884 11612 20896
rect 11664 20884 11670 20936
rect 12802 20924 12808 20936
rect 12715 20896 12808 20924
rect 12802 20884 12808 20896
rect 12860 20924 12866 20936
rect 13722 20924 13728 20936
rect 12860 20896 13728 20924
rect 12860 20884 12866 20896
rect 13722 20884 13728 20896
rect 13780 20884 13786 20936
rect 9674 20816 9680 20868
rect 9732 20856 9738 20868
rect 10134 20856 10140 20868
rect 9732 20828 10140 20856
rect 9732 20816 9738 20828
rect 10134 20816 10140 20828
rect 10192 20856 10198 20868
rect 10321 20859 10379 20865
rect 10321 20856 10333 20859
rect 10192 20828 10333 20856
rect 10192 20816 10198 20828
rect 10321 20825 10333 20828
rect 10367 20825 10379 20859
rect 10321 20819 10379 20825
rect 4522 20748 4528 20800
rect 4580 20788 4586 20800
rect 5261 20791 5319 20797
rect 5261 20788 5273 20791
rect 4580 20760 5273 20788
rect 4580 20748 4586 20760
rect 5261 20757 5273 20760
rect 5307 20788 5319 20791
rect 5442 20788 5448 20800
rect 5307 20760 5448 20788
rect 5307 20757 5319 20760
rect 5261 20751 5319 20757
rect 5442 20748 5448 20760
rect 5500 20748 5506 20800
rect 9766 20748 9772 20800
rect 9824 20797 9830 20800
rect 9824 20791 9873 20797
rect 9824 20757 9827 20791
rect 9861 20757 9873 20791
rect 14458 20788 14464 20800
rect 14419 20760 14464 20788
rect 9824 20751 9873 20757
rect 9824 20748 9830 20751
rect 14458 20748 14464 20760
rect 14516 20748 14522 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 6178 20584 6184 20596
rect 6139 20556 6184 20584
rect 6178 20544 6184 20556
rect 6236 20544 6242 20596
rect 6641 20587 6699 20593
rect 6641 20553 6653 20587
rect 6687 20584 6699 20587
rect 6822 20584 6828 20596
rect 6687 20556 6828 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 6822 20544 6828 20556
rect 6880 20544 6886 20596
rect 7282 20584 7288 20596
rect 7243 20556 7288 20584
rect 7282 20544 7288 20556
rect 7340 20544 7346 20596
rect 10045 20587 10103 20593
rect 10045 20553 10057 20587
rect 10091 20584 10103 20587
rect 11054 20584 11060 20596
rect 10091 20556 11060 20584
rect 10091 20553 10103 20556
rect 10045 20547 10103 20553
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 13722 20544 13728 20596
rect 13780 20584 13786 20596
rect 13817 20587 13875 20593
rect 13817 20584 13829 20587
rect 13780 20556 13829 20584
rect 13780 20544 13786 20556
rect 13817 20553 13829 20556
rect 13863 20553 13875 20587
rect 13817 20547 13875 20553
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 15749 20587 15807 20593
rect 15749 20584 15761 20587
rect 15436 20556 15761 20584
rect 15436 20544 15442 20556
rect 15749 20553 15761 20556
rect 15795 20553 15807 20587
rect 15749 20547 15807 20553
rect 8202 20516 8208 20528
rect 8163 20488 8208 20516
rect 8202 20476 8208 20488
rect 8260 20476 8266 20528
rect 9950 20476 9956 20528
rect 10008 20516 10014 20528
rect 12161 20519 12219 20525
rect 12161 20516 12173 20519
rect 10008 20488 12173 20516
rect 10008 20476 10014 20488
rect 12161 20485 12173 20488
rect 12207 20516 12219 20519
rect 12250 20516 12256 20528
rect 12207 20488 12256 20516
rect 12207 20485 12219 20488
rect 12161 20479 12219 20485
rect 12250 20476 12256 20488
rect 12308 20476 12314 20528
rect 15470 20516 15476 20528
rect 15431 20488 15476 20516
rect 15470 20476 15476 20488
rect 15528 20476 15534 20528
rect 5905 20451 5963 20457
rect 5905 20417 5917 20451
rect 5951 20448 5963 20451
rect 9122 20448 9128 20460
rect 5951 20420 9128 20448
rect 5951 20417 5963 20420
rect 5905 20411 5963 20417
rect 9122 20408 9128 20420
rect 9180 20408 9186 20460
rect 10781 20451 10839 20457
rect 10781 20417 10793 20451
rect 10827 20448 10839 20451
rect 11146 20448 11152 20460
rect 10827 20420 11152 20448
rect 10827 20417 10839 20420
rect 10781 20411 10839 20417
rect 11146 20408 11152 20420
rect 11204 20448 11210 20460
rect 11471 20451 11529 20457
rect 11471 20448 11483 20451
rect 11204 20420 11483 20448
rect 11204 20408 11210 20420
rect 11471 20417 11483 20420
rect 11517 20417 11529 20451
rect 11471 20411 11529 20417
rect 11609 20451 11667 20457
rect 11609 20417 11621 20451
rect 11655 20448 11667 20451
rect 14090 20448 14096 20460
rect 11655 20420 14096 20448
rect 11655 20417 11667 20420
rect 11609 20411 11667 20417
rect 14090 20408 14096 20420
rect 14148 20408 14154 20460
rect 14734 20448 14740 20460
rect 14695 20420 14740 20448
rect 14734 20408 14740 20420
rect 14792 20408 14798 20460
rect 15838 20408 15844 20460
rect 15896 20448 15902 20460
rect 15933 20451 15991 20457
rect 15933 20448 15945 20451
rect 15896 20420 15945 20448
rect 15896 20408 15902 20420
rect 15933 20417 15945 20420
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 5077 20383 5135 20389
rect 5077 20349 5089 20383
rect 5123 20380 5135 20383
rect 5350 20380 5356 20392
rect 5123 20352 5356 20380
rect 5123 20349 5135 20352
rect 5077 20343 5135 20349
rect 5350 20340 5356 20352
rect 5408 20340 5414 20392
rect 5442 20340 5448 20392
rect 5500 20380 5506 20392
rect 5718 20380 5724 20392
rect 5500 20352 5724 20380
rect 5500 20340 5506 20352
rect 5718 20340 5724 20352
rect 5776 20340 5782 20392
rect 10410 20380 10416 20392
rect 10323 20352 10416 20380
rect 10410 20340 10416 20352
rect 10468 20380 10474 20392
rect 11384 20383 11442 20389
rect 10468 20352 11284 20380
rect 10468 20340 10474 20352
rect 7653 20315 7711 20321
rect 7653 20281 7665 20315
rect 7699 20281 7711 20315
rect 7653 20275 7711 20281
rect 7668 20244 7696 20275
rect 7742 20272 7748 20324
rect 7800 20312 7806 20324
rect 9446 20315 9504 20321
rect 9446 20312 9458 20315
rect 7800 20284 7845 20312
rect 8956 20284 9458 20312
rect 7800 20272 7806 20284
rect 8570 20244 8576 20256
rect 7668 20216 8576 20244
rect 8570 20204 8576 20216
rect 8628 20204 8634 20256
rect 8754 20204 8760 20256
rect 8812 20244 8818 20256
rect 8956 20253 8984 20284
rect 9446 20281 9458 20284
rect 9492 20312 9504 20315
rect 9950 20312 9956 20324
rect 9492 20284 9956 20312
rect 9492 20281 9504 20284
rect 9446 20275 9504 20281
rect 9950 20272 9956 20284
rect 10008 20272 10014 20324
rect 11256 20312 11284 20352
rect 11384 20349 11396 20383
rect 11430 20380 11442 20383
rect 11430 20352 11928 20380
rect 11430 20349 11442 20352
rect 11384 20343 11442 20349
rect 11609 20315 11667 20321
rect 11609 20312 11621 20315
rect 11256 20284 11621 20312
rect 11609 20281 11621 20284
rect 11655 20281 11667 20315
rect 11609 20275 11667 20281
rect 11900 20253 11928 20352
rect 12250 20340 12256 20392
rect 12308 20340 12314 20392
rect 12434 20340 12440 20392
rect 12492 20380 12498 20392
rect 12621 20383 12679 20389
rect 12621 20380 12633 20383
rect 12492 20352 12633 20380
rect 12492 20340 12498 20352
rect 12621 20349 12633 20352
rect 12667 20380 12679 20383
rect 13262 20380 13268 20392
rect 12667 20352 13268 20380
rect 12667 20349 12679 20352
rect 12621 20343 12679 20349
rect 13262 20340 13268 20352
rect 13320 20340 13326 20392
rect 13541 20383 13599 20389
rect 13541 20349 13553 20383
rect 13587 20380 13599 20383
rect 13814 20380 13820 20392
rect 13587 20352 13820 20380
rect 13587 20349 13599 20352
rect 13541 20343 13599 20349
rect 13814 20340 13820 20352
rect 13872 20340 13878 20392
rect 12268 20312 12296 20340
rect 12942 20315 13000 20321
rect 12942 20312 12954 20315
rect 12268 20284 12954 20312
rect 12942 20281 12954 20284
rect 12988 20281 13000 20315
rect 14458 20312 14464 20324
rect 14419 20284 14464 20312
rect 12942 20275 13000 20281
rect 14458 20272 14464 20284
rect 14516 20272 14522 20324
rect 14553 20315 14611 20321
rect 14553 20281 14565 20315
rect 14599 20281 14611 20315
rect 14553 20275 14611 20281
rect 8941 20247 8999 20253
rect 8941 20244 8953 20247
rect 8812 20216 8953 20244
rect 8812 20204 8818 20216
rect 8941 20213 8953 20216
rect 8987 20213 8999 20247
rect 8941 20207 8999 20213
rect 11885 20247 11943 20253
rect 11885 20213 11897 20247
rect 11931 20244 11943 20247
rect 11974 20244 11980 20256
rect 11931 20216 11980 20244
rect 11931 20213 11943 20216
rect 11885 20207 11943 20213
rect 11974 20204 11980 20216
rect 12032 20204 12038 20256
rect 14182 20244 14188 20256
rect 14143 20216 14188 20244
rect 14182 20204 14188 20216
rect 14240 20244 14246 20256
rect 14568 20244 14596 20275
rect 14240 20216 14596 20244
rect 14240 20204 14246 20216
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 5534 20000 5540 20052
rect 5592 20040 5598 20052
rect 5629 20043 5687 20049
rect 5629 20040 5641 20043
rect 5592 20012 5641 20040
rect 5592 20000 5598 20012
rect 5629 20009 5641 20012
rect 5675 20009 5687 20043
rect 5629 20003 5687 20009
rect 7101 20043 7159 20049
rect 7101 20009 7113 20043
rect 7147 20040 7159 20043
rect 7190 20040 7196 20052
rect 7147 20012 7196 20040
rect 7147 20009 7159 20012
rect 7101 20003 7159 20009
rect 7190 20000 7196 20012
rect 7248 20000 7254 20052
rect 7653 20043 7711 20049
rect 7653 20009 7665 20043
rect 7699 20040 7711 20043
rect 7742 20040 7748 20052
rect 7699 20012 7748 20040
rect 7699 20009 7711 20012
rect 7653 20003 7711 20009
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 9122 20040 9128 20052
rect 9083 20012 9128 20040
rect 9122 20000 9128 20012
rect 9180 20000 9186 20052
rect 11057 20043 11115 20049
rect 11057 20009 11069 20043
rect 11103 20040 11115 20043
rect 11882 20040 11888 20052
rect 11103 20012 11888 20040
rect 11103 20009 11115 20012
rect 11057 20003 11115 20009
rect 11882 20000 11888 20012
rect 11940 20040 11946 20052
rect 13262 20040 13268 20052
rect 11940 20012 12112 20040
rect 13223 20012 13268 20040
rect 11940 20000 11946 20012
rect 6546 19981 6552 19984
rect 6543 19972 6552 19981
rect 6507 19944 6552 19972
rect 6543 19935 6552 19944
rect 6546 19932 6552 19935
rect 6604 19932 6610 19984
rect 7208 19972 7236 20000
rect 8018 19972 8024 19984
rect 7208 19944 8024 19972
rect 8018 19932 8024 19944
rect 8076 19972 8082 19984
rect 8113 19975 8171 19981
rect 8113 19972 8125 19975
rect 8076 19944 8125 19972
rect 8076 19932 8082 19944
rect 8113 19941 8125 19944
rect 8159 19941 8171 19975
rect 8113 19935 8171 19941
rect 9950 19932 9956 19984
rect 10008 19972 10014 19984
rect 12084 19981 12112 20012
rect 13262 20000 13268 20012
rect 13320 20000 13326 20052
rect 10458 19975 10516 19981
rect 10458 19972 10470 19975
rect 10008 19944 10470 19972
rect 10008 19932 10014 19944
rect 10458 19941 10470 19944
rect 10504 19941 10516 19975
rect 10458 19935 10516 19941
rect 12069 19975 12127 19981
rect 12069 19941 12081 19975
rect 12115 19941 12127 19975
rect 12618 19972 12624 19984
rect 12579 19944 12624 19972
rect 12069 19935 12127 19941
rect 12618 19932 12624 19944
rect 12676 19932 12682 19984
rect 13814 19972 13820 19984
rect 13775 19944 13820 19972
rect 13814 19932 13820 19944
rect 13872 19932 13878 19984
rect 14090 19932 14096 19984
rect 14148 19972 14154 19984
rect 14148 19944 15399 19972
rect 14148 19932 14154 19944
rect 5074 19864 5080 19916
rect 5132 19904 5138 19916
rect 15371 19913 15399 19944
rect 5204 19907 5262 19913
rect 5204 19904 5216 19907
rect 5132 19876 5216 19904
rect 5132 19864 5138 19876
rect 5204 19873 5216 19876
rect 5250 19873 5262 19907
rect 5204 19867 5262 19873
rect 5307 19907 5365 19913
rect 5307 19873 5319 19907
rect 5353 19904 5365 19907
rect 15340 19907 15399 19913
rect 5353 19876 7328 19904
rect 5353 19873 5365 19876
rect 5307 19867 5365 19873
rect 6181 19839 6239 19845
rect 6181 19836 6193 19839
rect 6012 19808 6193 19836
rect 6012 19712 6040 19808
rect 6181 19805 6193 19808
rect 6227 19805 6239 19839
rect 7300 19836 7328 19876
rect 15340 19873 15352 19907
rect 15386 19904 15399 19907
rect 16022 19904 16028 19916
rect 15386 19876 16028 19904
rect 15386 19873 15398 19876
rect 15340 19867 15398 19873
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 8021 19839 8079 19845
rect 8021 19836 8033 19839
rect 7300 19808 8033 19836
rect 6181 19799 6239 19805
rect 8021 19805 8033 19808
rect 8067 19836 8079 19839
rect 8294 19836 8300 19848
rect 8067 19808 8300 19836
rect 8067 19805 8079 19808
rect 8021 19799 8079 19805
rect 8294 19796 8300 19808
rect 8352 19796 8358 19848
rect 10137 19839 10195 19845
rect 10137 19805 10149 19839
rect 10183 19805 10195 19839
rect 11977 19839 12035 19845
rect 11977 19836 11989 19839
rect 10137 19799 10195 19805
rect 11716 19808 11989 19836
rect 8202 19728 8208 19780
rect 8260 19768 8266 19780
rect 8570 19768 8576 19780
rect 8260 19740 8576 19768
rect 8260 19728 8266 19740
rect 8570 19728 8576 19740
rect 8628 19728 8634 19780
rect 5994 19700 6000 19712
rect 5955 19672 6000 19700
rect 5994 19660 6000 19672
rect 6052 19660 6058 19712
rect 10042 19700 10048 19712
rect 10003 19672 10048 19700
rect 10042 19660 10048 19672
rect 10100 19700 10106 19712
rect 10152 19700 10180 19799
rect 10100 19672 10180 19700
rect 10100 19660 10106 19672
rect 11606 19660 11612 19712
rect 11664 19700 11670 19712
rect 11716 19709 11744 19808
rect 11977 19805 11989 19808
rect 12023 19805 12035 19839
rect 11977 19799 12035 19805
rect 12250 19796 12256 19848
rect 12308 19836 12314 19848
rect 12897 19839 12955 19845
rect 12897 19836 12909 19839
rect 12308 19808 12909 19836
rect 12308 19796 12314 19808
rect 12897 19805 12909 19808
rect 12943 19836 12955 19839
rect 12986 19836 12992 19848
rect 12943 19808 12992 19836
rect 12943 19805 12955 19808
rect 12897 19799 12955 19805
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19805 13783 19839
rect 14366 19836 14372 19848
rect 14327 19808 14372 19836
rect 13725 19799 13783 19805
rect 13740 19768 13768 19799
rect 14366 19796 14372 19808
rect 14424 19796 14430 19848
rect 13906 19768 13912 19780
rect 13740 19740 13912 19768
rect 13906 19728 13912 19740
rect 13964 19768 13970 19780
rect 15427 19771 15485 19777
rect 15427 19768 15439 19771
rect 13964 19740 15439 19768
rect 13964 19728 13970 19740
rect 15427 19737 15439 19740
rect 15473 19737 15485 19771
rect 15427 19731 15485 19737
rect 11701 19703 11759 19709
rect 11701 19700 11713 19703
rect 11664 19672 11713 19700
rect 11664 19660 11670 19672
rect 11701 19669 11713 19672
rect 11747 19669 11759 19703
rect 11701 19663 11759 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 6273 19499 6331 19505
rect 6273 19465 6285 19499
rect 6319 19496 6331 19499
rect 6546 19496 6552 19508
rect 6319 19468 6552 19496
rect 6319 19465 6331 19468
rect 6273 19459 6331 19465
rect 6546 19456 6552 19468
rect 6604 19456 6610 19508
rect 7742 19496 7748 19508
rect 7703 19468 7748 19496
rect 7742 19456 7748 19468
rect 7800 19456 7806 19508
rect 8018 19496 8024 19508
rect 7979 19468 8024 19496
rect 8018 19456 8024 19468
rect 8076 19456 8082 19508
rect 11882 19496 11888 19508
rect 11843 19468 11888 19496
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 12986 19496 12992 19508
rect 12947 19468 12992 19496
rect 12986 19456 12992 19468
rect 13044 19456 13050 19508
rect 14093 19499 14151 19505
rect 14093 19465 14105 19499
rect 14139 19496 14151 19499
rect 14182 19496 14188 19508
rect 14139 19468 14188 19496
rect 14139 19465 14151 19468
rect 14093 19459 14151 19465
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 13814 19388 13820 19440
rect 13872 19428 13878 19440
rect 14369 19431 14427 19437
rect 14369 19428 14381 19431
rect 13872 19400 14381 19428
rect 13872 19388 13878 19400
rect 14369 19397 14381 19400
rect 14415 19397 14427 19431
rect 16022 19428 16028 19440
rect 15983 19400 16028 19428
rect 14369 19391 14427 19397
rect 16022 19388 16028 19400
rect 16080 19388 16086 19440
rect 5905 19363 5963 19369
rect 5905 19329 5917 19363
rect 5951 19360 5963 19363
rect 5994 19360 6000 19372
rect 5951 19332 6000 19360
rect 5951 19329 5963 19332
rect 5905 19323 5963 19329
rect 5994 19320 6000 19332
rect 6052 19320 6058 19372
rect 9582 19360 9588 19372
rect 9543 19332 9588 19360
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 10244 19332 13860 19360
rect 4709 19295 4767 19301
rect 4709 19261 4721 19295
rect 4755 19292 4767 19295
rect 5445 19295 5503 19301
rect 5445 19292 5457 19295
rect 4755 19264 5457 19292
rect 4755 19261 4767 19264
rect 4709 19255 4767 19261
rect 5445 19261 5457 19264
rect 5491 19292 5503 19295
rect 5534 19292 5540 19304
rect 5491 19264 5540 19292
rect 5491 19261 5503 19264
rect 5445 19255 5503 19261
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 5718 19292 5724 19304
rect 5679 19264 5724 19292
rect 5718 19252 5724 19264
rect 5776 19252 5782 19304
rect 6822 19292 6828 19304
rect 6783 19264 6828 19292
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 8294 19252 8300 19304
rect 8352 19292 8358 19304
rect 8389 19295 8447 19301
rect 8389 19292 8401 19295
rect 8352 19264 8401 19292
rect 8352 19252 8358 19264
rect 8389 19261 8401 19264
rect 8435 19261 8447 19295
rect 9030 19292 9036 19304
rect 8991 19264 9036 19292
rect 8389 19255 8447 19261
rect 9030 19252 9036 19264
rect 9088 19252 9094 19304
rect 9401 19295 9459 19301
rect 9401 19261 9413 19295
rect 9447 19292 9459 19295
rect 10244 19292 10272 19332
rect 10686 19292 10692 19304
rect 9447 19264 10272 19292
rect 10647 19264 10692 19292
rect 9447 19261 9459 19264
rect 9401 19255 9459 19261
rect 5350 19184 5356 19236
rect 5408 19224 5414 19236
rect 5736 19224 5764 19252
rect 5408 19196 5764 19224
rect 5408 19184 5414 19196
rect 6546 19184 6552 19236
rect 6604 19224 6610 19236
rect 7146 19227 7204 19233
rect 7146 19224 7158 19227
rect 6604 19196 7158 19224
rect 6604 19184 6610 19196
rect 7146 19193 7158 19196
rect 7192 19193 7204 19227
rect 9416 19224 9444 19255
rect 10686 19252 10692 19264
rect 10744 19252 10750 19304
rect 11054 19292 11060 19304
rect 11015 19264 11060 19292
rect 11054 19252 11060 19264
rect 11112 19292 11118 19304
rect 11330 19292 11336 19304
rect 11112 19264 11336 19292
rect 11112 19252 11118 19264
rect 11330 19252 11336 19264
rect 11388 19292 11394 19304
rect 11517 19295 11575 19301
rect 11517 19292 11529 19295
rect 11388 19264 11529 19292
rect 11388 19252 11394 19264
rect 11517 19261 11529 19264
rect 11563 19261 11575 19295
rect 11517 19255 11575 19261
rect 12713 19295 12771 19301
rect 12713 19261 12725 19295
rect 12759 19292 12771 19295
rect 13078 19292 13084 19304
rect 12759 19264 13084 19292
rect 12759 19261 12771 19264
rect 12713 19255 12771 19261
rect 13078 19252 13084 19264
rect 13136 19292 13142 19304
rect 13173 19295 13231 19301
rect 13173 19292 13185 19295
rect 13136 19264 13185 19292
rect 13136 19252 13142 19264
rect 13173 19261 13185 19264
rect 13219 19261 13231 19295
rect 13832 19292 13860 19332
rect 21358 19320 21364 19372
rect 21416 19360 21422 19372
rect 21634 19360 21640 19372
rect 21416 19332 21640 19360
rect 21416 19320 21422 19332
rect 21634 19320 21640 19332
rect 21692 19320 21698 19372
rect 14737 19295 14795 19301
rect 14737 19292 14749 19295
rect 13832 19264 14749 19292
rect 13173 19255 13231 19261
rect 14737 19261 14749 19264
rect 14783 19261 14795 19295
rect 14918 19292 14924 19304
rect 14879 19264 14924 19292
rect 14737 19255 14795 19261
rect 7146 19187 7204 19193
rect 8864 19196 9444 19224
rect 11241 19227 11299 19233
rect 8864 19168 8892 19196
rect 11241 19193 11253 19227
rect 11287 19224 11299 19227
rect 12434 19224 12440 19236
rect 11287 19196 12440 19224
rect 11287 19193 11299 19196
rect 11241 19187 11299 19193
rect 12434 19184 12440 19196
rect 12492 19184 12498 19236
rect 12986 19184 12992 19236
rect 13044 19224 13050 19236
rect 13494 19227 13552 19233
rect 13494 19224 13506 19227
rect 13044 19196 13506 19224
rect 13044 19184 13050 19196
rect 13494 19193 13506 19196
rect 13540 19193 13552 19227
rect 14752 19224 14780 19255
rect 14918 19252 14924 19264
rect 14976 19252 14982 19304
rect 15381 19295 15439 19301
rect 15381 19261 15393 19295
rect 15427 19261 15439 19295
rect 15381 19255 15439 19261
rect 15396 19224 15424 19255
rect 14752 19196 15424 19224
rect 13494 19187 13552 19193
rect 5074 19156 5080 19168
rect 5035 19128 5080 19156
rect 5074 19116 5080 19128
rect 5132 19116 5138 19168
rect 8846 19156 8852 19168
rect 8807 19128 8852 19156
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 10134 19156 10140 19168
rect 10095 19128 10140 19156
rect 10134 19116 10140 19128
rect 10192 19116 10198 19168
rect 15194 19156 15200 19168
rect 15155 19128 15200 19156
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 7466 18912 7472 18964
rect 7524 18952 7530 18964
rect 7524 18924 7696 18952
rect 7524 18912 7530 18924
rect 6641 18887 6699 18893
rect 6641 18853 6653 18887
rect 6687 18884 6699 18887
rect 6822 18884 6828 18896
rect 6687 18856 6828 18884
rect 6687 18853 6699 18856
rect 6641 18847 6699 18853
rect 6822 18844 6828 18856
rect 6880 18884 6886 18896
rect 7668 18893 7696 18924
rect 9674 18912 9680 18964
rect 9732 18952 9738 18964
rect 10686 18952 10692 18964
rect 9732 18924 10692 18952
rect 9732 18912 9738 18924
rect 10686 18912 10692 18924
rect 10744 18912 10750 18964
rect 11054 18912 11060 18964
rect 11112 18952 11118 18964
rect 11112 18924 12296 18952
rect 11112 18912 11118 18924
rect 7285 18887 7343 18893
rect 7285 18884 7297 18887
rect 6880 18856 7297 18884
rect 6880 18844 6886 18856
rect 7285 18853 7297 18856
rect 7331 18853 7343 18887
rect 7285 18847 7343 18853
rect 7653 18887 7711 18893
rect 7653 18853 7665 18887
rect 7699 18853 7711 18887
rect 7653 18847 7711 18853
rect 10413 18887 10471 18893
rect 10413 18853 10425 18887
rect 10459 18884 10471 18887
rect 10962 18884 10968 18896
rect 10459 18856 10968 18884
rect 10459 18853 10471 18856
rect 10413 18847 10471 18853
rect 10962 18844 10968 18856
rect 11020 18844 11026 18896
rect 11146 18844 11152 18896
rect 11204 18884 11210 18896
rect 11425 18887 11483 18893
rect 11425 18884 11437 18887
rect 11204 18856 11437 18884
rect 11204 18844 11210 18856
rect 11425 18853 11437 18856
rect 11471 18884 11483 18887
rect 12158 18884 12164 18896
rect 11471 18856 12164 18884
rect 11471 18853 11483 18856
rect 11425 18847 11483 18853
rect 12158 18844 12164 18856
rect 12216 18844 12222 18896
rect 12268 18884 12296 18924
rect 12434 18912 12440 18964
rect 12492 18952 12498 18964
rect 13078 18952 13084 18964
rect 12492 18924 12537 18952
rect 13039 18924 13084 18952
rect 12492 18912 12498 18924
rect 13078 18912 13084 18924
rect 13136 18912 13142 18964
rect 13906 18952 13912 18964
rect 13867 18924 13912 18952
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 14918 18952 14924 18964
rect 14879 18924 14924 18952
rect 14918 18912 14924 18924
rect 14976 18912 14982 18964
rect 12268 18856 13400 18884
rect 13372 18828 13400 18856
rect 5534 18776 5540 18828
rect 5592 18816 5598 18828
rect 5905 18819 5963 18825
rect 5905 18816 5917 18819
rect 5592 18788 5917 18816
rect 5592 18776 5598 18788
rect 5905 18785 5917 18788
rect 5951 18785 5963 18819
rect 6454 18816 6460 18828
rect 6415 18788 6460 18816
rect 5905 18779 5963 18785
rect 6454 18776 6460 18788
rect 6512 18776 6518 18828
rect 9953 18819 10011 18825
rect 9953 18785 9965 18819
rect 9999 18785 10011 18819
rect 9953 18779 10011 18785
rect 10229 18819 10287 18825
rect 10229 18785 10241 18819
rect 10275 18816 10287 18819
rect 10686 18816 10692 18828
rect 10275 18788 10692 18816
rect 10275 18785 10287 18788
rect 10229 18779 10287 18785
rect 7558 18748 7564 18760
rect 7519 18720 7564 18748
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 8202 18748 8208 18760
rect 8163 18720 8208 18748
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 9030 18748 9036 18760
rect 8943 18720 9036 18748
rect 9030 18708 9036 18720
rect 9088 18748 9094 18760
rect 9968 18748 9996 18779
rect 10686 18776 10692 18788
rect 10744 18816 10750 18828
rect 11054 18816 11060 18828
rect 10744 18788 11060 18816
rect 10744 18776 10750 18788
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 13081 18819 13139 18825
rect 13081 18785 13093 18819
rect 13127 18785 13139 18819
rect 13354 18816 13360 18828
rect 13315 18788 13360 18816
rect 13081 18779 13139 18785
rect 10962 18748 10968 18760
rect 9088 18720 10968 18748
rect 9088 18708 9094 18720
rect 10962 18708 10968 18720
rect 11020 18708 11026 18760
rect 11330 18748 11336 18760
rect 11291 18720 11336 18748
rect 11330 18708 11336 18720
rect 11388 18708 11394 18760
rect 11606 18748 11612 18760
rect 11567 18720 11612 18748
rect 11606 18708 11612 18720
rect 11664 18708 11670 18760
rect 13096 18748 13124 18779
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 15378 18825 15384 18828
rect 15356 18819 15384 18825
rect 15356 18785 15368 18819
rect 15356 18779 15384 18785
rect 15378 18776 15384 18779
rect 15436 18776 15442 18828
rect 13170 18748 13176 18760
rect 13083 18720 13176 18748
rect 13170 18708 13176 18720
rect 13228 18748 13234 18760
rect 14918 18748 14924 18760
rect 13228 18720 14924 18748
rect 13228 18708 13234 18720
rect 14918 18708 14924 18720
rect 14976 18708 14982 18760
rect 5718 18640 5724 18692
rect 5776 18640 5782 18692
rect 5261 18615 5319 18621
rect 5261 18581 5273 18615
rect 5307 18612 5319 18615
rect 5736 18612 5764 18640
rect 6362 18612 6368 18624
rect 5307 18584 6368 18612
rect 5307 18581 5319 18584
rect 5261 18575 5319 18581
rect 6362 18572 6368 18584
rect 6420 18572 6426 18624
rect 6914 18612 6920 18624
rect 6875 18584 6920 18612
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 14274 18612 14280 18624
rect 14235 18584 14280 18612
rect 14274 18572 14280 18584
rect 14332 18572 14338 18624
rect 15427 18615 15485 18621
rect 15427 18581 15439 18615
rect 15473 18612 15485 18615
rect 15930 18612 15936 18624
rect 15473 18584 15936 18612
rect 15473 18581 15485 18584
rect 15427 18575 15485 18581
rect 15930 18572 15936 18584
rect 15988 18572 15994 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 5166 18368 5172 18420
rect 5224 18408 5230 18420
rect 5534 18408 5540 18420
rect 5224 18380 5540 18408
rect 5224 18368 5230 18380
rect 5534 18368 5540 18380
rect 5592 18408 5598 18420
rect 5905 18411 5963 18417
rect 5905 18408 5917 18411
rect 5592 18380 5917 18408
rect 5592 18368 5598 18380
rect 5905 18377 5917 18380
rect 5951 18377 5963 18411
rect 6546 18408 6552 18420
rect 6507 18380 6552 18408
rect 5905 18371 5963 18377
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 7466 18368 7472 18420
rect 7524 18408 7530 18420
rect 7745 18411 7803 18417
rect 7745 18408 7757 18411
rect 7524 18380 7757 18408
rect 7524 18368 7530 18380
rect 7745 18377 7757 18380
rect 7791 18408 7803 18411
rect 8021 18411 8079 18417
rect 8021 18408 8033 18411
rect 7791 18380 8033 18408
rect 7791 18377 7803 18380
rect 7745 18371 7803 18377
rect 8021 18377 8033 18380
rect 8067 18377 8079 18411
rect 8021 18371 8079 18377
rect 10045 18411 10103 18417
rect 10045 18377 10057 18411
rect 10091 18408 10103 18411
rect 11146 18408 11152 18420
rect 10091 18380 11152 18408
rect 10091 18377 10103 18380
rect 10045 18371 10103 18377
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 11330 18368 11336 18420
rect 11388 18408 11394 18420
rect 11471 18411 11529 18417
rect 11471 18408 11483 18411
rect 11388 18380 11483 18408
rect 11388 18368 11394 18380
rect 11471 18377 11483 18380
rect 11517 18377 11529 18411
rect 11882 18408 11888 18420
rect 11843 18380 11888 18408
rect 11471 18371 11529 18377
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 13354 18368 13360 18420
rect 13412 18408 13418 18420
rect 13633 18411 13691 18417
rect 13633 18408 13645 18411
rect 13412 18380 13645 18408
rect 13412 18368 13418 18380
rect 13633 18377 13645 18380
rect 13679 18377 13691 18411
rect 15378 18408 15384 18420
rect 15339 18380 15384 18408
rect 13633 18371 13691 18377
rect 15378 18368 15384 18380
rect 15436 18368 15442 18420
rect 5629 18275 5687 18281
rect 5629 18241 5641 18275
rect 5675 18272 5687 18275
rect 6454 18272 6460 18284
rect 5675 18244 6460 18272
rect 5675 18241 5687 18244
rect 5629 18235 5687 18241
rect 6454 18232 6460 18244
rect 6512 18232 6518 18284
rect 12434 18232 12440 18284
rect 12492 18272 12498 18284
rect 12492 18244 12537 18272
rect 12492 18232 12498 18244
rect 14366 18232 14372 18284
rect 14424 18272 14430 18284
rect 14553 18275 14611 18281
rect 14553 18272 14565 18275
rect 14424 18244 14565 18272
rect 14424 18232 14430 18244
rect 14553 18241 14565 18244
rect 14599 18241 14611 18275
rect 14553 18235 14611 18241
rect 5534 18164 5540 18216
rect 5592 18204 5598 18216
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 5592 18176 6837 18204
rect 5592 18164 5598 18176
rect 6825 18173 6837 18176
rect 6871 18204 6883 18207
rect 6914 18204 6920 18216
rect 6871 18176 6920 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 9125 18207 9183 18213
rect 9125 18173 9137 18207
rect 9171 18204 9183 18207
rect 9214 18204 9220 18216
rect 9171 18176 9220 18204
rect 9171 18173 9183 18176
rect 9125 18167 9183 18173
rect 9214 18164 9220 18176
rect 9272 18164 9278 18216
rect 10413 18207 10471 18213
rect 10413 18173 10425 18207
rect 10459 18204 10471 18207
rect 10686 18204 10692 18216
rect 10459 18176 10692 18204
rect 10459 18173 10471 18176
rect 10413 18167 10471 18173
rect 10686 18164 10692 18176
rect 10744 18164 10750 18216
rect 11400 18207 11458 18213
rect 11400 18173 11412 18207
rect 11446 18204 11458 18207
rect 11882 18204 11888 18216
rect 11446 18176 11888 18204
rect 11446 18173 11458 18176
rect 11400 18167 11458 18173
rect 11882 18164 11888 18176
rect 11940 18164 11946 18216
rect 12176 18176 12848 18204
rect 6546 18096 6552 18148
rect 6604 18136 6610 18148
rect 7146 18139 7204 18145
rect 7146 18136 7158 18139
rect 6604 18108 7158 18136
rect 6604 18096 6610 18108
rect 7146 18105 7158 18108
rect 7192 18136 7204 18139
rect 7834 18136 7840 18148
rect 7192 18108 7840 18136
rect 7192 18105 7204 18108
rect 7146 18099 7204 18105
rect 7834 18096 7840 18108
rect 7892 18136 7898 18148
rect 8754 18136 8760 18148
rect 7892 18108 8760 18136
rect 7892 18096 7898 18108
rect 8754 18096 8760 18108
rect 8812 18136 8818 18148
rect 8941 18139 8999 18145
rect 8941 18136 8953 18139
rect 8812 18108 8953 18136
rect 8812 18096 8818 18108
rect 8941 18105 8953 18108
rect 8987 18136 8999 18139
rect 9446 18139 9504 18145
rect 9446 18136 9458 18139
rect 8987 18108 9458 18136
rect 8987 18105 8999 18108
rect 8941 18099 8999 18105
rect 9446 18105 9458 18108
rect 9492 18136 9504 18139
rect 10134 18136 10140 18148
rect 9492 18108 10140 18136
rect 9492 18105 9504 18108
rect 9446 18099 9504 18105
rect 10134 18096 10140 18108
rect 10192 18096 10198 18148
rect 12176 18080 12204 18176
rect 12820 18145 12848 18176
rect 13262 18164 13268 18216
rect 13320 18204 13326 18216
rect 13357 18207 13415 18213
rect 13357 18204 13369 18207
rect 13320 18176 13369 18204
rect 13320 18164 13326 18176
rect 13357 18173 13369 18176
rect 13403 18204 13415 18207
rect 14001 18207 14059 18213
rect 14001 18204 14013 18207
rect 13403 18176 14013 18204
rect 13403 18173 13415 18176
rect 13357 18167 13415 18173
rect 12799 18139 12857 18145
rect 12799 18105 12811 18139
rect 12845 18105 12857 18139
rect 12799 18099 12857 18105
rect 10781 18071 10839 18077
rect 10781 18037 10793 18071
rect 10827 18068 10839 18071
rect 10962 18068 10968 18080
rect 10827 18040 10968 18068
rect 10827 18037 10839 18040
rect 10781 18031 10839 18037
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 12158 18068 12164 18080
rect 12119 18040 12164 18068
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 13740 18068 13768 18176
rect 14001 18173 14013 18176
rect 14047 18173 14059 18207
rect 14001 18167 14059 18173
rect 16117 18207 16175 18213
rect 16117 18173 16129 18207
rect 16163 18204 16175 18207
rect 16574 18204 16580 18216
rect 16163 18176 16580 18204
rect 16163 18173 16175 18176
rect 16117 18167 16175 18173
rect 16574 18164 16580 18176
rect 16632 18164 16638 18216
rect 13814 18096 13820 18148
rect 13872 18136 13878 18148
rect 14274 18136 14280 18148
rect 13872 18108 14280 18136
rect 13872 18096 13878 18108
rect 14274 18096 14280 18108
rect 14332 18096 14338 18148
rect 14369 18139 14427 18145
rect 14369 18105 14381 18139
rect 14415 18105 14427 18139
rect 14369 18099 14427 18105
rect 14384 18068 14412 18099
rect 13740 18040 14412 18068
rect 16669 18071 16727 18077
rect 16669 18037 16681 18071
rect 16715 18068 16727 18071
rect 16758 18068 16764 18080
rect 16715 18040 16764 18068
rect 16715 18037 16727 18040
rect 16669 18031 16727 18037
rect 16758 18028 16764 18040
rect 16816 18028 16822 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 7098 17824 7104 17876
rect 7156 17864 7162 17876
rect 7377 17867 7435 17873
rect 7377 17864 7389 17867
rect 7156 17836 7389 17864
rect 7156 17824 7162 17836
rect 7377 17833 7389 17836
rect 7423 17833 7435 17867
rect 7377 17827 7435 17833
rect 7558 17824 7564 17876
rect 7616 17864 7622 17876
rect 7653 17867 7711 17873
rect 7653 17864 7665 17867
rect 7616 17836 7665 17864
rect 7616 17824 7622 17836
rect 7653 17833 7665 17836
rect 7699 17864 7711 17867
rect 8343 17867 8401 17873
rect 8343 17864 8355 17867
rect 7699 17836 8355 17864
rect 7699 17833 7711 17836
rect 7653 17827 7711 17833
rect 8343 17833 8355 17836
rect 8389 17833 8401 17867
rect 8343 17827 8401 17833
rect 10597 17867 10655 17873
rect 10597 17833 10609 17867
rect 10643 17864 10655 17867
rect 10870 17864 10876 17876
rect 10643 17836 10876 17864
rect 10643 17833 10655 17836
rect 10597 17827 10655 17833
rect 10870 17824 10876 17836
rect 10928 17824 10934 17876
rect 11330 17864 11336 17876
rect 11291 17836 11336 17864
rect 11330 17824 11336 17836
rect 11388 17824 11394 17876
rect 12805 17867 12863 17873
rect 12805 17833 12817 17867
rect 12851 17833 12863 17867
rect 13170 17864 13176 17876
rect 13131 17836 13176 17864
rect 12805 17827 12863 17833
rect 6546 17756 6552 17808
rect 6604 17796 6610 17808
rect 6778 17799 6836 17805
rect 6778 17796 6790 17799
rect 6604 17768 6790 17796
rect 6604 17756 6610 17768
rect 6778 17765 6790 17768
rect 6824 17765 6836 17799
rect 6778 17759 6836 17765
rect 10039 17799 10097 17805
rect 10039 17765 10051 17799
rect 10085 17796 10097 17799
rect 10134 17796 10140 17808
rect 10085 17768 10140 17796
rect 10085 17765 10097 17768
rect 10039 17759 10097 17765
rect 10134 17756 10140 17768
rect 10192 17756 10198 17808
rect 12158 17756 12164 17808
rect 12216 17805 12222 17808
rect 12216 17799 12264 17805
rect 12216 17765 12218 17799
rect 12252 17765 12264 17799
rect 12820 17796 12848 17827
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 15470 17864 15476 17876
rect 13832 17836 15476 17864
rect 13446 17796 13452 17808
rect 12820 17768 13452 17796
rect 12216 17759 12264 17765
rect 12216 17756 12222 17759
rect 13446 17756 13452 17768
rect 13504 17796 13510 17808
rect 13832 17805 13860 17836
rect 15470 17824 15476 17836
rect 15528 17824 15534 17876
rect 16206 17864 16212 17876
rect 16167 17836 16212 17864
rect 16206 17824 16212 17836
rect 16264 17824 16270 17876
rect 13817 17799 13875 17805
rect 13817 17796 13829 17799
rect 13504 17768 13829 17796
rect 13504 17756 13510 17768
rect 13817 17765 13829 17768
rect 13863 17765 13875 17799
rect 14366 17796 14372 17808
rect 14327 17768 14372 17796
rect 13817 17759 13875 17765
rect 14366 17756 14372 17768
rect 14424 17756 14430 17808
rect 16574 17756 16580 17808
rect 16632 17796 16638 17808
rect 16669 17799 16727 17805
rect 16669 17796 16681 17799
rect 16632 17768 16681 17796
rect 16632 17756 16638 17768
rect 16669 17765 16681 17768
rect 16715 17765 16727 17799
rect 16669 17759 16727 17765
rect 5166 17728 5172 17740
rect 5127 17700 5172 17728
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 5350 17728 5356 17740
rect 5311 17700 5356 17728
rect 5350 17688 5356 17700
rect 5408 17688 5414 17740
rect 8272 17731 8330 17737
rect 8272 17697 8284 17731
rect 8318 17728 8330 17731
rect 8662 17728 8668 17740
rect 8318 17700 8668 17728
rect 8318 17697 8330 17700
rect 8272 17691 8330 17697
rect 8662 17688 8668 17700
rect 8720 17688 8726 17740
rect 15378 17737 15384 17740
rect 15356 17731 15384 17737
rect 15356 17697 15368 17731
rect 15356 17691 15384 17697
rect 15378 17688 15384 17691
rect 15436 17688 15442 17740
rect 5442 17660 5448 17672
rect 5403 17632 5448 17660
rect 5442 17620 5448 17632
rect 5500 17620 5506 17672
rect 6454 17660 6460 17672
rect 6415 17632 6460 17660
rect 6454 17620 6460 17632
rect 6512 17620 6518 17672
rect 9674 17660 9680 17672
rect 9635 17632 9680 17660
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 11790 17620 11796 17672
rect 11848 17660 11854 17672
rect 11885 17663 11943 17669
rect 11885 17660 11897 17663
rect 11848 17632 11897 17660
rect 11848 17620 11854 17632
rect 11885 17629 11897 17632
rect 11931 17629 11943 17663
rect 13722 17660 13728 17672
rect 13683 17632 13728 17660
rect 11885 17623 11943 17629
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 15746 17620 15752 17672
rect 15804 17660 15810 17672
rect 16577 17663 16635 17669
rect 16577 17660 16589 17663
rect 15804 17632 16589 17660
rect 15804 17620 15810 17632
rect 16577 17629 16589 17632
rect 16623 17629 16635 17663
rect 16577 17623 16635 17629
rect 16666 17620 16672 17672
rect 16724 17660 16730 17672
rect 18049 17663 18107 17669
rect 18049 17660 18061 17663
rect 16724 17632 18061 17660
rect 16724 17620 16730 17632
rect 18049 17629 18061 17632
rect 18095 17629 18107 17663
rect 18049 17623 18107 17629
rect 16942 17552 16948 17604
rect 17000 17592 17006 17604
rect 17129 17595 17187 17601
rect 17129 17592 17141 17595
rect 17000 17564 17141 17592
rect 17000 17552 17006 17564
rect 17129 17561 17141 17564
rect 17175 17561 17187 17595
rect 17129 17555 17187 17561
rect 9214 17524 9220 17536
rect 9175 17496 9220 17524
rect 9214 17484 9220 17496
rect 9272 17484 9278 17536
rect 10962 17524 10968 17536
rect 10923 17496 10968 17524
rect 10962 17484 10968 17496
rect 11020 17484 11026 17536
rect 15427 17527 15485 17533
rect 15427 17493 15439 17527
rect 15473 17524 15485 17527
rect 16114 17524 16120 17536
rect 15473 17496 16120 17524
rect 15473 17493 15485 17496
rect 15427 17487 15485 17493
rect 16114 17484 16120 17496
rect 16172 17484 16178 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 5166 17280 5172 17332
rect 5224 17320 5230 17332
rect 5261 17323 5319 17329
rect 5261 17320 5273 17323
rect 5224 17292 5273 17320
rect 5224 17280 5230 17292
rect 5261 17289 5273 17292
rect 5307 17289 5319 17323
rect 6270 17320 6276 17332
rect 6231 17292 6276 17320
rect 5261 17283 5319 17289
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 6638 17320 6644 17332
rect 6599 17292 6644 17320
rect 6638 17280 6644 17292
rect 6696 17280 6702 17332
rect 7098 17280 7104 17332
rect 7156 17320 7162 17332
rect 7377 17323 7435 17329
rect 7377 17320 7389 17323
rect 7156 17292 7389 17320
rect 7156 17280 7162 17292
rect 7377 17289 7389 17292
rect 7423 17320 7435 17323
rect 7742 17320 7748 17332
rect 7423 17292 7748 17320
rect 7423 17289 7435 17292
rect 7377 17283 7435 17289
rect 7742 17280 7748 17292
rect 7800 17280 7806 17332
rect 10134 17320 10140 17332
rect 10095 17292 10140 17320
rect 10134 17280 10140 17292
rect 10192 17280 10198 17332
rect 10689 17323 10747 17329
rect 10689 17289 10701 17323
rect 10735 17320 10747 17323
rect 10870 17320 10876 17332
rect 10735 17292 10876 17320
rect 10735 17289 10747 17292
rect 10689 17283 10747 17289
rect 10870 17280 10876 17292
rect 10928 17280 10934 17332
rect 11885 17323 11943 17329
rect 11885 17320 11897 17323
rect 11158 17292 11897 17320
rect 4985 17255 5043 17261
rect 4985 17221 4997 17255
rect 5031 17252 5043 17255
rect 5350 17252 5356 17264
rect 5031 17224 5356 17252
rect 5031 17221 5043 17224
rect 4985 17215 5043 17221
rect 5350 17212 5356 17224
rect 5408 17212 5414 17264
rect 6288 17184 6316 17280
rect 8202 17252 8208 17264
rect 8163 17224 8208 17252
rect 8202 17212 8208 17224
rect 8260 17212 8266 17264
rect 8662 17252 8668 17264
rect 8623 17224 8668 17252
rect 8662 17212 8668 17224
rect 8720 17212 8726 17264
rect 10152 17252 10180 17280
rect 11158 17252 11186 17292
rect 11885 17289 11897 17292
rect 11931 17320 11943 17323
rect 12158 17320 12164 17332
rect 11931 17292 12164 17320
rect 11931 17289 11943 17292
rect 11885 17283 11943 17289
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 13446 17320 13452 17332
rect 13407 17292 13452 17320
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 13679 17323 13737 17329
rect 13679 17289 13691 17323
rect 13725 17320 13737 17323
rect 13814 17320 13820 17332
rect 13725 17292 13820 17320
rect 13725 17289 13737 17292
rect 13679 17283 13737 17289
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 14461 17323 14519 17329
rect 14461 17289 14473 17323
rect 14507 17320 14519 17323
rect 14642 17320 14648 17332
rect 14507 17292 14648 17320
rect 14507 17289 14519 17292
rect 14461 17283 14519 17289
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 15378 17320 15384 17332
rect 15339 17292 15384 17320
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 10152 17224 11186 17252
rect 11425 17255 11483 17261
rect 11425 17221 11437 17255
rect 11471 17252 11483 17255
rect 11606 17252 11612 17264
rect 11471 17224 11612 17252
rect 11471 17221 11483 17224
rect 11425 17215 11483 17221
rect 11606 17212 11612 17224
rect 11664 17212 11670 17264
rect 16206 17212 16212 17264
rect 16264 17252 16270 17264
rect 16264 17224 16344 17252
rect 16264 17212 16270 17224
rect 5736 17156 6316 17184
rect 10873 17187 10931 17193
rect 5736 17125 5764 17156
rect 10873 17153 10885 17187
rect 10919 17184 10931 17187
rect 10962 17184 10968 17196
rect 10919 17156 10968 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 10962 17144 10968 17156
rect 11020 17184 11026 17196
rect 16316 17193 16344 17224
rect 12575 17187 12633 17193
rect 12575 17184 12587 17187
rect 11020 17156 12587 17184
rect 11020 17144 11026 17156
rect 12575 17153 12587 17156
rect 12621 17153 12633 17187
rect 12575 17147 12633 17153
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17153 16359 17187
rect 16301 17147 16359 17153
rect 5736 17119 5814 17125
rect 5736 17088 5768 17119
rect 5756 17085 5768 17088
rect 5802 17085 5814 17119
rect 5756 17079 5814 17085
rect 5859 17119 5917 17125
rect 5859 17085 5871 17119
rect 5905 17116 5917 17119
rect 6730 17116 6736 17128
rect 5905 17088 6736 17116
rect 5905 17085 5917 17088
rect 5859 17079 5917 17085
rect 6730 17076 6736 17088
rect 6788 17076 6794 17128
rect 9033 17119 9091 17125
rect 9033 17085 9045 17119
rect 9079 17116 9091 17119
rect 9401 17119 9459 17125
rect 9401 17116 9413 17119
rect 9079 17088 9413 17116
rect 9079 17085 9091 17088
rect 9033 17079 9091 17085
rect 9401 17085 9413 17088
rect 9447 17116 9459 17119
rect 9490 17116 9496 17128
rect 9447 17088 9496 17116
rect 9447 17085 9459 17088
rect 9401 17079 9459 17085
rect 9490 17076 9496 17088
rect 9548 17076 9554 17128
rect 9582 17076 9588 17128
rect 9640 17116 9646 17128
rect 13630 17125 13636 17128
rect 12488 17119 12546 17125
rect 9640 17088 9685 17116
rect 9640 17076 9646 17088
rect 12488 17085 12500 17119
rect 12534 17116 12546 17119
rect 13592 17119 13636 17125
rect 12534 17088 13032 17116
rect 12534 17085 12546 17088
rect 12488 17079 12546 17085
rect 6454 17008 6460 17060
rect 6512 17048 6518 17060
rect 7009 17051 7067 17057
rect 7009 17048 7021 17051
rect 6512 17020 7021 17048
rect 6512 17008 6518 17020
rect 7009 17017 7021 17020
rect 7055 17017 7067 17051
rect 7650 17048 7656 17060
rect 7611 17020 7656 17048
rect 7009 17011 7067 17017
rect 7650 17008 7656 17020
rect 7708 17008 7714 17060
rect 7742 17008 7748 17060
rect 7800 17048 7806 17060
rect 7800 17020 7845 17048
rect 7800 17008 7806 17020
rect 10870 17008 10876 17060
rect 10928 17048 10934 17060
rect 10965 17051 11023 17057
rect 10965 17048 10977 17051
rect 10928 17020 10977 17048
rect 10928 17008 10934 17020
rect 10965 17017 10977 17020
rect 11011 17017 11023 17051
rect 10965 17011 11023 17017
rect 13004 16992 13032 17088
rect 13592 17085 13604 17119
rect 13688 17116 13694 17128
rect 14090 17116 14096 17128
rect 13688 17088 14096 17116
rect 13592 17079 13636 17085
rect 13630 17076 13636 17079
rect 13688 17076 13694 17088
rect 14090 17076 14096 17088
rect 14148 17076 14154 17128
rect 14642 17125 14648 17128
rect 14620 17119 14648 17125
rect 14620 17085 14632 17119
rect 14620 17079 14648 17085
rect 14642 17076 14648 17079
rect 14700 17076 14706 17128
rect 17034 17076 17040 17128
rect 17092 17116 17098 17128
rect 17865 17119 17923 17125
rect 17865 17116 17877 17119
rect 17092 17088 17877 17116
rect 17092 17076 17098 17088
rect 17865 17085 17877 17088
rect 17911 17116 17923 17119
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 17911 17088 18153 17116
rect 17911 17085 17923 17088
rect 17865 17079 17923 17085
rect 18141 17085 18153 17088
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 16117 17051 16175 17057
rect 16117 17017 16129 17051
rect 16163 17048 16175 17051
rect 16393 17051 16451 17057
rect 16393 17048 16405 17051
rect 16163 17020 16405 17048
rect 16163 17017 16175 17020
rect 16117 17011 16175 17017
rect 16393 17017 16405 17020
rect 16439 17048 16451 17051
rect 16758 17048 16764 17060
rect 16439 17020 16764 17048
rect 16439 17017 16451 17020
rect 16393 17011 16451 17017
rect 16758 17008 16764 17020
rect 16816 17008 16822 17060
rect 16942 17048 16948 17060
rect 16903 17020 16948 17048
rect 16942 17008 16948 17020
rect 17000 17008 17006 17060
rect 18046 17048 18052 17060
rect 18007 17020 18052 17048
rect 18046 17008 18052 17020
rect 18104 17008 18110 17060
rect 9214 16980 9220 16992
rect 9175 16952 9220 16980
rect 9214 16940 9220 16952
rect 9272 16940 9278 16992
rect 12986 16980 12992 16992
rect 12947 16952 12992 16980
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 14458 16940 14464 16992
rect 14516 16980 14522 16992
rect 14691 16983 14749 16989
rect 14691 16980 14703 16983
rect 14516 16952 14703 16980
rect 14516 16940 14522 16952
rect 14691 16949 14703 16952
rect 14737 16949 14749 16983
rect 15746 16980 15752 16992
rect 15707 16952 15752 16980
rect 14691 16943 14749 16949
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 16482 16940 16488 16992
rect 16540 16980 16546 16992
rect 17313 16983 17371 16989
rect 17313 16980 17325 16983
rect 16540 16952 17325 16980
rect 16540 16940 16546 16952
rect 17313 16949 17325 16952
rect 17359 16980 17371 16983
rect 18322 16980 18328 16992
rect 17359 16952 18328 16980
rect 17359 16949 17371 16952
rect 17313 16943 17371 16949
rect 18322 16940 18328 16952
rect 18380 16940 18386 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 4338 16776 4344 16788
rect 4299 16748 4344 16776
rect 4338 16736 4344 16748
rect 4396 16736 4402 16788
rect 5166 16736 5172 16788
rect 5224 16776 5230 16788
rect 5997 16779 6055 16785
rect 5997 16776 6009 16779
rect 5224 16748 6009 16776
rect 5224 16736 5230 16748
rect 5997 16745 6009 16748
rect 6043 16776 6055 16779
rect 6178 16776 6184 16788
rect 6043 16748 6184 16776
rect 6043 16745 6055 16748
rect 5997 16739 6055 16745
rect 6178 16736 6184 16748
rect 6236 16736 6242 16788
rect 6454 16776 6460 16788
rect 6415 16748 6460 16776
rect 6454 16736 6460 16748
rect 6512 16736 6518 16788
rect 8846 16776 8852 16788
rect 8588 16748 8852 16776
rect 5307 16711 5365 16717
rect 5307 16677 5319 16711
rect 5353 16708 5365 16711
rect 7561 16711 7619 16717
rect 7561 16708 7573 16711
rect 5353 16680 7573 16708
rect 5353 16677 5365 16680
rect 5307 16671 5365 16677
rect 7561 16677 7573 16680
rect 7607 16708 7619 16711
rect 7650 16708 7656 16720
rect 7607 16680 7656 16708
rect 7607 16677 7619 16680
rect 7561 16671 7619 16677
rect 7650 16668 7656 16680
rect 7708 16668 7714 16720
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16640 4215 16643
rect 4246 16640 4252 16652
rect 4203 16612 4252 16640
rect 4203 16609 4215 16612
rect 4157 16603 4215 16609
rect 4246 16600 4252 16612
rect 4304 16600 4310 16652
rect 5166 16600 5172 16652
rect 5224 16649 5230 16652
rect 5224 16643 5262 16649
rect 5250 16609 5262 16643
rect 6178 16640 6184 16652
rect 6139 16612 6184 16640
rect 5224 16603 5262 16609
rect 5224 16600 5230 16603
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 6733 16643 6791 16649
rect 6733 16609 6745 16643
rect 6779 16640 6791 16643
rect 7926 16640 7932 16652
rect 6779 16612 7932 16640
rect 6779 16609 6791 16612
rect 6733 16603 6791 16609
rect 7926 16600 7932 16612
rect 7984 16640 7990 16652
rect 8021 16643 8079 16649
rect 8021 16640 8033 16643
rect 7984 16612 8033 16640
rect 7984 16600 7990 16612
rect 8021 16609 8033 16612
rect 8067 16609 8079 16643
rect 8021 16603 8079 16609
rect 8478 16600 8484 16652
rect 8536 16640 8542 16652
rect 8588 16649 8616 16748
rect 8846 16736 8852 16748
rect 8904 16776 8910 16788
rect 9217 16779 9275 16785
rect 9217 16776 9229 16779
rect 8904 16748 9229 16776
rect 8904 16736 8910 16748
rect 9217 16745 9229 16748
rect 9263 16776 9275 16779
rect 9582 16776 9588 16788
rect 9263 16748 9588 16776
rect 9263 16745 9275 16748
rect 9217 16739 9275 16745
rect 9582 16736 9588 16748
rect 9640 16776 9646 16788
rect 11146 16776 11152 16788
rect 9640 16748 11152 16776
rect 9640 16736 9646 16748
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 13587 16779 13645 16785
rect 13587 16745 13599 16779
rect 13633 16776 13645 16779
rect 13722 16776 13728 16788
rect 13633 16748 13728 16776
rect 13633 16745 13645 16748
rect 13587 16739 13645 16745
rect 13722 16736 13728 16748
rect 13780 16776 13786 16788
rect 13909 16779 13967 16785
rect 13909 16776 13921 16779
rect 13780 16748 13921 16776
rect 13780 16736 13786 16748
rect 13909 16745 13921 16748
rect 13955 16745 13967 16779
rect 18782 16776 18788 16788
rect 13909 16739 13967 16745
rect 18248 16748 18788 16776
rect 8757 16711 8815 16717
rect 8757 16677 8769 16711
rect 8803 16708 8815 16711
rect 9674 16708 9680 16720
rect 8803 16680 9680 16708
rect 8803 16677 8815 16680
rect 8757 16671 8815 16677
rect 9674 16668 9680 16680
rect 9732 16708 9738 16720
rect 9861 16711 9919 16717
rect 9861 16708 9873 16711
rect 9732 16680 9873 16708
rect 9732 16668 9738 16680
rect 9861 16677 9873 16680
rect 9907 16677 9919 16711
rect 9861 16671 9919 16677
rect 11057 16711 11115 16717
rect 11057 16677 11069 16711
rect 11103 16708 11115 16711
rect 11701 16711 11759 16717
rect 11701 16708 11713 16711
rect 11103 16680 11713 16708
rect 11103 16677 11115 16680
rect 11057 16671 11115 16677
rect 11701 16677 11713 16680
rect 11747 16708 11759 16711
rect 11790 16708 11796 16720
rect 11747 16680 11796 16708
rect 11747 16677 11759 16680
rect 11701 16671 11759 16677
rect 11790 16668 11796 16680
rect 11848 16668 11854 16720
rect 11974 16708 11980 16720
rect 11935 16680 11980 16708
rect 11974 16668 11980 16680
rect 12032 16668 12038 16720
rect 12069 16711 12127 16717
rect 12069 16677 12081 16711
rect 12115 16708 12127 16711
rect 12342 16708 12348 16720
rect 12115 16680 12348 16708
rect 12115 16677 12127 16680
rect 12069 16671 12127 16677
rect 12342 16668 12348 16680
rect 12400 16668 12406 16720
rect 15194 16668 15200 16720
rect 15252 16708 15258 16720
rect 15427 16711 15485 16717
rect 15427 16708 15439 16711
rect 15252 16680 15439 16708
rect 15252 16668 15258 16680
rect 15427 16677 15439 16680
rect 15473 16677 15485 16711
rect 16666 16708 16672 16720
rect 16627 16680 16672 16708
rect 15427 16671 15485 16677
rect 16666 16668 16672 16680
rect 16724 16668 16730 16720
rect 16758 16668 16764 16720
rect 16816 16708 16822 16720
rect 17310 16708 17316 16720
rect 16816 16680 17316 16708
rect 16816 16668 16822 16680
rect 17310 16668 17316 16680
rect 17368 16668 17374 16720
rect 18248 16717 18276 16748
rect 18782 16736 18788 16748
rect 18840 16776 18846 16788
rect 19843 16779 19901 16785
rect 19843 16776 19855 16779
rect 18840 16748 19855 16776
rect 18840 16736 18846 16748
rect 19843 16745 19855 16748
rect 19889 16745 19901 16779
rect 19843 16739 19901 16745
rect 18233 16711 18291 16717
rect 18233 16677 18245 16711
rect 18279 16677 18291 16711
rect 18233 16671 18291 16677
rect 18322 16668 18328 16720
rect 18380 16708 18386 16720
rect 18380 16680 18425 16708
rect 18380 16668 18386 16680
rect 8573 16643 8631 16649
rect 8573 16640 8585 16643
rect 8536 16612 8585 16640
rect 8536 16600 8542 16612
rect 8573 16609 8585 16612
rect 8619 16609 8631 16643
rect 8573 16603 8631 16609
rect 10134 16600 10140 16652
rect 10192 16640 10198 16652
rect 10321 16643 10379 16649
rect 10321 16640 10333 16643
rect 10192 16612 10333 16640
rect 10192 16600 10198 16612
rect 10321 16609 10333 16612
rect 10367 16609 10379 16643
rect 10321 16603 10379 16609
rect 10686 16600 10692 16652
rect 10744 16640 10750 16652
rect 10781 16643 10839 16649
rect 10781 16640 10793 16643
rect 10744 16612 10793 16640
rect 10744 16600 10750 16612
rect 10781 16609 10793 16612
rect 10827 16609 10839 16643
rect 10781 16603 10839 16609
rect 13446 16600 13452 16652
rect 13504 16649 13510 16652
rect 13504 16643 13542 16649
rect 13530 16609 13542 16643
rect 13504 16603 13542 16609
rect 13504 16600 13510 16603
rect 15286 16600 15292 16652
rect 15344 16649 15350 16652
rect 15344 16643 15382 16649
rect 15370 16609 15382 16643
rect 15344 16603 15382 16609
rect 15344 16600 15350 16603
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 19740 16643 19798 16649
rect 19740 16640 19752 16643
rect 19484 16612 19752 16640
rect 19484 16600 19490 16612
rect 19740 16609 19752 16612
rect 19786 16609 19798 16643
rect 19740 16603 19798 16609
rect 11330 16532 11336 16584
rect 11388 16572 11394 16584
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 11388 16544 12265 16572
rect 11388 16532 11394 16544
rect 12253 16541 12265 16544
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 17313 16575 17371 16581
rect 17313 16541 17325 16575
rect 17359 16572 17371 16575
rect 17957 16575 18015 16581
rect 17957 16572 17969 16575
rect 17359 16544 17969 16572
rect 17359 16541 17371 16544
rect 17313 16535 17371 16541
rect 17957 16541 17969 16544
rect 18003 16541 18015 16575
rect 17957 16535 18015 16541
rect 18509 16575 18567 16581
rect 18509 16541 18521 16575
rect 18555 16541 18567 16575
rect 18509 16535 18567 16541
rect 10778 16464 10784 16516
rect 10836 16504 10842 16516
rect 13722 16504 13728 16516
rect 10836 16476 13728 16504
rect 10836 16464 10842 16476
rect 13722 16464 13728 16476
rect 13780 16464 13786 16516
rect 17972 16504 18000 16535
rect 18138 16504 18144 16516
rect 17972 16476 18144 16504
rect 18138 16464 18144 16476
rect 18196 16504 18202 16516
rect 18524 16504 18552 16535
rect 18196 16476 18552 16504
rect 18196 16464 18202 16476
rect 12618 16396 12624 16448
rect 12676 16436 12682 16448
rect 12897 16439 12955 16445
rect 12897 16436 12909 16439
rect 12676 16408 12909 16436
rect 12676 16396 12682 16408
rect 12897 16405 12909 16408
rect 12943 16405 12955 16439
rect 13354 16436 13360 16448
rect 13315 16408 13360 16436
rect 12897 16399 12955 16405
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 15654 16396 15660 16448
rect 15712 16436 15718 16448
rect 15749 16439 15807 16445
rect 15749 16436 15761 16439
rect 15712 16408 15761 16436
rect 15712 16396 15718 16408
rect 15749 16405 15761 16408
rect 15795 16405 15807 16439
rect 16206 16436 16212 16448
rect 16167 16408 16212 16436
rect 15749 16399 15807 16405
rect 16206 16396 16212 16408
rect 16264 16396 16270 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 5905 16235 5963 16241
rect 5905 16201 5917 16235
rect 5951 16232 5963 16235
rect 6178 16232 6184 16244
rect 5951 16204 6184 16232
rect 5951 16201 5963 16204
rect 5905 16195 5963 16201
rect 6178 16192 6184 16204
rect 6236 16192 6242 16244
rect 8478 16232 8484 16244
rect 8439 16204 8484 16232
rect 8478 16192 8484 16204
rect 8536 16192 8542 16244
rect 10226 16192 10232 16244
rect 10284 16232 10290 16244
rect 10321 16235 10379 16241
rect 10321 16232 10333 16235
rect 10284 16204 10333 16232
rect 10284 16192 10290 16204
rect 10321 16201 10333 16204
rect 10367 16201 10379 16235
rect 10321 16195 10379 16201
rect 7926 16124 7932 16176
rect 7984 16164 7990 16176
rect 9953 16167 10011 16173
rect 9953 16164 9965 16167
rect 7984 16136 9965 16164
rect 7984 16124 7990 16136
rect 9953 16133 9965 16136
rect 9999 16164 10011 16167
rect 10134 16164 10140 16176
rect 9999 16136 10140 16164
rect 9999 16133 10011 16136
rect 9953 16127 10011 16133
rect 10134 16124 10140 16136
rect 10192 16124 10198 16176
rect 10336 16164 10364 16195
rect 13354 16192 13360 16244
rect 13412 16232 13418 16244
rect 15151 16235 15209 16241
rect 15151 16232 15163 16235
rect 13412 16204 15163 16232
rect 13412 16192 13418 16204
rect 15151 16201 15163 16204
rect 15197 16201 15209 16235
rect 15562 16232 15568 16244
rect 15523 16204 15568 16232
rect 15151 16195 15209 16201
rect 15562 16192 15568 16204
rect 15620 16192 15626 16244
rect 17034 16232 17040 16244
rect 16995 16204 17040 16232
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 17310 16232 17316 16244
rect 17271 16204 17316 16232
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 17865 16235 17923 16241
rect 17865 16201 17877 16235
rect 17911 16232 17923 16235
rect 18046 16232 18052 16244
rect 17911 16204 18052 16232
rect 17911 16201 17923 16204
rect 17865 16195 17923 16201
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 10336 16136 10456 16164
rect 5258 16028 5264 16040
rect 5219 16000 5264 16028
rect 5258 15988 5264 16000
rect 5316 15988 5322 16040
rect 5721 16031 5779 16037
rect 5721 16028 5733 16031
rect 5644 16000 5733 16028
rect 5644 15904 5672 16000
rect 5721 15997 5733 16000
rect 5767 15997 5779 16031
rect 5721 15991 5779 15997
rect 7285 16031 7343 16037
rect 7285 15997 7297 16031
rect 7331 15997 7343 16031
rect 7558 16028 7564 16040
rect 7471 16000 7564 16028
rect 7285 15991 7343 15997
rect 4246 15892 4252 15904
rect 4207 15864 4252 15892
rect 4246 15852 4252 15864
rect 4304 15852 4310 15904
rect 5626 15892 5632 15904
rect 5587 15864 5632 15892
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 6273 15895 6331 15901
rect 6273 15861 6285 15895
rect 6319 15892 6331 15895
rect 6641 15895 6699 15901
rect 6641 15892 6653 15895
rect 6319 15864 6653 15892
rect 6319 15861 6331 15864
rect 6273 15855 6331 15861
rect 6641 15861 6653 15864
rect 6687 15892 6699 15895
rect 7300 15892 7328 15991
rect 7558 15988 7564 16000
rect 7616 16028 7622 16040
rect 7616 16000 8248 16028
rect 7616 15988 7622 16000
rect 7742 15960 7748 15972
rect 7703 15932 7748 15960
rect 7742 15920 7748 15932
rect 7800 15920 7806 15972
rect 8220 15960 8248 16000
rect 8754 15988 8760 16040
rect 8812 16028 8818 16040
rect 8941 16031 8999 16037
rect 8941 16028 8953 16031
rect 8812 16000 8953 16028
rect 8812 15988 8818 16000
rect 8941 15997 8953 16000
rect 8987 15997 8999 16031
rect 8941 15991 8999 15997
rect 9030 15988 9036 16040
rect 9088 16028 9094 16040
rect 9493 16031 9551 16037
rect 9493 16028 9505 16031
rect 9088 16000 9505 16028
rect 9088 15988 9094 16000
rect 9493 15997 9505 16000
rect 9539 16028 9551 16031
rect 10428 16028 10456 16136
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16096 12587 16099
rect 13372 16096 13400 16192
rect 14182 16124 14188 16176
rect 14240 16164 14246 16176
rect 14461 16167 14519 16173
rect 14461 16164 14473 16167
rect 14240 16136 14473 16164
rect 14240 16124 14246 16136
rect 14461 16133 14473 16136
rect 14507 16133 14519 16167
rect 14461 16127 14519 16133
rect 15286 16124 15292 16176
rect 15344 16164 15350 16176
rect 15841 16167 15899 16173
rect 15841 16164 15853 16167
rect 15344 16136 15853 16164
rect 15344 16124 15350 16136
rect 15841 16133 15853 16136
rect 15887 16133 15899 16167
rect 15841 16127 15899 16133
rect 12575 16068 13400 16096
rect 12575 16065 12587 16068
rect 12529 16059 12587 16065
rect 10505 16031 10563 16037
rect 10505 16028 10517 16031
rect 9539 16000 9812 16028
rect 10428 16000 10517 16028
rect 9539 15997 9551 16000
rect 9493 15991 9551 15997
rect 9048 15960 9076 15988
rect 9674 15960 9680 15972
rect 8220 15932 9076 15960
rect 9635 15932 9680 15960
rect 9674 15920 9680 15932
rect 9732 15920 9738 15972
rect 9784 15960 9812 16000
rect 10505 15997 10517 16000
rect 10551 15997 10563 16031
rect 10505 15991 10563 15997
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 16028 11115 16031
rect 11517 16031 11575 16037
rect 11517 16028 11529 16031
rect 11103 16000 11529 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 11517 15997 11529 16000
rect 11563 15997 11575 16031
rect 11517 15991 11575 15997
rect 10134 15960 10140 15972
rect 9784 15932 10140 15960
rect 10134 15920 10140 15932
rect 10192 15960 10198 15972
rect 11072 15960 11100 15991
rect 13906 15988 13912 16040
rect 13964 16028 13970 16040
rect 14068 16031 14126 16037
rect 14068 16028 14080 16031
rect 13964 16000 14080 16028
rect 13964 15988 13970 16000
rect 14068 15997 14080 16000
rect 14114 16028 14126 16031
rect 14200 16028 14228 16124
rect 18138 16096 18144 16108
rect 18099 16068 18144 16096
rect 18138 16056 18144 16068
rect 18196 16056 18202 16108
rect 14114 16000 14228 16028
rect 15080 16031 15138 16037
rect 14114 15997 14126 16000
rect 14068 15991 14126 15997
rect 15080 15997 15092 16031
rect 15126 16028 15138 16031
rect 15562 16028 15568 16040
rect 15126 16000 15568 16028
rect 15126 15997 15138 16000
rect 15080 15991 15138 15997
rect 15562 15988 15568 16000
rect 15620 15988 15626 16040
rect 15654 15988 15660 16040
rect 15712 16028 15718 16040
rect 16117 16031 16175 16037
rect 16117 16028 16129 16031
rect 15712 16000 16129 16028
rect 15712 15988 15718 16000
rect 16117 15997 16129 16000
rect 16163 15997 16175 16031
rect 19705 16031 19763 16037
rect 19705 16028 19717 16031
rect 16117 15991 16175 15997
rect 19076 16000 19717 16028
rect 10192 15932 11100 15960
rect 10192 15920 10198 15932
rect 12618 15920 12624 15972
rect 12676 15960 12682 15972
rect 13170 15960 13176 15972
rect 12676 15932 12721 15960
rect 13131 15932 13176 15960
rect 12676 15920 12682 15932
rect 13170 15920 13176 15932
rect 13228 15920 13234 15972
rect 16206 15920 16212 15972
rect 16264 15960 16270 15972
rect 16438 15963 16496 15969
rect 16438 15960 16450 15963
rect 16264 15932 16450 15960
rect 16264 15920 16270 15932
rect 16438 15929 16450 15932
rect 16484 15929 16496 15963
rect 16438 15923 16496 15929
rect 18138 15920 18144 15972
rect 18196 15960 18202 15972
rect 18233 15963 18291 15969
rect 18233 15960 18245 15963
rect 18196 15932 18245 15960
rect 18196 15920 18202 15932
rect 18233 15929 18245 15932
rect 18279 15929 18291 15963
rect 18233 15923 18291 15929
rect 18785 15963 18843 15969
rect 18785 15929 18797 15963
rect 18831 15960 18843 15963
rect 18874 15960 18880 15972
rect 18831 15932 18880 15960
rect 18831 15929 18843 15932
rect 18785 15923 18843 15929
rect 18874 15920 18880 15932
rect 18932 15920 18938 15972
rect 19076 15904 19104 16000
rect 19705 15997 19717 16000
rect 19751 15997 19763 16031
rect 19705 15991 19763 15997
rect 19150 15920 19156 15972
rect 19208 15960 19214 15972
rect 19613 15963 19671 15969
rect 19613 15960 19625 15963
rect 19208 15932 19625 15960
rect 19208 15920 19214 15932
rect 19613 15929 19625 15932
rect 19659 15929 19671 15963
rect 19613 15923 19671 15929
rect 7926 15892 7932 15904
rect 6687 15864 7932 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 7926 15852 7932 15864
rect 7984 15892 7990 15904
rect 8021 15895 8079 15901
rect 8021 15892 8033 15895
rect 7984 15864 8033 15892
rect 7984 15852 7990 15864
rect 8021 15861 8033 15864
rect 8067 15861 8079 15895
rect 8754 15892 8760 15904
rect 8715 15864 8760 15892
rect 8021 15855 8079 15861
rect 8754 15852 8760 15864
rect 8812 15852 8818 15904
rect 10778 15892 10784 15904
rect 10739 15864 10784 15892
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 11977 15895 12035 15901
rect 11977 15861 11989 15895
rect 12023 15892 12035 15895
rect 12342 15892 12348 15904
rect 12023 15864 12348 15892
rect 12023 15861 12035 15864
rect 11977 15855 12035 15861
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 13446 15892 13452 15904
rect 13407 15864 13452 15892
rect 13446 15852 13452 15864
rect 13504 15852 13510 15904
rect 13538 15852 13544 15904
rect 13596 15892 13602 15904
rect 14139 15895 14197 15901
rect 14139 15892 14151 15895
rect 13596 15864 14151 15892
rect 13596 15852 13602 15864
rect 14139 15861 14151 15864
rect 14185 15861 14197 15895
rect 19058 15892 19064 15904
rect 19019 15864 19064 15892
rect 14139 15855 14197 15861
rect 19058 15852 19064 15864
rect 19116 15852 19122 15904
rect 19426 15892 19432 15904
rect 19387 15864 19432 15892
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 6365 15691 6423 15697
rect 6365 15688 6377 15691
rect 5684 15660 6377 15688
rect 5684 15648 5690 15660
rect 6365 15657 6377 15660
rect 6411 15657 6423 15691
rect 7098 15688 7104 15700
rect 7011 15660 7104 15688
rect 6365 15651 6423 15657
rect 7098 15648 7104 15660
rect 7156 15688 7162 15700
rect 7558 15688 7564 15700
rect 7156 15660 7564 15688
rect 7156 15648 7162 15660
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 9030 15688 9036 15700
rect 8991 15660 9036 15688
rect 9030 15648 9036 15660
rect 9088 15648 9094 15700
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9732 15660 9873 15688
rect 9732 15648 9738 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 9861 15651 9919 15657
rect 10413 15691 10471 15697
rect 10413 15657 10425 15691
rect 10459 15688 10471 15691
rect 10686 15688 10692 15700
rect 10459 15660 10692 15688
rect 10459 15657 10471 15660
rect 10413 15651 10471 15657
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 11701 15691 11759 15697
rect 11701 15657 11713 15691
rect 11747 15688 11759 15691
rect 11974 15688 11980 15700
rect 11747 15660 11980 15688
rect 11747 15657 11759 15660
rect 11701 15651 11759 15657
rect 11974 15648 11980 15660
rect 12032 15648 12038 15700
rect 13265 15691 13323 15697
rect 13265 15657 13277 15691
rect 13311 15688 13323 15691
rect 13538 15688 13544 15700
rect 13311 15660 13544 15688
rect 13311 15657 13323 15660
rect 13265 15651 13323 15657
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 16482 15688 16488 15700
rect 16443 15660 16488 15688
rect 16482 15648 16488 15660
rect 16540 15648 16546 15700
rect 16666 15648 16672 15700
rect 16724 15688 16730 15700
rect 16761 15691 16819 15697
rect 16761 15688 16773 15691
rect 16724 15660 16773 15688
rect 16724 15648 16730 15660
rect 16761 15657 16773 15660
rect 16807 15657 16819 15691
rect 16761 15651 16819 15657
rect 17954 15648 17960 15700
rect 18012 15648 18018 15700
rect 18322 15688 18328 15700
rect 18283 15660 18328 15688
rect 18322 15648 18328 15660
rect 18380 15648 18386 15700
rect 18782 15688 18788 15700
rect 18743 15660 18788 15688
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 7834 15629 7840 15632
rect 7831 15620 7840 15629
rect 7795 15592 7840 15620
rect 7831 15583 7840 15592
rect 7834 15580 7840 15583
rect 7892 15580 7898 15632
rect 10781 15623 10839 15629
rect 10781 15620 10793 15623
rect 8404 15592 10793 15620
rect 8404 15564 8432 15592
rect 10781 15589 10793 15592
rect 10827 15620 10839 15623
rect 10870 15620 10876 15632
rect 10827 15592 10876 15620
rect 10827 15589 10839 15592
rect 10781 15583 10839 15589
rect 10870 15580 10876 15592
rect 10928 15580 10934 15632
rect 11330 15620 11336 15632
rect 11291 15592 11336 15620
rect 11330 15580 11336 15592
rect 11388 15580 11394 15632
rect 12342 15620 12348 15632
rect 12303 15592 12348 15620
rect 12342 15580 12348 15592
rect 12400 15580 12406 15632
rect 15927 15623 15985 15629
rect 15927 15589 15939 15623
rect 15973 15620 15985 15623
rect 16206 15620 16212 15632
rect 15973 15592 16212 15620
rect 15973 15589 15985 15592
rect 15927 15583 15985 15589
rect 16206 15580 16212 15592
rect 16264 15580 16270 15632
rect 17034 15580 17040 15632
rect 17092 15620 17098 15632
rect 17494 15620 17500 15632
rect 17092 15592 17500 15620
rect 17092 15580 17098 15592
rect 17494 15580 17500 15592
rect 17552 15580 17558 15632
rect 17972 15620 18000 15648
rect 18966 15620 18972 15632
rect 17972 15592 18972 15620
rect 18966 15580 18972 15592
rect 19024 15580 19030 15632
rect 19061 15623 19119 15629
rect 19061 15589 19073 15623
rect 19107 15620 19119 15623
rect 19150 15620 19156 15632
rect 19107 15592 19156 15620
rect 19107 15589 19119 15592
rect 19061 15583 19119 15589
rect 19150 15580 19156 15592
rect 19208 15580 19214 15632
rect 5905 15555 5963 15561
rect 5905 15521 5917 15555
rect 5951 15552 5963 15555
rect 5994 15552 6000 15564
rect 5951 15524 6000 15552
rect 5951 15521 5963 15524
rect 5905 15515 5963 15521
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 6181 15555 6239 15561
rect 6181 15521 6193 15555
rect 6227 15521 6239 15555
rect 8386 15552 8392 15564
rect 8299 15524 8392 15552
rect 6181 15515 6239 15521
rect 5442 15444 5448 15496
rect 5500 15484 5506 15496
rect 6196 15484 6224 15515
rect 8386 15512 8392 15524
rect 8444 15512 8450 15564
rect 13722 15512 13728 15564
rect 13780 15561 13786 15564
rect 13780 15555 13818 15561
rect 13806 15521 13818 15555
rect 13780 15515 13818 15521
rect 13780 15512 13786 15515
rect 5500 15456 6224 15484
rect 5500 15444 5506 15456
rect 7006 15444 7012 15496
rect 7064 15484 7070 15496
rect 7469 15487 7527 15493
rect 7469 15484 7481 15487
rect 7064 15456 7481 15484
rect 7064 15444 7070 15456
rect 7469 15453 7481 15456
rect 7515 15484 7527 15487
rect 8202 15484 8208 15496
rect 7515 15456 8208 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 10686 15484 10692 15496
rect 10647 15456 10692 15484
rect 10686 15444 10692 15456
rect 10744 15444 10750 15496
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15484 12127 15487
rect 12253 15487 12311 15493
rect 12253 15484 12265 15487
rect 12115 15456 12265 15484
rect 12115 15453 12127 15456
rect 12069 15447 12127 15453
rect 12253 15453 12265 15456
rect 12299 15484 12311 15487
rect 13863 15487 13921 15493
rect 13863 15484 13875 15487
rect 12299 15456 13875 15484
rect 12299 15453 12311 15456
rect 12253 15447 12311 15453
rect 13863 15453 13875 15456
rect 13909 15453 13921 15487
rect 15562 15484 15568 15496
rect 15523 15456 15568 15484
rect 13863 15447 13921 15453
rect 15562 15444 15568 15456
rect 15620 15444 15626 15496
rect 16942 15444 16948 15496
rect 17000 15484 17006 15496
rect 17405 15487 17463 15493
rect 17405 15484 17417 15487
rect 17000 15456 17417 15484
rect 17000 15444 17006 15456
rect 17405 15453 17417 15456
rect 17451 15484 17463 15487
rect 17862 15484 17868 15496
rect 17451 15456 17868 15484
rect 17451 15453 17463 15456
rect 17405 15447 17463 15453
rect 17862 15444 17868 15456
rect 17920 15444 17926 15496
rect 5534 15376 5540 15428
rect 5592 15416 5598 15428
rect 5997 15419 6055 15425
rect 5997 15416 6009 15419
rect 5592 15388 6009 15416
rect 5592 15376 5598 15388
rect 5997 15385 6009 15388
rect 6043 15385 6055 15419
rect 5997 15379 6055 15385
rect 12434 15376 12440 15428
rect 12492 15416 12498 15428
rect 12805 15419 12863 15425
rect 12805 15416 12817 15419
rect 12492 15388 12817 15416
rect 12492 15376 12498 15388
rect 12805 15385 12817 15388
rect 12851 15385 12863 15419
rect 12805 15379 12863 15385
rect 17957 15419 18015 15425
rect 17957 15385 17969 15419
rect 18003 15416 18015 15419
rect 18874 15416 18880 15428
rect 18003 15388 18880 15416
rect 18003 15385 18015 15388
rect 17957 15379 18015 15385
rect 18874 15376 18880 15388
rect 18932 15376 18938 15428
rect 19518 15416 19524 15428
rect 19479 15388 19524 15416
rect 19518 15376 19524 15388
rect 19576 15376 19582 15428
rect 15105 15351 15163 15357
rect 15105 15317 15117 15351
rect 15151 15348 15163 15351
rect 15286 15348 15292 15360
rect 15151 15320 15292 15348
rect 15151 15317 15163 15320
rect 15105 15311 15163 15317
rect 15286 15308 15292 15320
rect 15344 15308 15350 15360
rect 19978 15348 19984 15360
rect 19939 15320 19984 15348
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 7285 15147 7343 15153
rect 7285 15113 7297 15147
rect 7331 15144 7343 15147
rect 7834 15144 7840 15156
rect 7331 15116 7840 15144
rect 7331 15113 7343 15116
rect 7285 15107 7343 15113
rect 7834 15104 7840 15116
rect 7892 15104 7898 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8941 15147 8999 15153
rect 8941 15144 8953 15147
rect 8352 15116 8953 15144
rect 8352 15104 8358 15116
rect 8941 15113 8953 15116
rect 8987 15113 8999 15147
rect 10502 15144 10508 15156
rect 10463 15116 10508 15144
rect 8941 15107 8999 15113
rect 10502 15104 10508 15116
rect 10560 15104 10566 15156
rect 11238 15144 11244 15156
rect 11199 15116 11244 15144
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 13722 15144 13728 15156
rect 13683 15116 13728 15144
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 14826 15144 14832 15156
rect 14787 15116 14832 15144
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 15289 15147 15347 15153
rect 15289 15113 15301 15147
rect 15335 15144 15347 15147
rect 16206 15144 16212 15156
rect 15335 15116 16212 15144
rect 15335 15113 15347 15116
rect 15289 15107 15347 15113
rect 16206 15104 16212 15116
rect 16264 15104 16270 15156
rect 17494 15144 17500 15156
rect 17455 15116 17500 15144
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18233 15147 18291 15153
rect 18233 15144 18245 15147
rect 18012 15116 18245 15144
rect 18012 15104 18018 15116
rect 18233 15113 18245 15116
rect 18279 15113 18291 15147
rect 18233 15107 18291 15113
rect 18969 15147 19027 15153
rect 18969 15113 18981 15147
rect 19015 15144 19027 15147
rect 19150 15144 19156 15156
rect 19015 15116 19156 15144
rect 19015 15113 19027 15116
rect 18969 15107 19027 15113
rect 19150 15104 19156 15116
rect 19208 15104 19214 15156
rect 19978 15104 19984 15156
rect 20036 15144 20042 15156
rect 21131 15147 21189 15153
rect 21131 15144 21143 15147
rect 20036 15116 21143 15144
rect 20036 15104 20042 15116
rect 21131 15113 21143 15116
rect 21177 15113 21189 15147
rect 21131 15107 21189 15113
rect 5905 15079 5963 15085
rect 5905 15045 5917 15079
rect 5951 15076 5963 15079
rect 7098 15076 7104 15088
rect 5951 15048 7104 15076
rect 5951 15045 5963 15048
rect 5905 15039 5963 15045
rect 7098 15036 7104 15048
rect 7156 15036 7162 15088
rect 7852 15076 7880 15104
rect 9401 15079 9459 15085
rect 9401 15076 9413 15079
rect 7852 15048 9413 15076
rect 9401 15045 9413 15048
rect 9447 15076 9459 15079
rect 10226 15076 10232 15088
rect 9447 15048 10232 15076
rect 9447 15045 9459 15048
rect 9401 15039 9459 15045
rect 10226 15036 10232 15048
rect 10284 15076 10290 15088
rect 11054 15076 11060 15088
rect 10284 15048 11060 15076
rect 10284 15036 10290 15048
rect 11054 15036 11060 15048
rect 11112 15036 11118 15088
rect 11146 15036 11152 15088
rect 11204 15076 11210 15088
rect 11517 15079 11575 15085
rect 11517 15076 11529 15079
rect 11204 15048 11529 15076
rect 11204 15036 11210 15048
rect 11517 15045 11529 15048
rect 11563 15045 11575 15079
rect 11517 15039 11575 15045
rect 12434 15036 12440 15088
rect 12492 15076 12498 15088
rect 13170 15076 13176 15088
rect 12492 15048 13176 15076
rect 12492 15036 12498 15048
rect 13170 15036 13176 15048
rect 13228 15076 13234 15088
rect 13357 15079 13415 15085
rect 13357 15076 13369 15079
rect 13228 15048 13369 15076
rect 13228 15036 13234 15048
rect 13357 15045 13369 15048
rect 13403 15045 13415 15079
rect 19996 15076 20024 15104
rect 13357 15039 13415 15045
rect 19536 15048 20024 15076
rect 5534 14968 5540 15020
rect 5592 15008 5598 15020
rect 6181 15011 6239 15017
rect 6181 15008 6193 15011
rect 5592 14980 6193 15008
rect 5592 14968 5598 14980
rect 6181 14977 6193 14980
rect 6227 14977 6239 15011
rect 6181 14971 6239 14977
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 15008 7435 15011
rect 7742 15008 7748 15020
rect 7423 14980 7748 15008
rect 7423 14977 7435 14980
rect 7377 14971 7435 14977
rect 7742 14968 7748 14980
rect 7800 15008 7806 15020
rect 8573 15011 8631 15017
rect 8573 15008 8585 15011
rect 7800 14980 8585 15008
rect 7800 14968 7806 14980
rect 8573 14977 8585 14980
rect 8619 14977 8631 15011
rect 9582 15008 9588 15020
rect 9543 14980 9588 15008
rect 8573 14971 8631 14977
rect 9582 14968 9588 14980
rect 9640 14968 9646 15020
rect 12161 15011 12219 15017
rect 12161 15008 12173 15011
rect 11072 14980 12173 15008
rect 5721 14943 5779 14949
rect 5721 14909 5733 14943
rect 5767 14940 5779 14943
rect 11072 14940 11100 14980
rect 12161 14977 12173 14980
rect 12207 15008 12219 15011
rect 12342 15008 12348 15020
rect 12207 14980 12348 15008
rect 12207 14977 12219 14980
rect 12161 14971 12219 14977
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 12805 15011 12863 15017
rect 12805 14977 12817 15011
rect 12851 15008 12863 15011
rect 13538 15008 13544 15020
rect 12851 14980 13544 15008
rect 12851 14977 12863 14980
rect 12805 14971 12863 14977
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 19536 15017 19564 15048
rect 19521 15011 19579 15017
rect 19521 14977 19533 15011
rect 19567 14977 19579 15011
rect 19978 15008 19984 15020
rect 19939 14980 19984 15008
rect 19521 14971 19579 14977
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 11330 14940 11336 14952
rect 5767 14912 6684 14940
rect 5767 14909 5779 14912
rect 5721 14903 5779 14909
rect 6656 14816 6684 14912
rect 8312 14912 11100 14940
rect 11291 14912 11336 14940
rect 7739 14875 7797 14881
rect 7739 14841 7751 14875
rect 7785 14872 7797 14875
rect 7834 14872 7840 14884
rect 7785 14844 7840 14872
rect 7785 14841 7797 14844
rect 7739 14835 7797 14841
rect 7834 14832 7840 14844
rect 7892 14832 7898 14884
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 5537 14807 5595 14813
rect 5537 14804 5549 14807
rect 5500 14776 5549 14804
rect 5500 14764 5506 14776
rect 5537 14773 5549 14776
rect 5583 14773 5595 14807
rect 6638 14804 6644 14816
rect 6599 14776 6644 14804
rect 5537 14767 5595 14773
rect 6638 14764 6644 14776
rect 6696 14764 6702 14816
rect 7558 14764 7564 14816
rect 7616 14804 7622 14816
rect 8312 14813 8340 14912
rect 11330 14900 11336 14912
rect 11388 14940 11394 14952
rect 11793 14943 11851 14949
rect 11793 14940 11805 14943
rect 11388 14912 11805 14940
rect 11388 14900 11394 14912
rect 11793 14909 11805 14912
rect 11839 14909 11851 14943
rect 11793 14903 11851 14909
rect 14344 14943 14402 14949
rect 14344 14909 14356 14943
rect 14390 14940 14402 14943
rect 14826 14940 14832 14952
rect 14390 14912 14832 14940
rect 14390 14909 14402 14912
rect 14344 14903 14402 14909
rect 14826 14900 14832 14912
rect 14884 14900 14890 14952
rect 15470 14940 15476 14952
rect 15431 14912 15476 14940
rect 15470 14900 15476 14912
rect 15528 14900 15534 14952
rect 15838 14940 15844 14952
rect 15799 14912 15844 14940
rect 15838 14900 15844 14912
rect 15896 14900 15902 14952
rect 16206 14940 16212 14952
rect 16167 14912 16212 14940
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 16761 14943 16819 14949
rect 16761 14909 16773 14943
rect 16807 14940 16819 14943
rect 16807 14912 17264 14940
rect 16807 14909 16819 14912
rect 16761 14903 16819 14909
rect 9926 14875 9984 14881
rect 9926 14841 9938 14875
rect 9972 14872 9984 14875
rect 10226 14872 10232 14884
rect 9972 14844 10232 14872
rect 9972 14841 9984 14844
rect 9926 14835 9984 14841
rect 10226 14832 10232 14844
rect 10284 14832 10290 14884
rect 10870 14872 10876 14884
rect 10783 14844 10876 14872
rect 10870 14832 10876 14844
rect 10928 14872 10934 14884
rect 12897 14875 12955 14881
rect 10928 14844 12756 14872
rect 10928 14832 10934 14844
rect 12728 14816 12756 14844
rect 12897 14841 12909 14875
rect 12943 14841 12955 14875
rect 12897 14835 12955 14841
rect 8297 14807 8355 14813
rect 8297 14804 8309 14807
rect 7616 14776 8309 14804
rect 7616 14764 7622 14776
rect 8297 14773 8309 14776
rect 8343 14773 8355 14807
rect 12710 14804 12716 14816
rect 12623 14776 12716 14804
rect 8297 14767 8355 14773
rect 12710 14764 12716 14776
rect 12768 14804 12774 14816
rect 12912 14804 12940 14835
rect 12768 14776 12940 14804
rect 12768 14764 12774 14776
rect 14090 14764 14096 14816
rect 14148 14804 14154 14816
rect 14415 14807 14473 14813
rect 14415 14804 14427 14807
rect 14148 14776 14427 14804
rect 14148 14764 14154 14776
rect 14415 14773 14427 14776
rect 14461 14773 14473 14807
rect 15654 14804 15660 14816
rect 15615 14776 15660 14804
rect 14415 14767 14473 14773
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 17236 14813 17264 14912
rect 20714 14900 20720 14952
rect 20772 14940 20778 14952
rect 21028 14943 21086 14949
rect 21028 14940 21040 14943
rect 20772 14912 21040 14940
rect 20772 14900 20778 14912
rect 21028 14909 21040 14912
rect 21074 14940 21086 14943
rect 21453 14943 21511 14949
rect 21453 14940 21465 14943
rect 21074 14912 21465 14940
rect 21074 14909 21086 14912
rect 21028 14903 21086 14909
rect 21453 14909 21465 14912
rect 21499 14909 21511 14943
rect 21453 14903 21511 14909
rect 23566 14900 23572 14952
rect 23624 14940 23630 14952
rect 23696 14943 23754 14949
rect 23696 14940 23708 14943
rect 23624 14912 23708 14940
rect 23624 14900 23630 14912
rect 23696 14909 23708 14912
rect 23742 14940 23754 14943
rect 24121 14943 24179 14949
rect 24121 14940 24133 14943
rect 23742 14912 24133 14940
rect 23742 14909 23754 14912
rect 23696 14903 23754 14909
rect 24121 14909 24133 14912
rect 24167 14909 24179 14943
rect 24121 14903 24179 14909
rect 19058 14832 19064 14884
rect 19116 14872 19122 14884
rect 19337 14875 19395 14881
rect 19337 14872 19349 14875
rect 19116 14844 19349 14872
rect 19116 14832 19122 14844
rect 19337 14841 19349 14844
rect 19383 14872 19395 14875
rect 19613 14875 19671 14881
rect 19613 14872 19625 14875
rect 19383 14844 19625 14872
rect 19383 14841 19395 14844
rect 19337 14835 19395 14841
rect 19613 14841 19625 14844
rect 19659 14872 19671 14875
rect 21174 14872 21180 14884
rect 19659 14844 21180 14872
rect 19659 14841 19671 14844
rect 19613 14835 19671 14841
rect 21174 14832 21180 14844
rect 21232 14832 21238 14884
rect 23799 14875 23857 14881
rect 23799 14841 23811 14875
rect 23845 14872 23857 14875
rect 24210 14872 24216 14884
rect 23845 14844 24216 14872
rect 23845 14841 23857 14844
rect 23799 14835 23857 14841
rect 24210 14832 24216 14844
rect 24268 14832 24274 14884
rect 17221 14807 17279 14813
rect 17221 14773 17233 14807
rect 17267 14804 17279 14807
rect 17586 14804 17592 14816
rect 17267 14776 17592 14804
rect 17267 14773 17279 14776
rect 17221 14767 17279 14773
rect 17586 14764 17592 14776
rect 17644 14764 17650 14816
rect 18414 14804 18420 14816
rect 18375 14776 18420 14804
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 7469 14603 7527 14609
rect 7469 14569 7481 14603
rect 7515 14600 7527 14603
rect 7834 14600 7840 14612
rect 7515 14572 7840 14600
rect 7515 14569 7527 14572
rect 7469 14563 7527 14569
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 10686 14560 10692 14612
rect 10744 14600 10750 14612
rect 10781 14603 10839 14609
rect 10781 14600 10793 14603
rect 10744 14572 10793 14600
rect 10744 14560 10750 14572
rect 10781 14569 10793 14572
rect 10827 14569 10839 14603
rect 12710 14600 12716 14612
rect 12671 14572 12716 14600
rect 10781 14563 10839 14569
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 15519 14603 15577 14609
rect 15519 14569 15531 14603
rect 15565 14600 15577 14603
rect 15746 14600 15752 14612
rect 15565 14572 15752 14600
rect 15565 14569 15577 14572
rect 15519 14563 15577 14569
rect 15746 14560 15752 14572
rect 15804 14560 15810 14612
rect 18966 14600 18972 14612
rect 18927 14572 18972 14600
rect 18966 14560 18972 14572
rect 19024 14560 19030 14612
rect 19150 14560 19156 14612
rect 19208 14600 19214 14612
rect 19208 14572 19472 14600
rect 19208 14560 19214 14572
rect 7006 14532 7012 14544
rect 6967 14504 7012 14532
rect 7006 14492 7012 14504
rect 7064 14492 7070 14544
rect 8021 14535 8079 14541
rect 8021 14501 8033 14535
rect 8067 14532 8079 14535
rect 8386 14532 8392 14544
rect 8067 14504 8392 14532
rect 8067 14501 8079 14504
rect 8021 14495 8079 14501
rect 8386 14492 8392 14504
rect 8444 14492 8450 14544
rect 9953 14535 10011 14541
rect 9953 14501 9965 14535
rect 9999 14532 10011 14535
rect 10704 14532 10732 14560
rect 9999 14504 10732 14532
rect 9999 14501 10011 14504
rect 9953 14495 10011 14501
rect 11054 14492 11060 14544
rect 11112 14532 11118 14544
rect 11698 14541 11704 14544
rect 11695 14532 11704 14541
rect 11112 14504 11704 14532
rect 11112 14492 11118 14504
rect 11695 14495 11704 14504
rect 11698 14492 11704 14495
rect 11756 14492 11762 14544
rect 13446 14541 13452 14544
rect 13443 14532 13452 14541
rect 13407 14504 13452 14532
rect 13443 14495 13452 14504
rect 13446 14492 13452 14495
rect 13504 14492 13510 14544
rect 18414 14492 18420 14544
rect 18472 14532 18478 14544
rect 19334 14532 19340 14544
rect 18472 14504 19340 14532
rect 18472 14492 18478 14504
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 19444 14541 19472 14572
rect 19429 14535 19487 14541
rect 19429 14501 19441 14535
rect 19475 14501 19487 14535
rect 19978 14532 19984 14544
rect 19939 14504 19984 14532
rect 19429 14495 19487 14501
rect 19978 14492 19984 14504
rect 20036 14492 20042 14544
rect 21085 14535 21143 14541
rect 21085 14501 21097 14535
rect 21131 14532 21143 14535
rect 21174 14532 21180 14544
rect 21131 14504 21180 14532
rect 21131 14501 21143 14504
rect 21085 14495 21143 14501
rect 21174 14492 21180 14504
rect 21232 14492 21238 14544
rect 5261 14467 5319 14473
rect 5261 14433 5273 14467
rect 5307 14464 5319 14467
rect 5350 14464 5356 14476
rect 5307 14436 5356 14464
rect 5307 14433 5319 14436
rect 5261 14427 5319 14433
rect 5350 14424 5356 14436
rect 5408 14424 5414 14476
rect 6546 14464 6552 14476
rect 6507 14436 6552 14464
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 6825 14467 6883 14473
rect 6825 14433 6837 14467
rect 6871 14464 6883 14467
rect 7098 14464 7104 14476
rect 6871 14436 7104 14464
rect 6871 14433 6883 14436
rect 6825 14427 6883 14433
rect 7098 14424 7104 14436
rect 7156 14424 7162 14476
rect 13078 14464 13084 14476
rect 13039 14436 13084 14464
rect 13078 14424 13084 14436
rect 13136 14424 13142 14476
rect 14642 14424 14648 14476
rect 14700 14464 14706 14476
rect 15416 14467 15474 14473
rect 15416 14464 15428 14467
rect 14700 14436 15428 14464
rect 14700 14424 14706 14436
rect 15416 14433 15428 14436
rect 15462 14433 15474 14467
rect 16574 14464 16580 14476
rect 16535 14436 16580 14464
rect 15416 14427 15474 14433
rect 16574 14424 16580 14436
rect 16632 14424 16638 14476
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 16853 14467 16911 14473
rect 16853 14464 16865 14467
rect 16724 14436 16865 14464
rect 16724 14424 16730 14436
rect 16853 14433 16865 14436
rect 16899 14433 16911 14467
rect 16853 14427 16911 14433
rect 17034 14424 17040 14476
rect 17092 14464 17098 14476
rect 17221 14467 17279 14473
rect 17221 14464 17233 14467
rect 17092 14436 17233 14464
rect 17092 14424 17098 14436
rect 17221 14433 17233 14436
rect 17267 14433 17279 14467
rect 17586 14464 17592 14476
rect 17547 14436 17592 14464
rect 17221 14427 17279 14433
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 7466 14356 7472 14408
rect 7524 14396 7530 14408
rect 7929 14399 7987 14405
rect 7929 14396 7941 14399
rect 7524 14368 7941 14396
rect 7524 14356 7530 14368
rect 7929 14365 7941 14368
rect 7975 14396 7987 14399
rect 8849 14399 8907 14405
rect 8849 14396 8861 14399
rect 7975 14368 8861 14396
rect 7975 14365 7987 14368
rect 7929 14359 7987 14365
rect 8849 14365 8861 14368
rect 8895 14365 8907 14399
rect 9858 14396 9864 14408
rect 9819 14368 9864 14396
rect 8849 14359 8907 14365
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14396 10563 14399
rect 10686 14396 10692 14408
rect 10551 14368 10692 14396
rect 10551 14365 10563 14368
rect 10505 14359 10563 14365
rect 8386 14288 8392 14340
rect 8444 14328 8450 14340
rect 8481 14331 8539 14337
rect 8481 14328 8493 14331
rect 8444 14300 8493 14328
rect 8444 14288 8450 14300
rect 8481 14297 8493 14300
rect 8527 14328 8539 14331
rect 10520 14328 10548 14359
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14396 11391 14399
rect 11974 14396 11980 14408
rect 11379 14368 11980 14396
rect 11379 14365 11391 14368
rect 11333 14359 11391 14365
rect 11974 14356 11980 14368
rect 12032 14356 12038 14408
rect 16301 14399 16359 14405
rect 16301 14365 16313 14399
rect 16347 14396 16359 14399
rect 17604 14396 17632 14424
rect 16347 14368 17632 14396
rect 17865 14399 17923 14405
rect 16347 14365 16359 14368
rect 16301 14359 16359 14365
rect 17865 14365 17877 14399
rect 17911 14396 17923 14399
rect 17954 14396 17960 14408
rect 17911 14368 17960 14396
rect 17911 14365 17923 14368
rect 17865 14359 17923 14365
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 20990 14396 20996 14408
rect 20951 14368 20996 14396
rect 20990 14356 20996 14368
rect 21048 14356 21054 14408
rect 21266 14396 21272 14408
rect 21227 14368 21272 14396
rect 21266 14356 21272 14368
rect 21324 14356 21330 14408
rect 8527 14300 10548 14328
rect 8527 14297 8539 14300
rect 8481 14291 8539 14297
rect 5445 14263 5503 14269
rect 5445 14229 5457 14263
rect 5491 14260 5503 14263
rect 5994 14260 6000 14272
rect 5491 14232 6000 14260
rect 5491 14229 5503 14232
rect 5445 14223 5503 14229
rect 5994 14220 6000 14232
rect 6052 14260 6058 14272
rect 6822 14260 6828 14272
rect 6052 14232 6828 14260
rect 6052 14220 6058 14232
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 9122 14220 9128 14272
rect 9180 14260 9186 14272
rect 9217 14263 9275 14269
rect 9217 14260 9229 14263
rect 9180 14232 9229 14260
rect 9180 14220 9186 14232
rect 9217 14229 9229 14232
rect 9263 14229 9275 14263
rect 11146 14260 11152 14272
rect 11107 14232 11152 14260
rect 9217 14223 9275 14229
rect 11146 14220 11152 14232
rect 11204 14220 11210 14272
rect 12250 14260 12256 14272
rect 12211 14232 12256 14260
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 14001 14263 14059 14269
rect 14001 14260 14013 14263
rect 12860 14232 14013 14260
rect 12860 14220 12866 14232
rect 14001 14229 14013 14232
rect 14047 14229 14059 14263
rect 14734 14260 14740 14272
rect 14695 14232 14740 14260
rect 14001 14223 14059 14229
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 15105 14263 15163 14269
rect 15105 14229 15117 14263
rect 15151 14260 15163 14263
rect 15470 14260 15476 14272
rect 15151 14232 15476 14260
rect 15151 14229 15163 14232
rect 15105 14223 15163 14229
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 15838 14220 15844 14272
rect 15896 14260 15902 14272
rect 15933 14263 15991 14269
rect 15933 14260 15945 14263
rect 15896 14232 15945 14260
rect 15896 14220 15902 14232
rect 15933 14229 15945 14232
rect 15979 14260 15991 14263
rect 16666 14260 16672 14272
rect 15979 14232 16672 14260
rect 15979 14229 15991 14232
rect 15933 14223 15991 14229
rect 16666 14220 16672 14232
rect 16724 14220 16730 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 4154 14056 4160 14068
rect 4115 14028 4160 14056
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 6270 14016 6276 14068
rect 6328 14056 6334 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 6328 14028 6377 14056
rect 6328 14016 6334 14028
rect 6365 14025 6377 14028
rect 6411 14056 6423 14059
rect 6546 14056 6552 14068
rect 6411 14028 6552 14056
rect 6411 14025 6423 14028
rect 6365 14019 6423 14025
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 7098 14056 7104 14068
rect 7059 14028 7104 14056
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 8665 14059 8723 14065
rect 8665 14056 8677 14059
rect 8536 14028 8677 14056
rect 8536 14016 8542 14028
rect 8665 14025 8677 14028
rect 8711 14025 8723 14059
rect 9030 14056 9036 14068
rect 8991 14028 9036 14056
rect 8665 14019 8723 14025
rect 9030 14016 9036 14028
rect 9088 14056 9094 14068
rect 9088 14028 9352 14056
rect 9088 14016 9094 14028
rect 9324 13997 9352 14028
rect 9858 14016 9864 14068
rect 9916 14056 9922 14068
rect 10229 14059 10287 14065
rect 10229 14056 10241 14059
rect 9916 14028 10241 14056
rect 9916 14016 9922 14028
rect 10229 14025 10241 14028
rect 10275 14025 10287 14059
rect 10594 14056 10600 14068
rect 10555 14028 10600 14056
rect 10229 14019 10287 14025
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 14642 14016 14648 14068
rect 14700 14056 14706 14068
rect 15013 14059 15071 14065
rect 15013 14056 15025 14059
rect 14700 14028 15025 14056
rect 14700 14016 14706 14028
rect 15013 14025 15025 14028
rect 15059 14025 15071 14059
rect 15013 14019 15071 14025
rect 16298 14016 16304 14068
rect 16356 14056 16362 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 16356 14028 17785 14056
rect 16356 14016 16362 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 17773 14019 17831 14025
rect 18969 14059 19027 14065
rect 18969 14025 18981 14059
rect 19015 14056 19027 14059
rect 19058 14056 19064 14068
rect 19015 14028 19064 14056
rect 19015 14025 19027 14028
rect 18969 14019 19027 14025
rect 9309 13991 9367 13997
rect 9309 13957 9321 13991
rect 9355 13957 9367 13991
rect 11422 13988 11428 14000
rect 11383 13960 11428 13988
rect 9309 13951 9367 13957
rect 11422 13948 11428 13960
rect 11480 13948 11486 14000
rect 14737 13991 14795 13997
rect 14737 13957 14749 13991
rect 14783 13988 14795 13991
rect 15838 13988 15844 14000
rect 14783 13960 15844 13988
rect 14783 13957 14795 13960
rect 14737 13951 14795 13957
rect 15838 13948 15844 13960
rect 15896 13948 15902 14000
rect 6362 13880 6368 13932
rect 6420 13920 6426 13932
rect 6546 13920 6552 13932
rect 6420 13892 6552 13920
rect 6420 13880 6426 13892
rect 6546 13880 6552 13892
rect 6604 13880 6610 13932
rect 7745 13923 7803 13929
rect 7745 13889 7757 13923
rect 7791 13920 7803 13923
rect 8018 13920 8024 13932
rect 7791 13892 8024 13920
rect 7791 13889 7803 13892
rect 7745 13883 7803 13889
rect 8018 13880 8024 13892
rect 8076 13880 8082 13932
rect 8386 13920 8392 13932
rect 8347 13892 8392 13920
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 9674 13920 9680 13932
rect 9635 13892 9680 13920
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 9950 13880 9956 13932
rect 10008 13920 10014 13932
rect 10873 13923 10931 13929
rect 10873 13920 10885 13923
rect 10008 13892 10885 13920
rect 10008 13880 10014 13892
rect 10873 13889 10885 13892
rect 10919 13920 10931 13923
rect 11146 13920 11152 13932
rect 10919 13892 11152 13920
rect 10919 13889 10931 13892
rect 10873 13883 10931 13889
rect 11146 13880 11152 13892
rect 11204 13880 11210 13932
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 12802 13920 12808 13932
rect 12299 13892 12808 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 12986 13920 12992 13932
rect 12947 13892 12992 13920
rect 12986 13880 12992 13892
rect 13044 13880 13050 13932
rect 13998 13880 14004 13932
rect 14056 13920 14062 13932
rect 14642 13920 14648 13932
rect 14056 13892 14648 13920
rect 14056 13880 14062 13892
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 15286 13880 15292 13932
rect 15344 13920 15350 13932
rect 16206 13920 16212 13932
rect 15344 13892 16212 13920
rect 15344 13880 15350 13892
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4433 13855 4491 13861
rect 4433 13852 4445 13855
rect 4212 13824 4445 13852
rect 4212 13812 4218 13824
rect 4433 13821 4445 13824
rect 4479 13852 4491 13855
rect 4890 13852 4896 13864
rect 4479 13824 4896 13852
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 5350 13852 5356 13864
rect 5311 13824 5356 13852
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 7558 13852 7564 13864
rect 7471 13824 7564 13852
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 9214 13852 9220 13864
rect 9175 13824 9220 13852
rect 9214 13812 9220 13824
rect 9272 13812 9278 13864
rect 9493 13855 9551 13861
rect 9493 13821 9505 13855
rect 9539 13821 9551 13855
rect 9493 13815 9551 13821
rect 4338 13784 4344 13796
rect 4299 13756 4344 13784
rect 4338 13744 4344 13756
rect 4396 13744 4402 13796
rect 7576 13784 7604 13812
rect 7837 13787 7895 13793
rect 7837 13784 7849 13787
rect 7576 13756 7849 13784
rect 7837 13753 7849 13756
rect 7883 13753 7895 13787
rect 7837 13747 7895 13753
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 9508 13784 9536 13815
rect 10594 13812 10600 13864
rect 10652 13852 10658 13864
rect 10652 13824 10732 13852
rect 10652 13812 10658 13824
rect 9180 13756 9536 13784
rect 10704 13784 10732 13824
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 15470 13852 15476 13864
rect 14792 13824 15148 13852
rect 15431 13824 15476 13852
rect 14792 13812 14798 13824
rect 10965 13787 11023 13793
rect 10965 13784 10977 13787
rect 10704 13756 10977 13784
rect 9180 13744 9186 13756
rect 10965 13753 10977 13756
rect 11011 13753 11023 13787
rect 10965 13747 11023 13753
rect 12434 13744 12440 13796
rect 12492 13784 12498 13796
rect 12713 13787 12771 13793
rect 12713 13784 12725 13787
rect 12492 13756 12725 13784
rect 12492 13744 12498 13756
rect 12713 13753 12725 13756
rect 12759 13753 12771 13787
rect 12713 13747 12771 13753
rect 12802 13744 12808 13796
rect 12860 13784 12866 13796
rect 15120 13784 15148 13824
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 15838 13852 15844 13864
rect 15799 13824 15844 13852
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 16040 13861 16068 13892
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13821 16083 13855
rect 16025 13815 16083 13821
rect 16485 13855 16543 13861
rect 16485 13821 16497 13855
rect 16531 13821 16543 13855
rect 16485 13815 16543 13821
rect 15562 13784 15568 13796
rect 12860 13756 12905 13784
rect 15120 13756 15568 13784
rect 12860 13744 12866 13756
rect 11238 13676 11244 13728
rect 11296 13716 11302 13728
rect 11698 13716 11704 13728
rect 11296 13688 11704 13716
rect 11296 13676 11302 13688
rect 11698 13676 11704 13688
rect 11756 13716 11762 13728
rect 11793 13719 11851 13725
rect 11793 13716 11805 13719
rect 11756 13688 11805 13716
rect 11756 13676 11762 13688
rect 11793 13685 11805 13688
rect 11839 13716 11851 13719
rect 13446 13716 13452 13728
rect 11839 13688 13452 13716
rect 11839 13685 11851 13688
rect 11793 13679 11851 13685
rect 13446 13676 13452 13688
rect 13504 13716 13510 13728
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 13504 13688 13645 13716
rect 13504 13676 13510 13688
rect 13633 13685 13645 13688
rect 13679 13685 13691 13719
rect 14366 13716 14372 13728
rect 14327 13688 14372 13716
rect 13633 13679 13691 13685
rect 14366 13676 14372 13688
rect 14424 13676 14430 13728
rect 15304 13725 15332 13756
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 16500 13784 16528 13815
rect 16666 13812 16672 13864
rect 16724 13852 16730 13864
rect 17313 13855 17371 13861
rect 17313 13852 17325 13855
rect 16724 13824 17325 13852
rect 16724 13812 16730 13824
rect 17313 13821 17325 13824
rect 17359 13821 17371 13855
rect 17313 13815 17371 13821
rect 16850 13784 16856 13796
rect 16500 13756 16856 13784
rect 16850 13744 16856 13756
rect 16908 13744 16914 13796
rect 17788 13784 17816 14019
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 19150 14016 19156 14068
rect 19208 14056 19214 14068
rect 19245 14059 19303 14065
rect 19245 14056 19257 14059
rect 19208 14028 19257 14056
rect 19208 14016 19214 14028
rect 19245 14025 19257 14028
rect 19291 14025 19303 14059
rect 19245 14019 19303 14025
rect 19334 14016 19340 14068
rect 19392 14056 19398 14068
rect 19613 14059 19671 14065
rect 19613 14056 19625 14059
rect 19392 14028 19625 14056
rect 19392 14016 19398 14028
rect 19613 14025 19625 14028
rect 19659 14025 19671 14059
rect 21174 14056 21180 14068
rect 21135 14028 21180 14056
rect 19613 14019 19671 14025
rect 21174 14016 21180 14028
rect 21232 14016 21238 14068
rect 19978 13880 19984 13932
rect 20036 13920 20042 13932
rect 20257 13923 20315 13929
rect 20257 13920 20269 13923
rect 20036 13892 20269 13920
rect 20036 13880 20042 13892
rect 20257 13889 20269 13892
rect 20303 13889 20315 13923
rect 20257 13883 20315 13889
rect 18046 13852 18052 13864
rect 18007 13824 18052 13852
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 20073 13855 20131 13861
rect 20073 13821 20085 13855
rect 20119 13821 20131 13855
rect 20073 13815 20131 13821
rect 18370 13787 18428 13793
rect 18370 13784 18382 13787
rect 17788 13756 18382 13784
rect 18370 13753 18382 13756
rect 18416 13784 18428 13787
rect 18874 13784 18880 13796
rect 18416 13756 18880 13784
rect 18416 13753 18428 13756
rect 18370 13747 18428 13753
rect 18874 13744 18880 13756
rect 18932 13744 18938 13796
rect 20088 13784 20116 13815
rect 20898 13812 20904 13864
rect 20956 13852 20962 13864
rect 21542 13852 21548 13864
rect 20956 13824 21001 13852
rect 21503 13824 21548 13852
rect 20956 13812 20962 13824
rect 21542 13812 21548 13824
rect 21600 13812 21606 13864
rect 20349 13787 20407 13793
rect 20349 13784 20361 13787
rect 20088 13756 20361 13784
rect 20349 13753 20361 13756
rect 20395 13784 20407 13787
rect 20714 13784 20720 13796
rect 20395 13756 20720 13784
rect 20395 13753 20407 13756
rect 20349 13747 20407 13753
rect 20714 13744 20720 13756
rect 20772 13744 20778 13796
rect 15289 13719 15347 13725
rect 15289 13685 15301 13719
rect 15335 13685 15347 13719
rect 17034 13716 17040 13728
rect 16995 13688 17040 13716
rect 15289 13679 15347 13685
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 9769 13515 9827 13521
rect 9769 13481 9781 13515
rect 9815 13512 9827 13515
rect 9858 13512 9864 13524
rect 9815 13484 9864 13512
rect 9815 13481 9827 13484
rect 9769 13475 9827 13481
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 10042 13472 10048 13524
rect 10100 13512 10106 13524
rect 10321 13515 10379 13521
rect 10321 13512 10333 13515
rect 10100 13484 10333 13512
rect 10100 13472 10106 13484
rect 10321 13481 10333 13484
rect 10367 13481 10379 13515
rect 10321 13475 10379 13481
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12492 13484 12537 13512
rect 12492 13472 12498 13484
rect 13078 13472 13084 13524
rect 13136 13512 13142 13524
rect 13541 13515 13599 13521
rect 13541 13512 13553 13515
rect 13136 13484 13553 13512
rect 13136 13472 13142 13484
rect 13541 13481 13553 13484
rect 13587 13481 13599 13515
rect 14366 13512 14372 13524
rect 14279 13484 14372 13512
rect 13541 13475 13599 13481
rect 14366 13472 14372 13484
rect 14424 13512 14430 13524
rect 15470 13512 15476 13524
rect 14424 13484 15476 13512
rect 14424 13472 14430 13484
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 19518 13472 19524 13524
rect 19576 13512 19582 13524
rect 19889 13515 19947 13521
rect 19889 13512 19901 13515
rect 19576 13484 19901 13512
rect 19576 13472 19582 13484
rect 19889 13481 19901 13484
rect 19935 13481 19947 13515
rect 19889 13475 19947 13481
rect 19978 13472 19984 13524
rect 20036 13512 20042 13524
rect 20257 13515 20315 13521
rect 20257 13512 20269 13515
rect 20036 13484 20269 13512
rect 20036 13472 20042 13484
rect 20257 13481 20269 13484
rect 20303 13481 20315 13515
rect 20257 13475 20315 13481
rect 4154 13404 4160 13456
rect 4212 13444 4218 13456
rect 11143 13447 11201 13453
rect 4212 13416 5120 13444
rect 4212 13404 4218 13416
rect 4614 13336 4620 13388
rect 4672 13376 4678 13388
rect 5092 13385 5120 13416
rect 11143 13413 11155 13447
rect 11189 13444 11201 13447
rect 11238 13444 11244 13456
rect 11189 13416 11244 13444
rect 11189 13413 11201 13416
rect 11143 13407 11201 13413
rect 11238 13404 11244 13416
rect 11296 13404 11302 13456
rect 12250 13404 12256 13456
rect 12308 13444 12314 13456
rect 12713 13447 12771 13453
rect 12713 13444 12725 13447
rect 12308 13416 12725 13444
rect 12308 13404 12314 13416
rect 12713 13413 12725 13416
rect 12759 13413 12771 13447
rect 12713 13407 12771 13413
rect 17773 13447 17831 13453
rect 17773 13413 17785 13447
rect 17819 13444 17831 13447
rect 18046 13444 18052 13456
rect 17819 13416 18052 13444
rect 17819 13413 17831 13416
rect 17773 13407 17831 13413
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 18874 13404 18880 13456
rect 18932 13453 18938 13456
rect 18932 13447 18980 13453
rect 18932 13413 18934 13447
rect 18968 13413 18980 13447
rect 18932 13407 18980 13413
rect 18932 13404 18938 13407
rect 20714 13404 20720 13456
rect 20772 13444 20778 13456
rect 20901 13447 20959 13453
rect 20901 13444 20913 13447
rect 20772 13416 20913 13444
rect 20772 13404 20778 13416
rect 20901 13413 20913 13416
rect 20947 13413 20959 13447
rect 20901 13407 20959 13413
rect 4801 13379 4859 13385
rect 4801 13376 4813 13379
rect 4672 13348 4813 13376
rect 4672 13336 4678 13348
rect 4801 13345 4813 13348
rect 4847 13345 4859 13379
rect 4801 13339 4859 13345
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13345 5135 13379
rect 7282 13376 7288 13388
rect 7243 13348 7288 13376
rect 5077 13339 5135 13345
rect 7282 13336 7288 13348
rect 7340 13376 7346 13388
rect 8573 13379 8631 13385
rect 8573 13376 8585 13379
rect 7340 13348 8585 13376
rect 7340 13336 7346 13348
rect 8573 13345 8585 13348
rect 8619 13376 8631 13379
rect 8754 13376 8760 13388
rect 8619 13348 8760 13376
rect 8619 13345 8631 13348
rect 8573 13339 8631 13345
rect 8754 13336 8760 13348
rect 8812 13336 8818 13388
rect 14185 13379 14243 13385
rect 14185 13345 14197 13379
rect 14231 13376 14243 13379
rect 14366 13376 14372 13388
rect 14231 13348 14372 13376
rect 14231 13345 14243 13348
rect 14185 13339 14243 13345
rect 14366 13336 14372 13348
rect 14424 13336 14430 13388
rect 15470 13336 15476 13388
rect 15528 13376 15534 13388
rect 16209 13379 16267 13385
rect 16209 13376 16221 13379
rect 15528 13348 16221 13376
rect 15528 13336 15534 13348
rect 16209 13345 16221 13348
rect 16255 13376 16267 13379
rect 16574 13376 16580 13388
rect 16255 13348 16580 13376
rect 16255 13345 16267 13348
rect 16209 13339 16267 13345
rect 16574 13336 16580 13348
rect 16632 13336 16638 13388
rect 16666 13336 16672 13388
rect 16724 13376 16730 13388
rect 16761 13379 16819 13385
rect 16761 13376 16773 13379
rect 16724 13348 16773 13376
rect 16724 13336 16730 13348
rect 16761 13345 16773 13348
rect 16807 13345 16819 13379
rect 16761 13339 16819 13345
rect 16850 13336 16856 13388
rect 16908 13376 16914 13388
rect 17034 13376 17040 13388
rect 16908 13348 17040 13376
rect 16908 13336 16914 13348
rect 17034 13336 17040 13348
rect 17092 13376 17098 13388
rect 17129 13379 17187 13385
rect 17129 13376 17141 13379
rect 17092 13348 17141 13376
rect 17092 13336 17098 13348
rect 17129 13345 17141 13348
rect 17175 13345 17187 13379
rect 17129 13339 17187 13345
rect 17497 13379 17555 13385
rect 17497 13345 17509 13379
rect 17543 13345 17555 13379
rect 17497 13339 17555 13345
rect 4338 13268 4344 13320
rect 4396 13308 4402 13320
rect 4893 13311 4951 13317
rect 4893 13308 4905 13311
rect 4396 13280 4905 13308
rect 4396 13268 4402 13280
rect 4893 13277 4905 13280
rect 4939 13308 4951 13311
rect 5258 13308 5264 13320
rect 4939 13280 5264 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13308 5503 13311
rect 5534 13308 5540 13320
rect 5491 13280 5540 13308
rect 5491 13277 5503 13280
rect 5445 13271 5503 13277
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 10778 13308 10784 13320
rect 10739 13280 10784 13308
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 12066 13308 12072 13320
rect 11480 13280 12072 13308
rect 11480 13268 11486 13280
rect 12066 13268 12072 13280
rect 12124 13308 12130 13320
rect 12621 13311 12679 13317
rect 12621 13308 12633 13311
rect 12124 13280 12633 13308
rect 12124 13268 12130 13280
rect 12621 13277 12633 13280
rect 12667 13277 12679 13311
rect 12621 13271 12679 13277
rect 12710 13268 12716 13320
rect 12768 13308 12774 13320
rect 12897 13311 12955 13317
rect 12897 13308 12909 13311
rect 12768 13280 12909 13308
rect 12768 13268 12774 13280
rect 12897 13277 12909 13280
rect 12943 13308 12955 13311
rect 12986 13308 12992 13320
rect 12943 13280 12992 13308
rect 12943 13277 12955 13280
rect 12897 13271 12955 13277
rect 12986 13268 12992 13280
rect 13044 13268 13050 13320
rect 13998 13268 14004 13320
rect 14056 13308 14062 13320
rect 15013 13311 15071 13317
rect 15013 13308 15025 13311
rect 14056 13280 15025 13308
rect 14056 13268 14062 13280
rect 15013 13277 15025 13280
rect 15059 13308 15071 13311
rect 15286 13308 15292 13320
rect 15059 13280 15292 13308
rect 15059 13277 15071 13280
rect 15013 13271 15071 13277
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17512 13308 17540 13339
rect 17954 13336 17960 13388
rect 18012 13376 18018 13388
rect 18601 13379 18659 13385
rect 18601 13376 18613 13379
rect 18012 13348 18613 13376
rect 18012 13336 18018 13348
rect 18601 13345 18613 13348
rect 18647 13345 18659 13379
rect 18601 13339 18659 13345
rect 19521 13379 19579 13385
rect 19521 13345 19533 13379
rect 19567 13376 19579 13379
rect 20990 13376 20996 13388
rect 19567 13348 20996 13376
rect 19567 13345 19579 13348
rect 19521 13339 19579 13345
rect 20990 13336 20996 13348
rect 21048 13336 21054 13388
rect 17000 13280 17540 13308
rect 17000 13268 17006 13280
rect 6917 13243 6975 13249
rect 6917 13209 6929 13243
rect 6963 13240 6975 13243
rect 8018 13240 8024 13252
rect 6963 13212 8024 13240
rect 6963 13209 6975 13212
rect 6917 13203 6975 13209
rect 8018 13200 8024 13212
rect 8076 13200 8082 13252
rect 8570 13200 8576 13252
rect 8628 13240 8634 13252
rect 9214 13240 9220 13252
rect 8628 13212 9220 13240
rect 8628 13200 8634 13212
rect 9214 13200 9220 13212
rect 9272 13200 9278 13252
rect 12526 13200 12532 13252
rect 12584 13240 12590 13252
rect 13909 13243 13967 13249
rect 13909 13240 13921 13243
rect 12584 13212 13921 13240
rect 12584 13200 12590 13212
rect 13909 13209 13921 13212
rect 13955 13209 13967 13243
rect 15473 13243 15531 13249
rect 15473 13240 15485 13243
rect 13909 13203 13967 13209
rect 14660 13212 15485 13240
rect 7469 13175 7527 13181
rect 7469 13141 7481 13175
rect 7515 13172 7527 13175
rect 8110 13172 8116 13184
rect 7515 13144 8116 13172
rect 7515 13141 7527 13144
rect 7469 13135 7527 13141
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 8478 13172 8484 13184
rect 8439 13144 8484 13172
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 8757 13175 8815 13181
rect 8757 13141 8769 13175
rect 8803 13172 8815 13175
rect 9122 13172 9128 13184
rect 8803 13144 9128 13172
rect 8803 13141 8815 13144
rect 8757 13135 8815 13141
rect 9122 13132 9128 13144
rect 9180 13132 9186 13184
rect 11698 13172 11704 13184
rect 11659 13144 11704 13172
rect 11698 13132 11704 13144
rect 11756 13132 11762 13184
rect 11974 13172 11980 13184
rect 11935 13144 11980 13172
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 14458 13132 14464 13184
rect 14516 13172 14522 13184
rect 14660 13181 14688 13212
rect 15473 13209 15485 13212
rect 15519 13240 15531 13243
rect 15562 13240 15568 13252
rect 15519 13212 15568 13240
rect 15519 13209 15531 13212
rect 15473 13203 15531 13209
rect 15562 13200 15568 13212
rect 15620 13200 15626 13252
rect 14645 13175 14703 13181
rect 14645 13172 14657 13175
rect 14516 13144 14657 13172
rect 14516 13132 14522 13144
rect 14645 13141 14657 13144
rect 14691 13141 14703 13175
rect 14645 13135 14703 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 4154 12928 4160 12980
rect 4212 12968 4218 12980
rect 4249 12971 4307 12977
rect 4249 12968 4261 12971
rect 4212 12940 4261 12968
rect 4212 12928 4218 12940
rect 4249 12937 4261 12940
rect 4295 12937 4307 12971
rect 4249 12931 4307 12937
rect 2409 12767 2467 12773
rect 2409 12733 2421 12767
rect 2455 12733 2467 12767
rect 2409 12727 2467 12733
rect 3421 12767 3479 12773
rect 3421 12733 3433 12767
rect 3467 12764 3479 12767
rect 4264 12764 4292 12931
rect 5258 12928 5264 12980
rect 5316 12968 5322 12980
rect 5813 12971 5871 12977
rect 5813 12968 5825 12971
rect 5316 12940 5825 12968
rect 5316 12928 5322 12940
rect 5813 12937 5825 12940
rect 5859 12937 5871 12971
rect 5813 12931 5871 12937
rect 7101 12971 7159 12977
rect 7101 12937 7113 12971
rect 7147 12968 7159 12971
rect 7282 12968 7288 12980
rect 7147 12940 7288 12968
rect 7147 12937 7159 12940
rect 7101 12931 7159 12937
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 8754 12968 8760 12980
rect 8715 12940 8760 12968
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 10134 12968 10140 12980
rect 10095 12940 10140 12968
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 11793 12971 11851 12977
rect 11793 12968 11805 12971
rect 11756 12940 11805 12968
rect 11756 12928 11762 12940
rect 11793 12937 11805 12940
rect 11839 12968 11851 12971
rect 12618 12968 12624 12980
rect 11839 12940 12624 12968
rect 11839 12937 11851 12940
rect 11793 12931 11851 12937
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 16022 12928 16028 12980
rect 16080 12968 16086 12980
rect 16574 12968 16580 12980
rect 16080 12940 16580 12968
rect 16080 12928 16086 12940
rect 16574 12928 16580 12940
rect 16632 12968 16638 12980
rect 17405 12971 17463 12977
rect 17405 12968 17417 12971
rect 16632 12940 17417 12968
rect 16632 12928 16638 12940
rect 17405 12937 17417 12940
rect 17451 12937 17463 12971
rect 17405 12931 17463 12937
rect 17954 12928 17960 12980
rect 18012 12968 18018 12980
rect 18233 12971 18291 12977
rect 18233 12968 18245 12971
rect 18012 12940 18245 12968
rect 18012 12928 18018 12940
rect 18233 12937 18245 12940
rect 18279 12937 18291 12971
rect 18233 12931 18291 12937
rect 18693 12971 18751 12977
rect 18693 12937 18705 12971
rect 18739 12968 18751 12971
rect 18782 12968 18788 12980
rect 18739 12940 18788 12968
rect 18739 12937 18751 12940
rect 18693 12931 18751 12937
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 18923 12971 18981 12977
rect 18923 12937 18935 12971
rect 18969 12968 18981 12971
rect 19242 12968 19248 12980
rect 18969 12940 19248 12968
rect 18969 12937 18981 12940
rect 18923 12931 18981 12937
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 20990 12968 20996 12980
rect 20951 12940 20996 12968
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 8478 12900 8484 12912
rect 6972 12872 8484 12900
rect 6972 12860 6978 12872
rect 4430 12764 4436 12776
rect 3467 12736 4016 12764
rect 4264 12736 4436 12764
rect 3467 12733 3479 12736
rect 3421 12727 3479 12733
rect 2424 12696 2452 12727
rect 2866 12696 2872 12708
rect 2424 12668 2872 12696
rect 2866 12656 2872 12668
rect 2924 12656 2930 12708
rect 2590 12628 2596 12640
rect 2551 12600 2596 12628
rect 2590 12588 2596 12600
rect 2648 12588 2654 12640
rect 3602 12628 3608 12640
rect 3563 12600 3608 12628
rect 3602 12588 3608 12600
rect 3660 12588 3666 12640
rect 3988 12637 4016 12736
rect 4430 12724 4436 12736
rect 4488 12764 4494 12776
rect 7760 12773 7788 12872
rect 8478 12860 8484 12872
rect 8536 12860 8542 12912
rect 8294 12832 8300 12844
rect 8255 12804 8300 12832
rect 8294 12792 8300 12804
rect 8352 12792 8358 12844
rect 9769 12835 9827 12841
rect 9769 12832 9781 12835
rect 9324 12804 9781 12832
rect 4525 12767 4583 12773
rect 4525 12764 4537 12767
rect 4488 12736 4537 12764
rect 4488 12724 4494 12736
rect 4525 12733 4537 12736
rect 4571 12764 4583 12767
rect 5445 12767 5503 12773
rect 5445 12764 5457 12767
rect 4571 12736 5457 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 5445 12733 5457 12736
rect 5491 12733 5503 12767
rect 5445 12727 5503 12733
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 8110 12764 8116 12776
rect 8067 12736 8116 12764
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 5166 12696 5172 12708
rect 5127 12668 5172 12696
rect 5166 12656 5172 12668
rect 5224 12656 5230 12708
rect 7558 12696 7564 12708
rect 7519 12668 7564 12696
rect 7558 12656 7564 12668
rect 7616 12696 7622 12708
rect 7852 12696 7880 12727
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 9030 12724 9036 12776
rect 9088 12764 9094 12776
rect 9324 12773 9352 12804
rect 9769 12801 9781 12804
rect 9815 12801 9827 12835
rect 10152 12832 10180 12928
rect 12250 12900 12256 12912
rect 12211 12872 12256 12900
rect 12250 12860 12256 12872
rect 12308 12860 12314 12912
rect 13722 12860 13728 12912
rect 13780 12900 13786 12912
rect 20254 12900 20260 12912
rect 13780 12872 18920 12900
rect 13780 12860 13786 12872
rect 11057 12835 11115 12841
rect 10152 12804 10824 12832
rect 9769 12795 9827 12801
rect 9309 12767 9367 12773
rect 9309 12764 9321 12767
rect 9088 12736 9321 12764
rect 9088 12724 9094 12736
rect 9309 12733 9321 12736
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 9398 12724 9404 12776
rect 9456 12764 9462 12776
rect 10042 12764 10048 12776
rect 9456 12736 10048 12764
rect 9456 12724 9462 12736
rect 10042 12724 10048 12736
rect 10100 12764 10106 12776
rect 10796 12773 10824 12804
rect 11057 12801 11069 12835
rect 11103 12832 11115 12835
rect 11974 12832 11980 12844
rect 11103 12804 11980 12832
rect 11103 12801 11115 12804
rect 11057 12795 11115 12801
rect 11974 12792 11980 12804
rect 12032 12792 12038 12844
rect 12526 12832 12532 12844
rect 12487 12804 12532 12832
rect 12526 12792 12532 12804
rect 12584 12792 12590 12844
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 12805 12835 12863 12841
rect 12805 12832 12817 12835
rect 12768 12804 12817 12832
rect 12768 12792 12774 12804
rect 12805 12801 12817 12804
rect 12851 12801 12863 12835
rect 13446 12832 13452 12844
rect 13407 12804 13452 12832
rect 12805 12795 12863 12801
rect 13446 12792 13452 12804
rect 13504 12832 13510 12844
rect 18892 12832 18920 12872
rect 19260 12872 20260 12900
rect 19260 12841 19288 12872
rect 20254 12860 20260 12872
rect 20312 12860 20318 12912
rect 19245 12835 19303 12841
rect 19245 12832 19257 12835
rect 13504 12804 14412 12832
rect 13504 12792 13510 12804
rect 14384 12776 14412 12804
rect 18892 12804 19257 12832
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 10100 12736 10333 12764
rect 10100 12724 10106 12736
rect 10321 12733 10333 12736
rect 10367 12733 10379 12767
rect 10321 12727 10379 12733
rect 10781 12767 10839 12773
rect 10781 12733 10793 12767
rect 10827 12733 10839 12767
rect 14366 12764 14372 12776
rect 14279 12736 14372 12764
rect 10781 12727 10839 12733
rect 14366 12724 14372 12736
rect 14424 12724 14430 12776
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12733 14887 12767
rect 15286 12764 15292 12776
rect 15247 12736 15292 12764
rect 14829 12727 14887 12733
rect 7616 12668 7880 12696
rect 7616 12656 7622 12668
rect 12618 12656 12624 12708
rect 12676 12696 12682 12708
rect 12676 12668 12721 12696
rect 12676 12656 12682 12668
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 4062 12628 4068 12640
rect 4019 12600 4068 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 6178 12628 6184 12640
rect 6139 12600 6184 12628
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 9490 12628 9496 12640
rect 9451 12600 9496 12628
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 10042 12588 10048 12640
rect 10100 12628 10106 12640
rect 10962 12628 10968 12640
rect 10100 12600 10968 12628
rect 10100 12588 10106 12600
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 11333 12631 11391 12637
rect 11333 12628 11345 12631
rect 11296 12600 11345 12628
rect 11296 12588 11302 12600
rect 11333 12597 11345 12600
rect 11379 12597 11391 12631
rect 13814 12628 13820 12640
rect 13775 12600 13820 12628
rect 11333 12591 11391 12597
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 14182 12628 14188 12640
rect 14143 12600 14188 12628
rect 14182 12588 14188 12600
rect 14240 12628 14246 12640
rect 14844 12628 14872 12727
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 15562 12764 15568 12776
rect 15523 12736 15568 12764
rect 15562 12724 15568 12736
rect 15620 12764 15626 12776
rect 16942 12764 16948 12776
rect 15620 12736 16948 12764
rect 15620 12724 15626 12736
rect 16942 12724 16948 12736
rect 17000 12764 17006 12776
rect 18892 12773 18920 12804
rect 19245 12801 19257 12804
rect 19291 12801 19303 12835
rect 19245 12795 19303 12801
rect 19518 12792 19524 12844
rect 19576 12832 19582 12844
rect 19981 12835 20039 12841
rect 19981 12832 19993 12835
rect 19576 12804 19993 12832
rect 19576 12792 19582 12804
rect 19981 12801 19993 12804
rect 20027 12801 20039 12835
rect 20622 12832 20628 12844
rect 20583 12804 20628 12832
rect 19981 12795 20039 12801
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 17037 12767 17095 12773
rect 17037 12764 17049 12767
rect 17000 12736 17049 12764
rect 17000 12724 17006 12736
rect 17037 12733 17049 12736
rect 17083 12733 17095 12767
rect 17037 12727 17095 12733
rect 18852 12767 18920 12773
rect 18852 12733 18864 12767
rect 18898 12736 18920 12767
rect 18898 12733 18910 12736
rect 18852 12727 18910 12733
rect 21358 12724 21364 12776
rect 21416 12764 21422 12776
rect 21488 12767 21546 12773
rect 21488 12764 21500 12767
rect 21416 12736 21500 12764
rect 21416 12724 21422 12736
rect 21488 12733 21500 12736
rect 21534 12764 21546 12767
rect 21913 12767 21971 12773
rect 21913 12764 21925 12767
rect 21534 12736 21925 12764
rect 21534 12733 21546 12736
rect 21488 12727 21546 12733
rect 21913 12733 21925 12736
rect 21959 12733 21971 12767
rect 21913 12727 21971 12733
rect 22462 12724 22468 12776
rect 22520 12773 22526 12776
rect 22520 12767 22558 12773
rect 22546 12764 22558 12767
rect 22925 12767 22983 12773
rect 22925 12764 22937 12767
rect 22546 12736 22937 12764
rect 22546 12733 22558 12736
rect 22520 12727 22558 12733
rect 22925 12733 22937 12736
rect 22971 12733 22983 12767
rect 22925 12727 22983 12733
rect 22520 12724 22526 12727
rect 15838 12696 15844 12708
rect 15799 12668 15844 12696
rect 15838 12656 15844 12668
rect 15896 12656 15902 12708
rect 16850 12696 16856 12708
rect 16316 12668 16856 12696
rect 14240 12600 14872 12628
rect 14240 12588 14246 12600
rect 15562 12588 15568 12640
rect 15620 12628 15626 12640
rect 16316 12637 16344 12668
rect 16850 12656 16856 12668
rect 16908 12656 16914 12708
rect 20073 12699 20131 12705
rect 20073 12665 20085 12699
rect 20119 12696 20131 12699
rect 20990 12696 20996 12708
rect 20119 12668 20996 12696
rect 20119 12665 20131 12668
rect 20073 12659 20131 12665
rect 16301 12631 16359 12637
rect 16301 12628 16313 12631
rect 15620 12600 16313 12628
rect 15620 12588 15626 12600
rect 16301 12597 16313 12600
rect 16347 12597 16359 12631
rect 16666 12628 16672 12640
rect 16627 12600 16672 12628
rect 16301 12591 16359 12597
rect 16666 12588 16672 12600
rect 16724 12588 16730 12640
rect 19797 12631 19855 12637
rect 19797 12597 19809 12631
rect 19843 12628 19855 12631
rect 20088 12628 20116 12659
rect 20990 12656 20996 12668
rect 21048 12656 21054 12708
rect 19843 12600 20116 12628
rect 19843 12597 19855 12600
rect 19797 12591 19855 12597
rect 21174 12588 21180 12640
rect 21232 12628 21238 12640
rect 22646 12637 22652 12640
rect 21591 12631 21649 12637
rect 21591 12628 21603 12631
rect 21232 12600 21603 12628
rect 21232 12588 21238 12600
rect 21591 12597 21603 12600
rect 21637 12597 21649 12631
rect 21591 12591 21649 12597
rect 22603 12631 22652 12637
rect 22603 12597 22615 12631
rect 22649 12597 22652 12631
rect 22603 12591 22652 12597
rect 22646 12588 22652 12591
rect 22704 12588 22710 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 5261 12427 5319 12433
rect 5261 12424 5273 12427
rect 4212 12396 5273 12424
rect 4212 12384 4218 12396
rect 5261 12393 5273 12396
rect 5307 12393 5319 12427
rect 12066 12424 12072 12436
rect 12027 12396 12072 12424
rect 5261 12387 5319 12393
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 15286 12424 15292 12436
rect 13872 12396 15292 12424
rect 13872 12384 13878 12396
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 20898 12384 20904 12436
rect 20956 12424 20962 12436
rect 24762 12424 24768 12436
rect 20956 12396 21128 12424
rect 24723 12396 24768 12424
rect 20956 12384 20962 12396
rect 6178 12356 6184 12368
rect 2424 12328 6184 12356
rect 2424 12297 2452 12328
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12288 2375 12291
rect 2409 12291 2467 12297
rect 2409 12288 2421 12291
rect 2363 12260 2421 12288
rect 2363 12257 2375 12260
rect 2317 12251 2375 12257
rect 2409 12257 2421 12260
rect 2455 12257 2467 12291
rect 2682 12288 2688 12300
rect 2643 12260 2688 12288
rect 2409 12251 2467 12257
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 4614 12248 4620 12300
rect 4672 12288 4678 12300
rect 4816 12297 4844 12328
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 7558 12356 7564 12368
rect 7519 12328 7564 12356
rect 7558 12316 7564 12328
rect 7616 12316 7622 12368
rect 12805 12359 12863 12365
rect 12805 12325 12817 12359
rect 12851 12356 12863 12359
rect 14458 12356 14464 12368
rect 12851 12328 14464 12356
rect 12851 12325 12863 12328
rect 12805 12319 12863 12325
rect 4709 12291 4767 12297
rect 4709 12288 4721 12291
rect 4672 12260 4721 12288
rect 4672 12248 4678 12260
rect 4709 12257 4721 12260
rect 4755 12288 4767 12291
rect 4801 12291 4859 12297
rect 4801 12288 4813 12291
rect 4755 12260 4813 12288
rect 4755 12257 4767 12260
rect 4709 12251 4767 12257
rect 4801 12257 4813 12260
rect 4847 12257 4859 12291
rect 4801 12251 4859 12257
rect 4890 12248 4896 12300
rect 4948 12288 4954 12300
rect 5077 12291 5135 12297
rect 4948 12260 4993 12288
rect 4948 12248 4954 12260
rect 5077 12257 5089 12291
rect 5123 12288 5135 12291
rect 5166 12288 5172 12300
rect 5123 12260 5172 12288
rect 5123 12257 5135 12260
rect 5077 12251 5135 12257
rect 2038 12180 2044 12232
rect 2096 12220 2102 12232
rect 2869 12223 2927 12229
rect 2869 12220 2881 12223
rect 2096 12192 2881 12220
rect 2096 12180 2102 12192
rect 2869 12189 2881 12192
rect 2915 12189 2927 12223
rect 2869 12183 2927 12189
rect 4154 12180 4160 12232
rect 4212 12220 4218 12232
rect 5092 12220 5120 12251
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 6362 12288 6368 12300
rect 5592 12260 6368 12288
rect 5592 12248 5598 12260
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 7190 12288 7196 12300
rect 7151 12260 7196 12288
rect 7190 12248 7196 12260
rect 7248 12248 7254 12300
rect 8205 12291 8263 12297
rect 8205 12257 8217 12291
rect 8251 12288 8263 12291
rect 8294 12288 8300 12300
rect 8251 12260 8300 12288
rect 8251 12257 8263 12260
rect 8205 12251 8263 12257
rect 8294 12248 8300 12260
rect 8352 12288 8358 12300
rect 9030 12288 9036 12300
rect 8352 12260 9036 12288
rect 8352 12248 8358 12260
rect 9030 12248 9036 12260
rect 9088 12248 9094 12300
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 9953 12291 10011 12297
rect 9953 12288 9965 12291
rect 9732 12260 9965 12288
rect 9732 12248 9738 12260
rect 9953 12257 9965 12260
rect 9999 12288 10011 12291
rect 10042 12288 10048 12300
rect 9999 12260 10048 12288
rect 9999 12257 10011 12260
rect 9953 12251 10011 12257
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 10134 12248 10140 12300
rect 10192 12288 10198 12300
rect 10410 12288 10416 12300
rect 10192 12260 10416 12288
rect 10192 12248 10198 12260
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 11514 12248 11520 12300
rect 11572 12297 11578 12300
rect 11572 12291 11610 12297
rect 11598 12257 11610 12291
rect 11572 12251 11610 12257
rect 11572 12248 11578 12251
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 12897 12291 12955 12297
rect 12897 12288 12909 12291
rect 12216 12260 12909 12288
rect 12216 12248 12222 12260
rect 12897 12257 12909 12260
rect 12943 12257 12955 12291
rect 13354 12288 13360 12300
rect 13315 12260 13360 12288
rect 12897 12251 12955 12257
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12288 13783 12291
rect 13998 12288 14004 12300
rect 13771 12260 14004 12288
rect 13771 12257 13783 12260
rect 13725 12251 13783 12257
rect 4212 12192 5120 12220
rect 10689 12223 10747 12229
rect 4212 12180 4218 12192
rect 10689 12189 10701 12223
rect 10735 12220 10747 12223
rect 10778 12220 10784 12232
rect 10735 12192 10784 12220
rect 10735 12189 10747 12192
rect 10689 12183 10747 12189
rect 10778 12180 10784 12192
rect 10836 12220 10842 12232
rect 10965 12223 11023 12229
rect 10965 12220 10977 12223
rect 10836 12192 10977 12220
rect 10836 12180 10842 12192
rect 10965 12189 10977 12192
rect 11011 12189 11023 12223
rect 10965 12183 11023 12189
rect 11425 12223 11483 12229
rect 11425 12189 11437 12223
rect 11471 12220 11483 12223
rect 11698 12220 11704 12232
rect 11471 12192 11704 12220
rect 11471 12189 11483 12192
rect 11425 12183 11483 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 13740 12220 13768 12251
rect 13998 12248 14004 12260
rect 14056 12248 14062 12300
rect 14108 12297 14136 12328
rect 14458 12316 14464 12328
rect 14516 12316 14522 12368
rect 18874 12316 18880 12368
rect 18932 12356 18938 12368
rect 21100 12365 21128 12396
rect 24762 12384 24768 12396
rect 24820 12384 24826 12436
rect 19106 12359 19164 12365
rect 19106 12356 19118 12359
rect 18932 12328 19118 12356
rect 18932 12316 18938 12328
rect 19106 12325 19118 12328
rect 19152 12325 19164 12359
rect 19106 12319 19164 12325
rect 21085 12359 21143 12365
rect 21085 12325 21097 12359
rect 21131 12325 21143 12359
rect 21085 12319 21143 12325
rect 14093 12291 14151 12297
rect 14093 12257 14105 12291
rect 14139 12257 14151 12291
rect 15286 12288 15292 12300
rect 15247 12260 15292 12288
rect 14093 12251 14151 12257
rect 15286 12248 15292 12260
rect 15344 12288 15350 12300
rect 15749 12291 15807 12297
rect 15749 12288 15761 12291
rect 15344 12260 15761 12288
rect 15344 12248 15350 12260
rect 15749 12257 15761 12260
rect 15795 12257 15807 12291
rect 15749 12251 15807 12257
rect 16301 12291 16359 12297
rect 16301 12257 16313 12291
rect 16347 12257 16359 12291
rect 16758 12288 16764 12300
rect 16719 12260 16764 12288
rect 16301 12251 16359 12257
rect 12636 12192 13768 12220
rect 2498 12152 2504 12164
rect 2459 12124 2504 12152
rect 2498 12112 2504 12124
rect 2556 12112 2562 12164
rect 8754 12152 8760 12164
rect 8715 12124 8760 12152
rect 8754 12112 8760 12124
rect 8812 12112 8818 12164
rect 12636 12096 12664 12192
rect 15470 12180 15476 12232
rect 15528 12220 15534 12232
rect 16022 12220 16028 12232
rect 15528 12192 16028 12220
rect 15528 12180 15534 12192
rect 16022 12180 16028 12192
rect 16080 12220 16086 12232
rect 16117 12223 16175 12229
rect 16117 12220 16129 12223
rect 16080 12192 16129 12220
rect 16080 12180 16086 12192
rect 16117 12189 16129 12192
rect 16163 12220 16175 12223
rect 16316 12220 16344 12251
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 17126 12288 17132 12300
rect 17087 12260 17132 12288
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17494 12288 17500 12300
rect 17455 12260 17500 12288
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 18782 12288 18788 12300
rect 18743 12260 18788 12288
rect 18782 12248 18788 12260
rect 18840 12248 18846 12300
rect 22462 12248 22468 12300
rect 22520 12297 22526 12300
rect 22520 12291 22558 12297
rect 22546 12257 22558 12291
rect 22520 12251 22558 12257
rect 22520 12248 22526 12251
rect 20990 12220 20996 12232
rect 16163 12192 16344 12220
rect 20951 12192 20996 12220
rect 16163 12189 16175 12192
rect 16117 12183 16175 12189
rect 20990 12180 20996 12192
rect 21048 12180 21054 12232
rect 21082 12180 21088 12232
rect 21140 12220 21146 12232
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 21140 12192 21281 12220
rect 21140 12180 21146 12192
rect 21269 12189 21281 12192
rect 21315 12220 21327 12223
rect 21913 12223 21971 12229
rect 21913 12220 21925 12223
rect 21315 12192 21925 12220
rect 21315 12189 21327 12192
rect 21269 12183 21327 12189
rect 21913 12189 21925 12192
rect 21959 12189 21971 12223
rect 21913 12183 21971 12189
rect 14274 12152 14280 12164
rect 14235 12124 14280 12152
rect 14274 12112 14280 12124
rect 14332 12112 14338 12164
rect 17678 12152 17684 12164
rect 17639 12124 17684 12152
rect 17678 12112 17684 12124
rect 17736 12112 17742 12164
rect 6546 12084 6552 12096
rect 6507 12056 6552 12084
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 11422 12044 11428 12096
rect 11480 12084 11486 12096
rect 11655 12087 11713 12093
rect 11655 12084 11667 12087
rect 11480 12056 11667 12084
rect 11480 12044 11486 12056
rect 11655 12053 11667 12056
rect 11701 12053 11713 12087
rect 11655 12047 11713 12053
rect 12434 12044 12440 12096
rect 12492 12084 12498 12096
rect 12618 12084 12624 12096
rect 12492 12056 12624 12084
rect 12492 12044 12498 12056
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 14642 12084 14648 12096
rect 14424 12056 14648 12084
rect 14424 12044 14430 12056
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 15473 12087 15531 12093
rect 15473 12053 15485 12087
rect 15519 12084 15531 12087
rect 16390 12084 16396 12096
rect 15519 12056 16396 12084
rect 15519 12053 15531 12056
rect 15473 12047 15531 12053
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 19518 12044 19524 12096
rect 19576 12084 19582 12096
rect 19705 12087 19763 12093
rect 19705 12084 19717 12087
rect 19576 12056 19717 12084
rect 19576 12044 19582 12056
rect 19705 12053 19717 12056
rect 19751 12053 19763 12087
rect 19705 12047 19763 12053
rect 22186 12044 22192 12096
rect 22244 12084 22250 12096
rect 22603 12087 22661 12093
rect 22603 12084 22615 12087
rect 22244 12056 22615 12084
rect 22244 12044 22250 12056
rect 22603 12053 22615 12056
rect 22649 12053 22661 12087
rect 22603 12047 22661 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1949 11883 2007 11889
rect 1949 11849 1961 11883
rect 1995 11880 2007 11883
rect 2498 11880 2504 11892
rect 1995 11852 2504 11880
rect 1995 11849 2007 11852
rect 1949 11843 2007 11849
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 2593 11883 2651 11889
rect 2593 11849 2605 11883
rect 2639 11880 2651 11883
rect 2682 11880 2688 11892
rect 2639 11852 2688 11880
rect 2639 11849 2651 11852
rect 2593 11843 2651 11849
rect 2682 11840 2688 11852
rect 2740 11880 2746 11892
rect 4154 11880 4160 11892
rect 2740 11852 4160 11880
rect 2740 11840 2746 11852
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 4430 11880 4436 11892
rect 4391 11852 4436 11880
rect 4430 11840 4436 11852
rect 4488 11880 4494 11892
rect 6089 11883 6147 11889
rect 4488 11852 4936 11880
rect 4488 11840 4494 11852
rect 4709 11815 4767 11821
rect 4709 11781 4721 11815
rect 4755 11812 4767 11815
rect 4798 11812 4804 11824
rect 4755 11784 4804 11812
rect 4755 11781 4767 11784
rect 4709 11775 4767 11781
rect 4798 11772 4804 11784
rect 4856 11772 4862 11824
rect 2038 11676 2044 11688
rect 1999 11648 2044 11676
rect 2038 11636 2044 11648
rect 2096 11636 2102 11688
rect 3145 11679 3203 11685
rect 3145 11676 3157 11679
rect 2884 11648 3157 11676
rect 2884 11552 2912 11648
rect 3145 11645 3157 11648
rect 3191 11645 3203 11679
rect 3145 11639 3203 11645
rect 3789 11679 3847 11685
rect 3789 11645 3801 11679
rect 3835 11676 3847 11679
rect 4614 11676 4620 11688
rect 3835 11648 4620 11676
rect 3835 11645 3847 11648
rect 3789 11639 3847 11645
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 4908 11685 4936 11852
rect 6089 11849 6101 11883
rect 6135 11880 6147 11883
rect 6178 11880 6184 11892
rect 6135 11852 6184 11880
rect 6135 11849 6147 11852
rect 6089 11843 6147 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 6362 11880 6368 11892
rect 6323 11852 6368 11880
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 8294 11880 8300 11892
rect 8255 11852 8300 11880
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 8570 11880 8576 11892
rect 8531 11852 8576 11880
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 10045 11883 10103 11889
rect 10045 11849 10057 11883
rect 10091 11880 10103 11883
rect 10410 11880 10416 11892
rect 10091 11852 10416 11880
rect 10091 11849 10103 11852
rect 10045 11843 10103 11849
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11572 11852 11805 11880
rect 11572 11840 11578 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 11793 11843 11851 11849
rect 12713 11883 12771 11889
rect 12713 11849 12725 11883
rect 12759 11880 12771 11883
rect 12894 11880 12900 11892
rect 12759 11852 12900 11880
rect 12759 11849 12771 11852
rect 12713 11843 12771 11849
rect 12894 11840 12900 11852
rect 12952 11880 12958 11892
rect 13354 11880 13360 11892
rect 12952 11852 13360 11880
rect 12952 11840 12958 11852
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 14182 11880 14188 11892
rect 14143 11852 14188 11880
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 18417 11883 18475 11889
rect 18417 11849 18429 11883
rect 18463 11880 18475 11883
rect 18693 11883 18751 11889
rect 18693 11880 18705 11883
rect 18463 11852 18705 11880
rect 18463 11849 18475 11852
rect 18417 11843 18475 11849
rect 18693 11849 18705 11852
rect 18739 11880 18751 11883
rect 18874 11880 18880 11892
rect 18739 11852 18880 11880
rect 18739 11849 18751 11852
rect 18693 11843 18751 11849
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 20625 11883 20683 11889
rect 20625 11849 20637 11883
rect 20671 11880 20683 11883
rect 20990 11880 20996 11892
rect 20671 11852 20996 11880
rect 20671 11849 20683 11852
rect 20625 11843 20683 11849
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 7101 11815 7159 11821
rect 7101 11781 7113 11815
rect 7147 11812 7159 11815
rect 7285 11815 7343 11821
rect 7285 11812 7297 11815
rect 7147 11784 7297 11812
rect 7147 11781 7159 11784
rect 7101 11775 7159 11781
rect 7285 11781 7297 11784
rect 7331 11812 7343 11815
rect 7834 11812 7840 11824
rect 7331 11784 7840 11812
rect 7331 11781 7343 11784
rect 7285 11775 7343 11781
rect 7834 11772 7840 11784
rect 7892 11772 7898 11824
rect 8754 11772 8760 11824
rect 8812 11812 8818 11824
rect 8849 11815 8907 11821
rect 8849 11812 8861 11815
rect 8812 11784 8861 11812
rect 8812 11772 8818 11784
rect 8849 11781 8861 11784
rect 8895 11781 8907 11815
rect 8849 11775 8907 11781
rect 5350 11744 5356 11756
rect 5311 11716 5356 11744
rect 5350 11704 5356 11716
rect 5408 11704 5414 11756
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11744 7987 11747
rect 8202 11744 8208 11756
rect 7975 11716 8208 11744
rect 7975 11713 7987 11716
rect 7929 11707 7987 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 14200 11744 14228 11840
rect 17494 11812 17500 11824
rect 15764 11784 17500 11812
rect 14200 11716 14872 11744
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11645 4951 11679
rect 7190 11676 7196 11688
rect 7151 11648 7196 11676
rect 4893 11639 4951 11645
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 7374 11636 7380 11688
rect 7432 11676 7438 11688
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 7432 11648 7481 11676
rect 7432 11636 7438 11648
rect 7469 11645 7481 11648
rect 7515 11645 7527 11679
rect 7469 11639 7527 11645
rect 8570 11636 8576 11688
rect 8628 11676 8634 11688
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 8628 11648 8769 11676
rect 8628 11636 8634 11648
rect 8757 11645 8769 11648
rect 8803 11645 8815 11679
rect 9030 11676 9036 11688
rect 8991 11648 9036 11676
rect 8757 11639 8815 11645
rect 9030 11636 9036 11648
rect 9088 11636 9094 11688
rect 11425 11679 11483 11685
rect 11425 11645 11437 11679
rect 11471 11676 11483 11679
rect 11698 11676 11704 11688
rect 11471 11648 11704 11676
rect 11471 11645 11483 11648
rect 11425 11639 11483 11645
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 12066 11636 12072 11688
rect 12124 11676 12130 11688
rect 13449 11679 13507 11685
rect 13449 11676 13461 11679
rect 12124 11648 13461 11676
rect 12124 11636 12130 11648
rect 13449 11645 13461 11648
rect 13495 11676 13507 11679
rect 13630 11676 13636 11688
rect 13495 11648 13636 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 14642 11676 14648 11688
rect 13955 11648 14648 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 14844 11685 14872 11716
rect 15764 11688 15792 11784
rect 17494 11772 17500 11784
rect 17552 11772 17558 11824
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 18877 11747 18935 11753
rect 18877 11744 18889 11747
rect 15887 11716 18889 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 18877 11713 18889 11716
rect 18923 11744 18935 11747
rect 20073 11747 20131 11753
rect 20073 11744 20085 11747
rect 18923 11716 20085 11744
rect 18923 11713 18935 11716
rect 18877 11707 18935 11713
rect 20073 11713 20085 11716
rect 20119 11713 20131 11747
rect 20073 11707 20131 11713
rect 14829 11679 14887 11685
rect 14829 11645 14841 11679
rect 14875 11645 14887 11679
rect 15378 11676 15384 11688
rect 15339 11648 15384 11676
rect 14829 11639 14887 11645
rect 4798 11568 4804 11620
rect 4856 11608 4862 11620
rect 5629 11611 5687 11617
rect 5629 11608 5641 11611
rect 4856 11580 5641 11608
rect 4856 11568 4862 11580
rect 5629 11577 5641 11580
rect 5675 11577 5687 11611
rect 5629 11571 5687 11577
rect 2222 11540 2228 11552
rect 2183 11512 2228 11540
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 2866 11540 2872 11552
rect 2827 11512 2872 11540
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 7208 11540 7236 11636
rect 9490 11608 9496 11620
rect 9451 11580 9496 11608
rect 9490 11568 9496 11580
rect 9548 11568 9554 11620
rect 13541 11611 13599 11617
rect 13541 11577 13553 11611
rect 13587 11608 13599 11611
rect 13722 11608 13728 11620
rect 13587 11580 13728 11608
rect 13587 11577 13599 11580
rect 13541 11571 13599 11577
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 14844 11608 14872 11639
rect 15378 11636 15384 11648
rect 15436 11636 15442 11688
rect 15746 11676 15752 11688
rect 15707 11648 15752 11676
rect 15746 11636 15752 11648
rect 15804 11636 15810 11688
rect 16669 11679 16727 11685
rect 16669 11676 16681 11679
rect 16316 11648 16681 11676
rect 16114 11608 16120 11620
rect 14844 11580 16120 11608
rect 16114 11568 16120 11580
rect 16172 11608 16178 11620
rect 16316 11617 16344 11648
rect 16669 11645 16681 11648
rect 16715 11676 16727 11679
rect 16758 11676 16764 11688
rect 16715 11648 16764 11676
rect 16715 11645 16727 11648
rect 16669 11639 16727 11645
rect 16758 11636 16764 11648
rect 16816 11676 16822 11688
rect 17129 11679 17187 11685
rect 17129 11676 17141 11679
rect 16816 11648 17141 11676
rect 16816 11636 16822 11648
rect 17129 11645 17141 11648
rect 17175 11645 17187 11679
rect 17129 11639 17187 11645
rect 19797 11679 19855 11685
rect 19797 11645 19809 11679
rect 19843 11676 19855 11679
rect 19843 11648 21036 11676
rect 19843 11645 19855 11648
rect 19797 11639 19855 11645
rect 16301 11611 16359 11617
rect 16301 11608 16313 11611
rect 16172 11580 16313 11608
rect 16172 11568 16178 11580
rect 16301 11577 16313 11580
rect 16347 11577 16359 11611
rect 16301 11571 16359 11577
rect 18874 11568 18880 11620
rect 18932 11608 18938 11620
rect 19198 11611 19256 11617
rect 19198 11608 19210 11611
rect 18932 11580 19210 11608
rect 18932 11568 18938 11580
rect 19198 11577 19210 11580
rect 19244 11577 19256 11611
rect 19198 11571 19256 11577
rect 8386 11540 8392 11552
rect 7208 11512 8392 11540
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 10321 11543 10379 11549
rect 10321 11540 10333 11543
rect 9732 11512 10333 11540
rect 9732 11500 9738 11512
rect 10321 11509 10333 11512
rect 10367 11509 10379 11543
rect 10321 11503 10379 11509
rect 10962 11500 10968 11552
rect 11020 11540 11026 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 11020 11512 11069 11540
rect 11020 11500 11026 11512
rect 11057 11509 11069 11512
rect 11103 11509 11115 11543
rect 12158 11540 12164 11552
rect 12119 11512 12164 11540
rect 11057 11503 11115 11509
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 16853 11543 16911 11549
rect 16853 11540 16865 11543
rect 16632 11512 16865 11540
rect 16632 11500 16638 11512
rect 16853 11509 16865 11512
rect 16899 11509 16911 11543
rect 20898 11540 20904 11552
rect 20859 11512 20904 11540
rect 16853 11503 16911 11509
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 21008 11540 21036 11648
rect 21082 11568 21088 11620
rect 21140 11608 21146 11620
rect 21453 11611 21511 11617
rect 21453 11608 21465 11611
rect 21140 11580 21465 11608
rect 21140 11568 21146 11580
rect 21453 11577 21465 11580
rect 21499 11577 21511 11611
rect 21453 11571 21511 11577
rect 21545 11611 21603 11617
rect 21545 11577 21557 11611
rect 21591 11577 21603 11611
rect 22094 11608 22100 11620
rect 22055 11580 22100 11608
rect 21545 11571 21603 11577
rect 21358 11540 21364 11552
rect 21008 11512 21364 11540
rect 21358 11500 21364 11512
rect 21416 11540 21422 11552
rect 21560 11540 21588 11571
rect 22094 11568 22100 11580
rect 22152 11568 22158 11620
rect 22462 11540 22468 11552
rect 21416 11512 21588 11540
rect 22423 11512 22468 11540
rect 21416 11500 21422 11512
rect 22462 11500 22468 11512
rect 22520 11500 22526 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 4709 11339 4767 11345
rect 4709 11305 4721 11339
rect 4755 11336 4767 11339
rect 4798 11336 4804 11348
rect 4755 11308 4804 11336
rect 4755 11305 4767 11308
rect 4709 11299 4767 11305
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 6512 11308 6745 11336
rect 6512 11296 6518 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 7926 11336 7932 11348
rect 7887 11308 7932 11336
rect 6733 11299 6791 11305
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 9030 11336 9036 11348
rect 8680 11308 9036 11336
rect 5442 11268 5448 11280
rect 2700 11240 5448 11268
rect 2222 11160 2228 11212
rect 2280 11200 2286 11212
rect 2409 11203 2467 11209
rect 2409 11200 2421 11203
rect 2280 11172 2421 11200
rect 2280 11160 2286 11172
rect 2409 11169 2421 11172
rect 2455 11169 2467 11203
rect 2409 11163 2467 11169
rect 2501 11203 2559 11209
rect 2501 11169 2513 11203
rect 2547 11200 2559 11203
rect 2590 11200 2596 11212
rect 2547 11172 2596 11200
rect 2547 11169 2559 11172
rect 2501 11163 2559 11169
rect 2590 11160 2596 11172
rect 2648 11160 2654 11212
rect 2700 11209 2728 11240
rect 5442 11228 5448 11240
rect 5500 11268 5506 11280
rect 7374 11268 7380 11280
rect 5500 11240 7380 11268
rect 5500 11228 5506 11240
rect 7374 11228 7380 11240
rect 7432 11268 7438 11280
rect 8680 11268 8708 11308
rect 9030 11296 9036 11308
rect 9088 11296 9094 11348
rect 10134 11336 10140 11348
rect 10095 11308 10140 11336
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 12066 11336 12072 11348
rect 12027 11308 12072 11336
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 14461 11339 14519 11345
rect 12492 11308 12537 11336
rect 12492 11296 12498 11308
rect 14461 11305 14473 11339
rect 14507 11336 14519 11339
rect 15378 11336 15384 11348
rect 14507 11308 15384 11336
rect 14507 11305 14519 11308
rect 14461 11299 14519 11305
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 15654 11296 15660 11348
rect 15712 11336 15718 11348
rect 15749 11339 15807 11345
rect 15749 11336 15761 11339
rect 15712 11308 15761 11336
rect 15712 11296 15718 11308
rect 15749 11305 15761 11308
rect 15795 11336 15807 11339
rect 16301 11339 16359 11345
rect 16301 11336 16313 11339
rect 15795 11308 16313 11336
rect 15795 11305 15807 11308
rect 15749 11299 15807 11305
rect 16301 11305 16313 11308
rect 16347 11336 16359 11339
rect 16666 11336 16672 11348
rect 16347 11308 16672 11336
rect 16347 11305 16359 11308
rect 16301 11299 16359 11305
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 18782 11336 18788 11348
rect 18743 11308 18788 11336
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 21358 11336 21364 11348
rect 21319 11308 21364 11336
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 7432 11240 8708 11268
rect 7432 11228 7438 11240
rect 8754 11228 8760 11280
rect 8812 11268 8818 11280
rect 9858 11268 9864 11280
rect 8812 11240 9864 11268
rect 8812 11228 8818 11240
rect 9858 11228 9864 11240
rect 9916 11268 9922 11280
rect 9916 11240 10364 11268
rect 9916 11228 9922 11240
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11169 2743 11203
rect 2685 11163 2743 11169
rect 2038 11092 2044 11144
rect 2096 11132 2102 11144
rect 2700 11132 2728 11163
rect 4890 11160 4896 11212
rect 4948 11200 4954 11212
rect 4985 11203 5043 11209
rect 4985 11200 4997 11203
rect 4948 11172 4997 11200
rect 4948 11160 4954 11172
rect 4985 11169 4997 11172
rect 5031 11169 5043 11203
rect 5258 11200 5264 11212
rect 5219 11172 5264 11200
rect 4985 11163 5043 11169
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 6454 11160 6460 11212
rect 6512 11200 6518 11212
rect 6549 11203 6607 11209
rect 6549 11200 6561 11203
rect 6512 11172 6561 11200
rect 6512 11160 6518 11172
rect 6549 11169 6561 11172
rect 6595 11200 6607 11203
rect 7009 11203 7067 11209
rect 7009 11200 7021 11203
rect 6595 11172 7021 11200
rect 6595 11169 6607 11172
rect 6549 11163 6607 11169
rect 7009 11169 7021 11172
rect 7055 11169 7067 11203
rect 7009 11163 7067 11169
rect 7834 11160 7840 11212
rect 7892 11200 7898 11212
rect 8021 11203 8079 11209
rect 8021 11200 8033 11203
rect 7892 11172 8033 11200
rect 7892 11160 7898 11172
rect 8021 11169 8033 11172
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11169 8539 11203
rect 10042 11200 10048 11212
rect 10003 11172 10048 11200
rect 8481 11163 8539 11169
rect 3142 11132 3148 11144
rect 2096 11104 2728 11132
rect 3103 11104 3148 11132
rect 2096 11092 2102 11104
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11132 5779 11135
rect 6822 11132 6828 11144
rect 5767 11104 6828 11132
rect 5767 11101 5779 11104
rect 5721 11095 5779 11101
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 5074 11064 5080 11076
rect 5035 11036 5080 11064
rect 5074 11024 5080 11036
rect 5132 11024 5138 11076
rect 8496 11064 8524 11163
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10336 11209 10364 11240
rect 12250 11228 12256 11280
rect 12308 11268 12314 11280
rect 15562 11268 15568 11280
rect 12308 11240 15568 11268
rect 12308 11228 12314 11240
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11169 10379 11203
rect 10689 11203 10747 11209
rect 10689 11200 10701 11203
rect 10321 11163 10379 11169
rect 10612 11172 10701 11200
rect 8757 11135 8815 11141
rect 8757 11101 8769 11135
rect 8803 11132 8815 11135
rect 9582 11132 9588 11144
rect 8803 11104 9588 11132
rect 8803 11101 8815 11104
rect 8757 11095 8815 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 10612 11064 10640 11172
rect 10689 11169 10701 11172
rect 10735 11169 10747 11203
rect 11054 11200 11060 11212
rect 11015 11172 11060 11200
rect 10689 11163 10747 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 12158 11200 12164 11212
rect 12119 11172 12164 11200
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 12894 11200 12900 11212
rect 12855 11172 12900 11200
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 13004 11209 13032 11240
rect 15562 11228 15568 11240
rect 15620 11228 15626 11280
rect 16684 11268 16712 11296
rect 17126 11268 17132 11280
rect 16684 11240 17132 11268
rect 17126 11228 17132 11240
rect 17184 11268 17190 11280
rect 19981 11271 20039 11277
rect 17184 11240 17356 11268
rect 17184 11228 17190 11240
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11169 13047 11203
rect 13538 11200 13544 11212
rect 13499 11172 13544 11200
rect 12989 11163 13047 11169
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 15286 11200 15292 11212
rect 15247 11172 15292 11200
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 16390 11160 16396 11212
rect 16448 11200 16454 11212
rect 16485 11203 16543 11209
rect 16485 11200 16497 11203
rect 16448 11172 16497 11200
rect 16448 11160 16454 11172
rect 16485 11169 16497 11172
rect 16531 11169 16543 11203
rect 16485 11163 16543 11169
rect 16574 11160 16580 11212
rect 16632 11200 16638 11212
rect 17328 11209 17356 11240
rect 19981 11237 19993 11271
rect 20027 11268 20039 11271
rect 20898 11268 20904 11280
rect 20027 11240 20904 11268
rect 20027 11237 20039 11240
rect 19981 11231 20039 11237
rect 20898 11228 20904 11240
rect 20956 11228 20962 11280
rect 21910 11268 21916 11280
rect 21871 11240 21916 11268
rect 21910 11228 21916 11240
rect 21968 11228 21974 11280
rect 22094 11228 22100 11280
rect 22152 11268 22158 11280
rect 22465 11271 22523 11277
rect 22465 11268 22477 11271
rect 22152 11240 22477 11268
rect 22152 11228 22158 11240
rect 22465 11237 22477 11240
rect 22511 11237 22523 11271
rect 22465 11231 22523 11237
rect 16945 11203 17003 11209
rect 16945 11200 16957 11203
rect 16632 11172 16957 11200
rect 16632 11160 16638 11172
rect 16945 11169 16957 11172
rect 16991 11169 17003 11203
rect 16945 11163 17003 11169
rect 17313 11203 17371 11209
rect 17313 11169 17325 11203
rect 17359 11169 17371 11203
rect 17313 11163 17371 11169
rect 17494 11160 17500 11212
rect 17552 11200 17558 11212
rect 17681 11203 17739 11209
rect 17681 11200 17693 11203
rect 17552 11172 17693 11200
rect 17552 11160 17558 11172
rect 17681 11169 17693 11172
rect 17727 11169 17739 11203
rect 19518 11200 19524 11212
rect 19479 11172 19524 11200
rect 17681 11163 17739 11169
rect 19518 11160 19524 11172
rect 19576 11160 19582 11212
rect 24118 11160 24124 11212
rect 24176 11200 24182 11212
rect 24340 11203 24398 11209
rect 24340 11200 24352 11203
rect 24176 11172 24352 11200
rect 24176 11160 24182 11172
rect 24340 11169 24352 11172
rect 24386 11169 24398 11203
rect 24340 11163 24398 11169
rect 21450 11092 21456 11144
rect 21508 11132 21514 11144
rect 21821 11135 21879 11141
rect 21821 11132 21833 11135
rect 21508 11104 21833 11132
rect 21508 11092 21514 11104
rect 21821 11101 21833 11104
rect 21867 11132 21879 11135
rect 23293 11135 23351 11141
rect 23293 11132 23305 11135
rect 21867 11104 23305 11132
rect 21867 11101 21879 11104
rect 21821 11095 21879 11101
rect 23293 11101 23305 11104
rect 23339 11101 23351 11135
rect 23293 11095 23351 11101
rect 12250 11064 12256 11076
rect 8312 11036 8524 11064
rect 9600 11036 12256 11064
rect 7926 10956 7932 11008
rect 7984 10996 7990 11008
rect 8312 10996 8340 11036
rect 7984 10968 8340 10996
rect 7984 10956 7990 10968
rect 9398 10956 9404 11008
rect 9456 10996 9462 11008
rect 9600 10996 9628 11036
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 15473 11067 15531 11073
rect 15473 11064 15485 11067
rect 14884 11036 15485 11064
rect 14884 11024 14890 11036
rect 15473 11033 15485 11036
rect 15519 11064 15531 11067
rect 17865 11067 17923 11073
rect 15519 11036 16620 11064
rect 15519 11033 15531 11036
rect 15473 11027 15531 11033
rect 13998 10996 14004 11008
rect 9456 10968 9628 10996
rect 13959 10968 14004 10996
rect 9456 10956 9462 10968
rect 13998 10956 14004 10968
rect 14056 10996 14062 11008
rect 14737 10999 14795 11005
rect 14737 10996 14749 10999
rect 14056 10968 14749 10996
rect 14056 10956 14062 10968
rect 14737 10965 14749 10968
rect 14783 10965 14795 10999
rect 16592 10996 16620 11036
rect 17865 11033 17877 11067
rect 17911 11064 17923 11067
rect 18046 11064 18052 11076
rect 17911 11036 18052 11064
rect 17911 11033 17923 11036
rect 17865 11027 17923 11033
rect 18046 11024 18052 11036
rect 18104 11024 18110 11076
rect 16942 10996 16948 11008
rect 16592 10968 16948 10996
rect 14737 10959 14795 10965
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 24443 10999 24501 11005
rect 24443 10965 24455 10999
rect 24489 10996 24501 10999
rect 24670 10996 24676 11008
rect 24489 10968 24676 10996
rect 24489 10965 24501 10968
rect 24443 10959 24501 10965
rect 24670 10956 24676 10968
rect 24728 10956 24734 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2038 10792 2044 10804
rect 1999 10764 2044 10792
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 2317 10795 2375 10801
rect 2317 10792 2329 10795
rect 2280 10764 2329 10792
rect 2280 10752 2286 10764
rect 2317 10761 2329 10764
rect 2363 10761 2375 10795
rect 2317 10755 2375 10761
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 2961 10795 3019 10801
rect 2961 10792 2973 10795
rect 2832 10764 2973 10792
rect 2832 10752 2838 10764
rect 2961 10761 2973 10764
rect 3007 10761 3019 10795
rect 2961 10755 3019 10761
rect 3142 10752 3148 10804
rect 3200 10792 3206 10804
rect 3329 10795 3387 10801
rect 3329 10792 3341 10795
rect 3200 10764 3341 10792
rect 3200 10752 3206 10764
rect 3329 10761 3341 10764
rect 3375 10761 3387 10795
rect 3329 10755 3387 10761
rect 7834 10752 7840 10804
rect 7892 10792 7898 10804
rect 8021 10795 8079 10801
rect 8021 10792 8033 10795
rect 7892 10764 8033 10792
rect 7892 10752 7898 10764
rect 8021 10761 8033 10764
rect 8067 10761 8079 10795
rect 8021 10755 8079 10761
rect 8386 10752 8392 10804
rect 8444 10792 8450 10804
rect 9398 10792 9404 10804
rect 8444 10764 9404 10792
rect 8444 10752 8450 10764
rect 9398 10752 9404 10764
rect 9456 10792 9462 10804
rect 9493 10795 9551 10801
rect 9493 10792 9505 10795
rect 9456 10764 9505 10792
rect 9456 10752 9462 10764
rect 9493 10761 9505 10764
rect 9539 10761 9551 10795
rect 9493 10755 9551 10761
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 10100 10764 11805 10792
rect 10100 10752 10106 10764
rect 11793 10761 11805 10764
rect 11839 10792 11851 10795
rect 12158 10792 12164 10804
rect 11839 10764 12164 10792
rect 11839 10761 11851 10764
rect 11793 10755 11851 10761
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12250 10752 12256 10804
rect 12308 10792 12314 10804
rect 12713 10795 12771 10801
rect 12308 10764 12353 10792
rect 12308 10752 12314 10764
rect 12713 10761 12725 10795
rect 12759 10792 12771 10795
rect 12894 10792 12900 10804
rect 12759 10764 12900 10792
rect 12759 10761 12771 10764
rect 12713 10755 12771 10761
rect 12894 10752 12900 10764
rect 12952 10792 12958 10804
rect 13173 10795 13231 10801
rect 13173 10792 13185 10795
rect 12952 10764 13185 10792
rect 12952 10752 12958 10764
rect 13173 10761 13185 10764
rect 13219 10761 13231 10795
rect 13173 10755 13231 10761
rect 3694 10724 3700 10736
rect 3655 10696 3700 10724
rect 3694 10684 3700 10696
rect 3752 10684 3758 10736
rect 8294 10684 8300 10736
rect 8352 10724 8358 10736
rect 8352 10696 8800 10724
rect 8352 10684 8358 10696
rect 8478 10656 8484 10668
rect 6564 10628 7144 10656
rect 8439 10628 8484 10656
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 3142 10588 3148 10600
rect 2547 10560 3148 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 3142 10548 3148 10560
rect 3200 10548 3206 10600
rect 3513 10591 3571 10597
rect 3513 10557 3525 10591
rect 3559 10588 3571 10591
rect 4893 10591 4951 10597
rect 3559 10560 4108 10588
rect 3559 10557 3571 10560
rect 3513 10551 3571 10557
rect 4080 10464 4108 10560
rect 4893 10557 4905 10591
rect 4939 10557 4951 10591
rect 4893 10551 4951 10557
rect 4908 10464 4936 10551
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 6564 10597 6592 10628
rect 5905 10591 5963 10597
rect 5905 10588 5917 10591
rect 5592 10560 5917 10588
rect 5592 10548 5598 10560
rect 5905 10557 5917 10560
rect 5951 10588 5963 10591
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 5951 10560 6561 10588
rect 5951 10557 5963 10560
rect 5905 10551 5963 10557
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 5166 10480 5172 10532
rect 5224 10520 5230 10532
rect 5261 10523 5319 10529
rect 5261 10520 5273 10523
rect 5224 10492 5273 10520
rect 5224 10480 5230 10492
rect 5261 10489 5273 10492
rect 5307 10520 5319 10523
rect 6840 10520 6868 10551
rect 6914 10548 6920 10600
rect 6972 10588 6978 10600
rect 7116 10597 7144 10628
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 8772 10665 8800 10696
rect 8757 10659 8815 10665
rect 8757 10625 8769 10659
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10413 10659 10471 10665
rect 10413 10656 10425 10659
rect 10192 10628 10425 10656
rect 10192 10616 10198 10628
rect 10413 10625 10425 10628
rect 10459 10625 10471 10659
rect 13188 10656 13216 10755
rect 16574 10752 16580 10804
rect 16632 10792 16638 10804
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 16632 10764 18245 10792
rect 16632 10752 16638 10764
rect 18233 10761 18245 10764
rect 18279 10761 18291 10795
rect 18233 10755 18291 10761
rect 19518 10752 19524 10804
rect 19576 10792 19582 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 19576 10764 19809 10792
rect 19576 10752 19582 10764
rect 19797 10761 19809 10764
rect 19843 10792 19855 10795
rect 20165 10795 20223 10801
rect 20165 10792 20177 10795
rect 19843 10764 20177 10792
rect 19843 10761 19855 10764
rect 19797 10755 19855 10761
rect 20165 10761 20177 10764
rect 20211 10792 20223 10795
rect 20530 10792 20536 10804
rect 20211 10764 20536 10792
rect 20211 10761 20223 10764
rect 20165 10755 20223 10761
rect 20530 10752 20536 10764
rect 20588 10752 20594 10804
rect 21450 10792 21456 10804
rect 21411 10764 21456 10792
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 21821 10795 21879 10801
rect 21821 10761 21833 10795
rect 21867 10792 21879 10795
rect 21910 10792 21916 10804
rect 21867 10764 21916 10792
rect 21867 10761 21879 10764
rect 21821 10755 21879 10761
rect 21910 10752 21916 10764
rect 21968 10752 21974 10804
rect 24762 10792 24768 10804
rect 24723 10764 24768 10792
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 15286 10724 15292 10736
rect 15247 10696 15292 10724
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 13188 10628 13860 10656
rect 10413 10619 10471 10625
rect 7101 10591 7159 10597
rect 6972 10560 7017 10588
rect 6972 10548 6978 10560
rect 7101 10557 7113 10591
rect 7147 10557 7159 10591
rect 7101 10551 7159 10557
rect 12158 10548 12164 10600
rect 12216 10588 12222 10600
rect 13354 10588 13360 10600
rect 12216 10560 13360 10588
rect 12216 10548 12222 10560
rect 13354 10548 13360 10560
rect 13412 10548 13418 10600
rect 13832 10597 13860 10628
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 17218 10656 17224 10668
rect 14056 10628 14596 10656
rect 14056 10616 14062 10628
rect 14568 10597 14596 10628
rect 16684 10628 17224 10656
rect 16684 10600 16712 10628
rect 17218 10616 17224 10628
rect 17276 10656 17282 10668
rect 17405 10659 17463 10665
rect 17405 10656 17417 10659
rect 17276 10628 17417 10656
rect 17276 10616 17282 10628
rect 17405 10625 17417 10628
rect 17451 10625 17463 10659
rect 20438 10656 20444 10668
rect 20399 10628 20444 10656
rect 17405 10619 17463 10625
rect 20438 10616 20444 10628
rect 20496 10616 20502 10668
rect 21082 10656 21088 10668
rect 21043 10628 21088 10656
rect 21082 10616 21088 10628
rect 21140 10616 21146 10668
rect 21928 10665 21956 10752
rect 21913 10659 21971 10665
rect 21913 10625 21925 10659
rect 21959 10625 21971 10659
rect 21913 10619 21971 10625
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 7558 10520 7564 10532
rect 5307 10492 7564 10520
rect 5307 10489 5319 10492
rect 5261 10483 5319 10489
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 8478 10480 8484 10532
rect 8536 10520 8542 10532
rect 8573 10523 8631 10529
rect 8573 10520 8585 10523
rect 8536 10492 8585 10520
rect 8536 10480 8542 10492
rect 8573 10489 8585 10492
rect 8619 10489 8631 10523
rect 8573 10483 8631 10489
rect 10321 10523 10379 10529
rect 10321 10489 10333 10523
rect 10367 10520 10379 10523
rect 10775 10523 10833 10529
rect 10775 10520 10787 10523
rect 10367 10492 10787 10520
rect 10367 10489 10379 10492
rect 10321 10483 10379 10489
rect 10775 10489 10787 10492
rect 10821 10520 10833 10523
rect 11238 10520 11244 10532
rect 10821 10492 11244 10520
rect 10821 10489 10833 10492
rect 10775 10483 10833 10489
rect 11238 10480 11244 10492
rect 11296 10520 11302 10532
rect 11296 10492 11836 10520
rect 11296 10480 11302 10492
rect 2682 10452 2688 10464
rect 2643 10424 2688 10452
rect 2682 10412 2688 10424
rect 2740 10412 2746 10464
rect 4062 10452 4068 10464
rect 4023 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 4890 10452 4896 10464
rect 4479 10424 4896 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 4890 10412 4896 10424
rect 4948 10452 4954 10464
rect 5537 10455 5595 10461
rect 5537 10452 5549 10455
rect 4948 10424 5549 10452
rect 4948 10412 4954 10424
rect 5537 10421 5549 10424
rect 5583 10452 5595 10455
rect 6638 10452 6644 10464
rect 5583 10424 6644 10452
rect 5583 10421 5595 10424
rect 5537 10415 5595 10421
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 7282 10452 7288 10464
rect 7243 10424 7288 10452
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 9861 10455 9919 10461
rect 9861 10452 9873 10455
rect 9732 10424 9873 10452
rect 9732 10412 9738 10424
rect 9861 10421 9873 10424
rect 9907 10452 9919 10455
rect 11054 10452 11060 10464
rect 9907 10424 11060 10452
rect 9907 10421 9919 10424
rect 9861 10415 9919 10421
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 11333 10455 11391 10461
rect 11333 10421 11345 10455
rect 11379 10452 11391 10455
rect 11698 10452 11704 10464
rect 11379 10424 11704 10452
rect 11379 10421 11391 10424
rect 11333 10415 11391 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 11808 10452 11836 10492
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 14200 10520 14228 10551
rect 15470 10548 15476 10600
rect 15528 10588 15534 10600
rect 15657 10591 15715 10597
rect 15657 10588 15669 10591
rect 15528 10560 15669 10588
rect 15528 10548 15534 10560
rect 15657 10557 15669 10560
rect 15703 10557 15715 10591
rect 16114 10588 16120 10600
rect 16075 10560 16120 10588
rect 15657 10551 15715 10557
rect 16114 10548 16120 10560
rect 16172 10548 16178 10600
rect 16666 10588 16672 10600
rect 16627 10560 16672 10588
rect 16666 10548 16672 10560
rect 16724 10548 16730 10600
rect 16942 10588 16948 10600
rect 16903 10560 16948 10588
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 18693 10591 18751 10597
rect 18693 10557 18705 10591
rect 18739 10588 18751 10591
rect 18877 10591 18935 10597
rect 18877 10588 18889 10591
rect 18739 10560 18889 10588
rect 18739 10557 18751 10560
rect 18693 10551 18751 10557
rect 18877 10557 18889 10560
rect 18923 10588 18935 10591
rect 18966 10588 18972 10600
rect 18923 10560 18972 10588
rect 18923 10557 18935 10560
rect 18877 10551 18935 10557
rect 18966 10548 18972 10560
rect 19024 10548 19030 10600
rect 21358 10548 21364 10600
rect 21416 10588 21422 10600
rect 22002 10588 22008 10600
rect 21416 10560 22008 10588
rect 21416 10548 21422 10560
rect 22002 10548 22008 10560
rect 22060 10548 22066 10600
rect 24118 10548 24124 10600
rect 24176 10588 24182 10600
rect 24302 10588 24308 10600
rect 24176 10560 24308 10588
rect 24176 10548 24182 10560
rect 24302 10548 24308 10560
rect 24360 10548 24366 10600
rect 24581 10591 24639 10597
rect 24581 10557 24593 10591
rect 24627 10588 24639 10591
rect 24670 10588 24676 10600
rect 24627 10560 24676 10588
rect 24627 10557 24639 10560
rect 24581 10551 24639 10557
rect 24670 10548 24676 10560
rect 24728 10588 24734 10600
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24728 10560 25145 10588
rect 24728 10548 24734 10560
rect 25133 10557 25145 10560
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 14826 10520 14832 10532
rect 12676 10492 14228 10520
rect 14787 10492 14832 10520
rect 12676 10480 12682 10492
rect 14826 10480 14832 10492
rect 14884 10480 14890 10532
rect 16390 10480 16396 10532
rect 16448 10520 16454 10532
rect 17773 10523 17831 10529
rect 17773 10520 17785 10523
rect 16448 10492 17785 10520
rect 16448 10480 16454 10492
rect 17773 10489 17785 10492
rect 17819 10489 17831 10523
rect 17773 10483 17831 10489
rect 20530 10480 20536 10532
rect 20588 10520 20594 10532
rect 20588 10492 20633 10520
rect 20588 10480 20594 10492
rect 13078 10452 13084 10464
rect 11808 10424 13084 10452
rect 13078 10412 13084 10424
rect 13136 10412 13142 10464
rect 16850 10452 16856 10464
rect 16811 10424 16856 10452
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 19058 10452 19064 10464
rect 19019 10424 19064 10452
rect 19058 10412 19064 10424
rect 19116 10412 19122 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 4893 10251 4951 10257
rect 4893 10217 4905 10251
rect 4939 10248 4951 10251
rect 5074 10248 5080 10260
rect 4939 10220 5080 10248
rect 4939 10217 4951 10220
rect 4893 10211 4951 10217
rect 5074 10208 5080 10220
rect 5132 10208 5138 10260
rect 7926 10248 7932 10260
rect 7887 10220 7932 10248
rect 7926 10208 7932 10220
rect 7984 10248 7990 10260
rect 8386 10248 8392 10260
rect 7984 10220 8392 10248
rect 7984 10208 7990 10220
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 10192 10220 10885 10248
rect 10192 10208 10198 10220
rect 10873 10217 10885 10220
rect 10919 10217 10931 10251
rect 12066 10248 12072 10260
rect 10873 10211 10931 10217
rect 11348 10220 12072 10248
rect 5721 10183 5779 10189
rect 5721 10149 5733 10183
rect 5767 10180 5779 10183
rect 6454 10180 6460 10192
rect 5767 10152 6460 10180
rect 5767 10149 5779 10152
rect 5721 10143 5779 10149
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 6730 10140 6736 10192
rect 6788 10180 6794 10192
rect 8110 10180 8116 10192
rect 6788 10152 8116 10180
rect 6788 10140 6794 10152
rect 8110 10140 8116 10152
rect 8168 10140 8174 10192
rect 8202 10140 8208 10192
rect 8260 10180 8266 10192
rect 8260 10152 8305 10180
rect 8260 10140 8266 10152
rect 10042 10140 10048 10192
rect 10100 10180 10106 10192
rect 11348 10189 11376 10220
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 12618 10248 12624 10260
rect 12579 10220 12624 10248
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13630 10248 13636 10260
rect 13591 10220 13636 10248
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 14918 10208 14924 10260
rect 14976 10248 14982 10260
rect 15013 10251 15071 10257
rect 15013 10248 15025 10251
rect 14976 10220 15025 10248
rect 14976 10208 14982 10220
rect 15013 10217 15025 10220
rect 15059 10217 15071 10251
rect 15013 10211 15071 10217
rect 15841 10251 15899 10257
rect 15841 10217 15853 10251
rect 15887 10248 15899 10251
rect 16114 10248 16120 10260
rect 15887 10220 16120 10248
rect 15887 10217 15899 10220
rect 15841 10211 15899 10217
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 20438 10248 20444 10260
rect 20399 10220 20444 10248
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 22002 10248 22008 10260
rect 21963 10220 22008 10248
rect 22002 10208 22008 10220
rect 22060 10208 22066 10260
rect 10505 10183 10563 10189
rect 10505 10180 10517 10183
rect 10100 10152 10517 10180
rect 10100 10140 10106 10152
rect 10505 10149 10517 10152
rect 10551 10149 10563 10183
rect 10505 10143 10563 10149
rect 11333 10183 11391 10189
rect 11333 10149 11345 10183
rect 11379 10149 11391 10183
rect 11882 10180 11888 10192
rect 11843 10152 11888 10180
rect 11333 10143 11391 10149
rect 11882 10140 11888 10152
rect 11940 10140 11946 10192
rect 13078 10189 13084 10192
rect 13075 10180 13084 10189
rect 13039 10152 13084 10180
rect 13075 10143 13084 10152
rect 13078 10140 13084 10143
rect 13136 10140 13142 10192
rect 13354 10140 13360 10192
rect 13412 10180 13418 10192
rect 13909 10183 13967 10189
rect 13909 10180 13921 10183
rect 13412 10152 13921 10180
rect 13412 10140 13418 10152
rect 13909 10149 13921 10152
rect 13955 10149 13967 10183
rect 13909 10143 13967 10149
rect 2130 10072 2136 10124
rect 2188 10112 2194 10124
rect 2409 10115 2467 10121
rect 2409 10112 2421 10115
rect 2188 10084 2421 10112
rect 2188 10072 2194 10084
rect 2409 10081 2421 10084
rect 2455 10081 2467 10115
rect 2409 10075 2467 10081
rect 2424 10044 2452 10075
rect 2590 10072 2596 10124
rect 2648 10112 2654 10124
rect 2685 10115 2743 10121
rect 2685 10112 2697 10115
rect 2648 10084 2697 10112
rect 2648 10072 2654 10084
rect 2685 10081 2697 10084
rect 2731 10081 2743 10115
rect 3142 10112 3148 10124
rect 3103 10084 3148 10112
rect 2685 10075 2743 10081
rect 3142 10072 3148 10084
rect 3200 10072 3206 10124
rect 4890 10072 4896 10124
rect 4948 10112 4954 10124
rect 4985 10115 5043 10121
rect 4985 10112 4997 10115
rect 4948 10084 4997 10112
rect 4948 10072 4954 10084
rect 4985 10081 4997 10084
rect 5031 10081 5043 10115
rect 4985 10075 5043 10081
rect 5261 10115 5319 10121
rect 5261 10081 5273 10115
rect 5307 10112 5319 10115
rect 5350 10112 5356 10124
rect 5307 10084 5356 10112
rect 5307 10081 5319 10084
rect 5261 10075 5319 10081
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 6549 10115 6607 10121
rect 6549 10081 6561 10115
rect 6595 10112 6607 10115
rect 6638 10112 6644 10124
rect 6595 10084 6644 10112
rect 6595 10081 6607 10084
rect 6549 10075 6607 10081
rect 6638 10072 6644 10084
rect 6696 10112 6702 10124
rect 7282 10112 7288 10124
rect 6696 10084 7288 10112
rect 6696 10072 6702 10084
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 9674 10112 9680 10124
rect 9635 10084 9680 10112
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 9858 10072 9864 10124
rect 9916 10112 9922 10124
rect 10137 10115 10195 10121
rect 10137 10112 10149 10115
rect 9916 10084 10149 10112
rect 9916 10072 9922 10084
rect 10137 10081 10149 10084
rect 10183 10081 10195 10115
rect 10137 10075 10195 10081
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 12713 10115 12771 10121
rect 12713 10112 12725 10115
rect 12492 10084 12725 10112
rect 12492 10072 12498 10084
rect 12713 10081 12725 10084
rect 12759 10112 12771 10115
rect 13262 10112 13268 10124
rect 12759 10084 13268 10112
rect 12759 10081 12771 10084
rect 12713 10075 12771 10081
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13924 10112 13952 10143
rect 13998 10140 14004 10192
rect 14056 10180 14062 10192
rect 15746 10180 15752 10192
rect 14056 10152 15752 10180
rect 14056 10140 14062 10152
rect 15746 10140 15752 10152
rect 15804 10180 15810 10192
rect 16209 10183 16267 10189
rect 16209 10180 16221 10183
rect 15804 10152 16221 10180
rect 15804 10140 15810 10152
rect 16209 10149 16221 10152
rect 16255 10149 16267 10183
rect 16209 10143 16267 10149
rect 16942 10140 16948 10192
rect 17000 10180 17006 10192
rect 17310 10180 17316 10192
rect 17000 10152 17316 10180
rect 17000 10140 17006 10152
rect 17310 10140 17316 10152
rect 17368 10180 17374 10192
rect 17368 10152 17632 10180
rect 17368 10140 17374 10152
rect 16390 10112 16396 10124
rect 13924 10084 16396 10112
rect 16390 10072 16396 10084
rect 16448 10072 16454 10124
rect 16574 10072 16580 10124
rect 16632 10112 16638 10124
rect 16853 10115 16911 10121
rect 16853 10112 16865 10115
rect 16632 10084 16865 10112
rect 16632 10072 16638 10084
rect 16853 10081 16865 10084
rect 16899 10081 16911 10115
rect 17218 10112 17224 10124
rect 17179 10084 17224 10112
rect 16853 10075 16911 10081
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 17604 10121 17632 10152
rect 18874 10140 18880 10192
rect 18932 10180 18938 10192
rect 19014 10183 19072 10189
rect 19014 10180 19026 10183
rect 18932 10152 19026 10180
rect 18932 10140 18938 10152
rect 19014 10149 19026 10152
rect 19060 10149 19072 10183
rect 19014 10143 19072 10149
rect 20806 10140 20812 10192
rect 20864 10180 20870 10192
rect 21085 10183 21143 10189
rect 21085 10180 21097 10183
rect 20864 10152 21097 10180
rect 20864 10140 20870 10152
rect 21085 10149 21097 10152
rect 21131 10149 21143 10183
rect 21085 10143 21143 10149
rect 17589 10115 17647 10121
rect 17589 10081 17601 10115
rect 17635 10081 17647 10115
rect 17589 10075 17647 10081
rect 18046 10072 18052 10124
rect 18104 10112 18110 10124
rect 18598 10112 18604 10124
rect 18104 10084 18604 10112
rect 18104 10072 18110 10084
rect 18598 10072 18604 10084
rect 18656 10112 18662 10124
rect 18693 10115 18751 10121
rect 18693 10112 18705 10115
rect 18656 10084 18705 10112
rect 18656 10072 18662 10084
rect 18693 10081 18705 10084
rect 18739 10081 18751 10115
rect 18693 10075 18751 10081
rect 22094 10072 22100 10124
rect 22152 10112 22158 10124
rect 23106 10112 23112 10124
rect 23164 10121 23170 10124
rect 23164 10115 23202 10121
rect 22152 10084 23112 10112
rect 22152 10072 22158 10084
rect 23106 10072 23112 10084
rect 23190 10081 23202 10115
rect 23164 10075 23202 10081
rect 23164 10072 23170 10075
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 2424 10016 4537 10044
rect 4525 10013 4537 10016
rect 4571 10044 4583 10047
rect 5166 10044 5172 10056
rect 4571 10016 5172 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 8352 10016 8401 10044
rect 8352 10004 8358 10016
rect 8389 10013 8401 10016
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 11241 10047 11299 10053
rect 11241 10013 11253 10047
rect 11287 10044 11299 10047
rect 11514 10044 11520 10056
rect 11287 10016 11520 10044
rect 11287 10013 11299 10016
rect 11241 10007 11299 10013
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 15286 10044 15292 10056
rect 15247 10016 15292 10044
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 17865 10047 17923 10053
rect 17865 10013 17877 10047
rect 17911 10044 17923 10047
rect 17954 10044 17960 10056
rect 17911 10016 17960 10044
rect 17911 10013 17923 10016
rect 17865 10007 17923 10013
rect 17954 10004 17960 10016
rect 18012 10004 18018 10056
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 20993 10047 21051 10053
rect 20993 10044 21005 10047
rect 20772 10016 21005 10044
rect 20772 10004 20778 10016
rect 20993 10013 21005 10016
rect 21039 10013 21051 10047
rect 20993 10007 21051 10013
rect 21637 10047 21695 10053
rect 21637 10013 21649 10047
rect 21683 10044 21695 10047
rect 21726 10044 21732 10056
rect 21683 10016 21732 10044
rect 21683 10013 21695 10016
rect 21637 10007 21695 10013
rect 21726 10004 21732 10016
rect 21784 10004 21790 10056
rect 2498 9976 2504 9988
rect 2459 9948 2504 9976
rect 2498 9936 2504 9948
rect 2556 9936 2562 9988
rect 4982 9936 4988 9988
rect 5040 9976 5046 9988
rect 5077 9979 5135 9985
rect 5077 9976 5089 9979
rect 5040 9948 5089 9976
rect 5040 9936 5046 9948
rect 5077 9945 5089 9948
rect 5123 9945 5135 9979
rect 5077 9939 5135 9945
rect 6270 9936 6276 9988
rect 6328 9976 6334 9988
rect 6733 9979 6791 9985
rect 6733 9976 6745 9979
rect 6328 9948 6745 9976
rect 6328 9936 6334 9948
rect 6733 9945 6745 9948
rect 6779 9945 6791 9979
rect 6733 9939 6791 9945
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7009 9911 7067 9917
rect 7009 9908 7021 9911
rect 6972 9880 7021 9908
rect 6972 9868 6978 9880
rect 7009 9877 7021 9880
rect 7055 9877 7067 9911
rect 7009 9871 7067 9877
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9908 7527 9911
rect 7558 9908 7564 9920
rect 7515 9880 7564 9908
rect 7515 9877 7527 9880
rect 7469 9871 7527 9877
rect 7558 9868 7564 9880
rect 7616 9868 7622 9920
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 9033 9911 9091 9917
rect 9033 9908 9045 9911
rect 8536 9880 9045 9908
rect 8536 9868 8542 9880
rect 9033 9877 9045 9880
rect 9079 9877 9091 9911
rect 9858 9908 9864 9920
rect 9819 9880 9864 9908
rect 9033 9871 9091 9877
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 12158 9908 12164 9920
rect 12119 9880 12164 9908
rect 12158 9868 12164 9880
rect 12216 9908 12222 9920
rect 13538 9908 13544 9920
rect 12216 9880 13544 9908
rect 12216 9868 12222 9880
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 19613 9911 19671 9917
rect 19613 9877 19625 9911
rect 19659 9908 19671 9911
rect 20806 9908 20812 9920
rect 19659 9880 20812 9908
rect 19659 9877 19671 9880
rect 19613 9871 19671 9877
rect 20806 9868 20812 9880
rect 20864 9868 20870 9920
rect 23247 9911 23305 9917
rect 23247 9877 23259 9911
rect 23293 9908 23305 9911
rect 23382 9908 23388 9920
rect 23293 9880 23388 9908
rect 23293 9877 23305 9880
rect 23247 9871 23305 9877
rect 23382 9868 23388 9880
rect 23440 9868 23446 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2130 9704 2136 9716
rect 2091 9676 2136 9704
rect 2130 9664 2136 9676
rect 2188 9664 2194 9716
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 5074 9704 5080 9716
rect 2556 9676 2820 9704
rect 2556 9664 2562 9676
rect 2792 9636 2820 9676
rect 4080 9676 5080 9704
rect 2869 9639 2927 9645
rect 2869 9636 2881 9639
rect 2792 9608 2881 9636
rect 2869 9605 2881 9608
rect 2915 9636 2927 9639
rect 3973 9639 4031 9645
rect 3973 9636 3985 9639
rect 2915 9608 3985 9636
rect 2915 9605 2927 9608
rect 2869 9599 2927 9605
rect 3973 9605 3985 9608
rect 4019 9636 4031 9639
rect 4080 9636 4108 9676
rect 5074 9664 5080 9676
rect 5132 9664 5138 9716
rect 6638 9704 6644 9716
rect 6599 9676 6644 9704
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 6914 9664 6920 9716
rect 6972 9664 6978 9716
rect 8110 9664 8116 9716
rect 8168 9704 8174 9716
rect 8168 9676 8248 9704
rect 8168 9664 8174 9676
rect 6932 9636 6960 9664
rect 4019 9608 4108 9636
rect 5184 9608 6960 9636
rect 8220 9636 8248 9676
rect 9674 9664 9680 9716
rect 9732 9704 9738 9716
rect 9769 9707 9827 9713
rect 9769 9704 9781 9707
rect 9732 9676 9781 9704
rect 9732 9664 9738 9676
rect 9769 9673 9781 9676
rect 9815 9673 9827 9707
rect 9769 9667 9827 9673
rect 11885 9707 11943 9713
rect 11885 9673 11897 9707
rect 11931 9704 11943 9707
rect 12066 9704 12072 9716
rect 11931 9676 12072 9704
rect 11931 9673 11943 9676
rect 11885 9667 11943 9673
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 15286 9704 15292 9716
rect 15120 9676 15292 9704
rect 9125 9639 9183 9645
rect 9125 9636 9137 9639
rect 8220 9608 9137 9636
rect 4019 9605 4031 9608
rect 3973 9599 4031 9605
rect 3326 9568 3332 9580
rect 3287 9540 3332 9568
rect 3326 9528 3332 9540
rect 3384 9568 3390 9580
rect 4982 9568 4988 9580
rect 3384 9540 3648 9568
rect 3384 9528 3390 9540
rect 3620 9509 3648 9540
rect 4540 9540 4988 9568
rect 4540 9509 4568 9540
rect 4982 9528 4988 9540
rect 5040 9568 5046 9580
rect 5184 9577 5212 9608
rect 9125 9605 9137 9608
rect 9171 9605 9183 9639
rect 9125 9599 9183 9605
rect 9398 9596 9404 9648
rect 9456 9636 9462 9648
rect 9493 9639 9551 9645
rect 9493 9636 9505 9639
rect 9456 9608 9505 9636
rect 9456 9596 9462 9608
rect 9493 9605 9505 9608
rect 9539 9605 9551 9639
rect 9493 9599 9551 9605
rect 10689 9639 10747 9645
rect 10689 9605 10701 9639
rect 10735 9636 10747 9639
rect 10962 9636 10968 9648
rect 10735 9608 10968 9636
rect 10735 9605 10747 9608
rect 10689 9599 10747 9605
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 13814 9636 13820 9648
rect 13775 9608 13820 9636
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14642 9636 14648 9648
rect 14603 9608 14648 9636
rect 14642 9596 14648 9608
rect 14700 9596 14706 9648
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 5040 9540 5181 9568
rect 5040 9528 5046 9540
rect 5169 9537 5181 9540
rect 5215 9537 5227 9571
rect 5534 9568 5540 9580
rect 5495 9540 5540 9568
rect 5169 9531 5227 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 12526 9568 12532 9580
rect 12487 9540 12532 9568
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12986 9568 12992 9580
rect 12947 9540 12992 9568
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 14093 9571 14151 9577
rect 14093 9537 14105 9571
rect 14139 9568 14151 9571
rect 14366 9568 14372 9580
rect 14139 9540 14372 9568
rect 14139 9537 14151 9540
rect 14093 9531 14151 9537
rect 14366 9528 14372 9540
rect 14424 9568 14430 9580
rect 15120 9568 15148 9676
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 15470 9704 15476 9716
rect 15431 9676 15476 9704
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 17310 9704 17316 9716
rect 17271 9676 17316 9704
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 18966 9704 18972 9716
rect 18927 9676 18972 9704
rect 18966 9664 18972 9676
rect 19024 9664 19030 9716
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 23106 9704 23112 9716
rect 20772 9676 22048 9704
rect 23067 9676 23112 9704
rect 20772 9664 20778 9676
rect 15841 9639 15899 9645
rect 15841 9605 15853 9639
rect 15887 9636 15899 9639
rect 16482 9636 16488 9648
rect 15887 9608 16488 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 16482 9596 16488 9608
rect 16540 9596 16546 9648
rect 17037 9639 17095 9645
rect 17037 9605 17049 9639
rect 17083 9636 17095 9639
rect 17218 9636 17224 9648
rect 17083 9608 17224 9636
rect 17083 9605 17095 9608
rect 17037 9599 17095 9605
rect 17218 9596 17224 9608
rect 17276 9596 17282 9648
rect 18984 9636 19012 9664
rect 19613 9639 19671 9645
rect 19613 9636 19625 9639
rect 18984 9608 19625 9636
rect 19613 9605 19625 9608
rect 19659 9636 19671 9639
rect 19978 9636 19984 9648
rect 19659 9608 19984 9636
rect 19659 9605 19671 9608
rect 19613 9599 19671 9605
rect 19978 9596 19984 9608
rect 20036 9596 20042 9648
rect 20806 9636 20812 9648
rect 20767 9608 20812 9636
rect 20806 9596 20812 9608
rect 20864 9596 20870 9648
rect 22020 9636 22048 9676
rect 23106 9664 23112 9676
rect 23164 9664 23170 9716
rect 22373 9639 22431 9645
rect 22373 9636 22385 9639
rect 22020 9608 22385 9636
rect 22373 9605 22385 9608
rect 22419 9605 22431 9639
rect 24762 9636 24768 9648
rect 24723 9608 24768 9636
rect 22373 9599 22431 9605
rect 24762 9596 24768 9608
rect 24820 9596 24826 9648
rect 14424 9540 15148 9568
rect 14424 9528 14430 9540
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18049 9571 18107 9577
rect 18049 9568 18061 9571
rect 18012 9540 18061 9568
rect 18012 9528 18018 9540
rect 18049 9537 18061 9540
rect 18095 9537 18107 9571
rect 18049 9531 18107 9537
rect 18874 9528 18880 9580
rect 18932 9568 18938 9580
rect 19245 9571 19303 9577
rect 19245 9568 19257 9571
rect 18932 9540 19257 9568
rect 18932 9528 18938 9540
rect 19245 9537 19257 9540
rect 19291 9537 19303 9571
rect 20162 9568 20168 9580
rect 20123 9540 20168 9568
rect 19245 9531 19303 9537
rect 20162 9528 20168 9540
rect 20220 9568 20226 9580
rect 20714 9568 20720 9580
rect 20220 9540 20720 9568
rect 20220 9528 20226 9540
rect 20714 9528 20720 9540
rect 20772 9528 20778 9580
rect 21266 9528 21272 9580
rect 21324 9568 21330 9580
rect 21453 9571 21511 9577
rect 21453 9568 21465 9571
rect 21324 9540 21465 9568
rect 21324 9528 21330 9540
rect 21453 9537 21465 9540
rect 21499 9537 21511 9571
rect 21726 9568 21732 9580
rect 21687 9540 21732 9568
rect 21453 9531 21511 9537
rect 21726 9528 21732 9540
rect 21784 9528 21790 9580
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 4525 9503 4583 9509
rect 4525 9500 4537 9503
rect 3651 9472 4537 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 4525 9469 4537 9472
rect 4571 9469 4583 9503
rect 5074 9500 5080 9512
rect 5035 9472 5080 9500
rect 4525 9463 4583 9469
rect 5074 9460 5080 9472
rect 5132 9460 5138 9512
rect 5350 9500 5356 9512
rect 5311 9472 5356 9500
rect 5350 9460 5356 9472
rect 5408 9500 5414 9512
rect 6089 9503 6147 9509
rect 6089 9500 6101 9503
rect 5408 9472 6101 9500
rect 5408 9460 5414 9472
rect 6089 9469 6101 9472
rect 6135 9469 6147 9503
rect 7561 9503 7619 9509
rect 7561 9500 7573 9503
rect 6089 9463 6147 9469
rect 7024 9472 7573 9500
rect 7024 9376 7052 9472
rect 7561 9469 7573 9472
rect 7607 9469 7619 9503
rect 9306 9500 9312 9512
rect 9267 9472 9312 9500
rect 7561 9463 7619 9469
rect 9306 9460 9312 9472
rect 9364 9500 9370 9512
rect 10137 9503 10195 9509
rect 10137 9500 10149 9503
rect 9364 9472 10149 9500
rect 9364 9460 9370 9472
rect 10137 9469 10149 9472
rect 10183 9469 10195 9503
rect 10137 9463 10195 9469
rect 7923 9435 7981 9441
rect 7923 9401 7935 9435
rect 7969 9401 7981 9435
rect 10873 9435 10931 9441
rect 10873 9432 10885 9435
rect 7923 9395 7981 9401
rect 10796 9404 10885 9432
rect 2501 9367 2559 9373
rect 2501 9333 2513 9367
rect 2547 9364 2559 9367
rect 2590 9364 2596 9376
rect 2547 9336 2596 9364
rect 2547 9333 2559 9336
rect 2501 9327 2559 9333
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 4890 9364 4896 9376
rect 4851 9336 4896 9364
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 7006 9364 7012 9376
rect 6967 9336 7012 9364
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 7469 9367 7527 9373
rect 7469 9333 7481 9367
rect 7515 9364 7527 9367
rect 7944 9364 7972 9395
rect 10796 9376 10824 9404
rect 10873 9401 10885 9404
rect 10919 9401 10931 9435
rect 10873 9395 10931 9401
rect 10962 9392 10968 9444
rect 11020 9432 11026 9444
rect 11514 9432 11520 9444
rect 11020 9404 11065 9432
rect 11475 9404 11520 9432
rect 11020 9392 11026 9404
rect 11514 9392 11520 9404
rect 11572 9392 11578 9444
rect 12621 9435 12679 9441
rect 12621 9401 12633 9435
rect 12667 9401 12679 9435
rect 12621 9395 12679 9401
rect 8110 9364 8116 9376
rect 7515 9336 8116 9364
rect 7515 9333 7527 9336
rect 7469 9327 7527 9333
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 8478 9364 8484 9376
rect 8439 9336 8484 9364
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 8754 9364 8760 9376
rect 8715 9336 8760 9364
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 10778 9324 10784 9376
rect 10836 9324 10842 9376
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 12250 9364 12256 9376
rect 11388 9336 12256 9364
rect 11388 9324 11394 9336
rect 12250 9324 12256 9336
rect 12308 9364 12314 9376
rect 12636 9364 12664 9395
rect 13814 9392 13820 9444
rect 13872 9432 13878 9444
rect 14185 9435 14243 9441
rect 14185 9432 14197 9435
rect 13872 9404 14197 9432
rect 13872 9392 13878 9404
rect 14185 9401 14197 9404
rect 14231 9401 14243 9435
rect 14185 9395 14243 9401
rect 15105 9435 15163 9441
rect 15105 9401 15117 9435
rect 15151 9432 15163 9435
rect 16022 9432 16028 9444
rect 15151 9404 15884 9432
rect 15983 9404 16028 9432
rect 15151 9401 15163 9404
rect 15105 9395 15163 9401
rect 12308 9336 12664 9364
rect 12308 9324 12314 9336
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 13541 9367 13599 9373
rect 13541 9364 13553 9367
rect 13136 9336 13553 9364
rect 13136 9324 13142 9336
rect 13541 9333 13553 9336
rect 13587 9364 13599 9367
rect 13722 9364 13728 9376
rect 13587 9336 13728 9364
rect 13587 9333 13599 9336
rect 13541 9327 13599 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 15856 9364 15884 9404
rect 16022 9392 16028 9404
rect 16080 9392 16086 9444
rect 16117 9435 16175 9441
rect 16117 9401 16129 9435
rect 16163 9401 16175 9435
rect 16666 9432 16672 9444
rect 16627 9404 16672 9432
rect 16117 9395 16175 9401
rect 16132 9364 16160 9395
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 17862 9432 17868 9444
rect 17775 9404 17868 9432
rect 17862 9392 17868 9404
rect 17920 9432 17926 9444
rect 18411 9435 18469 9441
rect 18411 9432 18423 9435
rect 17920 9404 18423 9432
rect 17920 9392 17926 9404
rect 18411 9401 18423 9404
rect 18457 9432 18469 9435
rect 18892 9432 18920 9528
rect 24578 9500 24584 9512
rect 24491 9472 24584 9500
rect 24578 9460 24584 9472
rect 24636 9500 24642 9512
rect 25133 9503 25191 9509
rect 25133 9500 25145 9503
rect 24636 9472 25145 9500
rect 24636 9460 24642 9472
rect 25133 9469 25145 9472
rect 25179 9469 25191 9503
rect 25133 9463 25191 9469
rect 18457 9404 18920 9432
rect 18457 9401 18469 9404
rect 18411 9395 18469 9401
rect 19518 9392 19524 9444
rect 19576 9432 19582 9444
rect 19889 9435 19947 9441
rect 19889 9432 19901 9435
rect 19576 9404 19901 9432
rect 19576 9392 19582 9404
rect 19889 9401 19901 9404
rect 19935 9401 19947 9435
rect 19889 9395 19947 9401
rect 19978 9392 19984 9444
rect 20036 9432 20042 9444
rect 20036 9404 20081 9432
rect 20036 9392 20042 9404
rect 21542 9392 21548 9444
rect 21600 9432 21606 9444
rect 21600 9404 21645 9432
rect 21600 9392 21606 9404
rect 16206 9364 16212 9376
rect 15856 9336 16212 9364
rect 16206 9324 16212 9336
rect 16264 9324 16270 9376
rect 21269 9367 21327 9373
rect 21269 9333 21281 9367
rect 21315 9364 21327 9367
rect 21560 9364 21588 9392
rect 21315 9336 21588 9364
rect 21315 9333 21327 9336
rect 21269 9327 21327 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 4982 9120 4988 9172
rect 5040 9160 5046 9172
rect 5537 9163 5595 9169
rect 5537 9160 5549 9163
rect 5040 9132 5549 9160
rect 5040 9120 5046 9132
rect 5537 9129 5549 9132
rect 5583 9129 5595 9163
rect 5537 9123 5595 9129
rect 6273 9163 6331 9169
rect 6273 9129 6285 9163
rect 6319 9160 6331 9163
rect 7193 9163 7251 9169
rect 7193 9160 7205 9163
rect 6319 9132 7205 9160
rect 6319 9129 6331 9132
rect 6273 9123 6331 9129
rect 7193 9129 7205 9132
rect 7239 9160 7251 9163
rect 7374 9160 7380 9172
rect 7239 9132 7380 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 7374 9120 7380 9132
rect 7432 9160 7438 9172
rect 7742 9160 7748 9172
rect 7432 9132 7748 9160
rect 7432 9120 7438 9132
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 8481 9163 8539 9169
rect 8481 9160 8493 9163
rect 8260 9132 8493 9160
rect 8260 9120 8266 9132
rect 8481 9129 8493 9132
rect 8527 9160 8539 9163
rect 8570 9160 8576 9172
rect 8527 9132 8576 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 8570 9120 8576 9132
rect 8628 9160 8634 9172
rect 8754 9160 8760 9172
rect 8628 9132 8760 9160
rect 8628 9120 8634 9132
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 11330 9160 11336 9172
rect 11291 9132 11336 9160
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 13262 9160 13268 9172
rect 13223 9132 13268 9160
rect 13262 9120 13268 9132
rect 13320 9120 13326 9172
rect 13998 9160 14004 9172
rect 13959 9132 14004 9160
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14366 9160 14372 9172
rect 14327 9132 14372 9160
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 15105 9163 15163 9169
rect 15105 9129 15117 9163
rect 15151 9160 15163 9163
rect 16022 9160 16028 9172
rect 15151 9132 16028 9160
rect 15151 9129 15163 9132
rect 15105 9123 15163 9129
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 16206 9160 16212 9172
rect 16167 9132 16212 9160
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 16574 9160 16580 9172
rect 16535 9132 16580 9160
rect 16574 9120 16580 9132
rect 16632 9120 16638 9172
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 18012 9132 18061 9160
rect 18012 9120 18018 9132
rect 18049 9129 18061 9132
rect 18095 9129 18107 9163
rect 18598 9160 18604 9172
rect 18559 9132 18604 9160
rect 18049 9123 18107 9129
rect 18598 9120 18604 9132
rect 18656 9120 18662 9172
rect 23707 9163 23765 9169
rect 23707 9129 23719 9163
rect 23753 9160 23765 9163
rect 24578 9160 24584 9172
rect 23753 9132 24584 9160
rect 23753 9129 23765 9132
rect 23707 9123 23765 9129
rect 24578 9120 24584 9132
rect 24636 9120 24642 9172
rect 5261 9095 5319 9101
rect 5261 9061 5273 9095
rect 5307 9092 5319 9095
rect 5350 9092 5356 9104
rect 5307 9064 5356 9092
rect 5307 9061 5319 9064
rect 5261 9055 5319 9061
rect 5350 9052 5356 9064
rect 5408 9092 5414 9104
rect 5905 9095 5963 9101
rect 5905 9092 5917 9095
rect 5408 9064 5917 9092
rect 5408 9052 5414 9064
rect 5905 9061 5917 9064
rect 5951 9061 5963 9095
rect 5905 9055 5963 9061
rect 7923 9095 7981 9101
rect 7923 9061 7935 9095
rect 7969 9092 7981 9095
rect 8110 9092 8116 9104
rect 7969 9064 8116 9092
rect 7969 9061 7981 9064
rect 7923 9055 7981 9061
rect 8110 9052 8116 9064
rect 8168 9052 8174 9104
rect 8386 9052 8392 9104
rect 8444 9092 8450 9104
rect 8849 9095 8907 9101
rect 8849 9092 8861 9095
rect 8444 9064 8861 9092
rect 8444 9052 8450 9064
rect 8849 9061 8861 9064
rect 8895 9092 8907 9095
rect 9306 9092 9312 9104
rect 8895 9064 9312 9092
rect 8895 9061 8907 9064
rect 8849 9055 8907 9061
rect 9306 9052 9312 9064
rect 9364 9052 9370 9104
rect 10134 9052 10140 9104
rect 10192 9092 10198 9104
rect 10734 9095 10792 9101
rect 10734 9092 10746 9095
rect 10192 9064 10746 9092
rect 10192 9052 10198 9064
rect 10734 9061 10746 9064
rect 10780 9061 10792 9095
rect 10734 9055 10792 9061
rect 12158 9052 12164 9104
rect 12216 9092 12222 9104
rect 12437 9095 12495 9101
rect 12437 9092 12449 9095
rect 12216 9064 12449 9092
rect 12216 9052 12222 9064
rect 12437 9061 12449 9064
rect 12483 9061 12495 9095
rect 12986 9092 12992 9104
rect 12947 9064 12992 9092
rect 12437 9055 12495 9061
rect 12986 9052 12992 9064
rect 13044 9052 13050 9104
rect 15378 9052 15384 9104
rect 15436 9092 15442 9104
rect 15651 9095 15709 9101
rect 15651 9092 15663 9095
rect 15436 9064 15663 9092
rect 15436 9052 15442 9064
rect 15651 9061 15663 9064
rect 15697 9092 15709 9095
rect 15697 9064 16160 9092
rect 15697 9061 15709 9064
rect 15651 9055 15709 9061
rect 4614 9024 4620 9036
rect 4575 8996 4620 9024
rect 4614 8984 4620 8996
rect 4672 9024 4678 9036
rect 5166 9024 5172 9036
rect 4672 8996 5172 9024
rect 4672 8984 4678 8996
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 6086 9024 6092 9036
rect 6047 8996 6092 9024
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 10321 9027 10379 9033
rect 10321 8993 10333 9027
rect 10367 9024 10379 9027
rect 11514 9024 11520 9036
rect 10367 8996 11520 9024
rect 10367 8993 10379 8996
rect 10321 8987 10379 8993
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 13538 8984 13544 9036
rect 13596 9024 13602 9036
rect 13817 9027 13875 9033
rect 13817 9024 13829 9027
rect 13596 8996 13829 9024
rect 13596 8984 13602 8996
rect 13817 8993 13829 8996
rect 13863 8993 13875 9027
rect 13817 8987 13875 8993
rect 14826 8984 14832 9036
rect 14884 9024 14890 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 14884 8996 15301 9024
rect 14884 8984 14890 8996
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 7561 8959 7619 8965
rect 7561 8925 7573 8959
rect 7607 8956 7619 8959
rect 7834 8956 7840 8968
rect 7607 8928 7840 8956
rect 7607 8925 7619 8928
rect 7561 8919 7619 8925
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 10042 8916 10048 8968
rect 10100 8956 10106 8968
rect 10413 8959 10471 8965
rect 10413 8956 10425 8959
rect 10100 8928 10425 8956
rect 10100 8916 10106 8928
rect 10413 8925 10425 8928
rect 10459 8925 10471 8959
rect 12342 8956 12348 8968
rect 12303 8928 12348 8956
rect 10413 8919 10471 8925
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 10778 8848 10784 8900
rect 10836 8888 10842 8900
rect 11609 8891 11667 8897
rect 11609 8888 11621 8891
rect 10836 8860 11621 8888
rect 10836 8848 10842 8860
rect 11609 8857 11621 8860
rect 11655 8857 11667 8891
rect 11609 8851 11667 8857
rect 12161 8891 12219 8897
rect 12161 8857 12173 8891
rect 12207 8888 12219 8891
rect 12526 8888 12532 8900
rect 12207 8860 12532 8888
rect 12207 8857 12219 8860
rect 12161 8851 12219 8857
rect 12526 8848 12532 8860
rect 12584 8848 12590 8900
rect 16132 8888 16160 9064
rect 16224 9024 16252 9120
rect 18506 9052 18512 9104
rect 18564 9092 18570 9104
rect 18877 9095 18935 9101
rect 18877 9092 18889 9095
rect 18564 9064 18889 9092
rect 18564 9052 18570 9064
rect 18877 9061 18889 9064
rect 18923 9061 18935 9095
rect 18877 9055 18935 9061
rect 18969 9095 19027 9101
rect 18969 9061 18981 9095
rect 19015 9092 19027 9095
rect 19058 9092 19064 9104
rect 19015 9064 19064 9092
rect 19015 9061 19027 9064
rect 18969 9055 19027 9061
rect 19058 9052 19064 9064
rect 19116 9052 19122 9104
rect 19521 9095 19579 9101
rect 19521 9061 19533 9095
rect 19567 9092 19579 9095
rect 20162 9092 20168 9104
rect 19567 9064 20168 9092
rect 19567 9061 19579 9064
rect 19521 9055 19579 9061
rect 20162 9052 20168 9064
rect 20220 9052 20226 9104
rect 21082 9092 21088 9104
rect 21043 9064 21088 9092
rect 21082 9052 21088 9064
rect 21140 9052 21146 9104
rect 17126 9024 17132 9036
rect 16224 8996 17132 9024
rect 17126 8984 17132 8996
rect 17184 8984 17190 9036
rect 23566 8984 23572 9036
rect 23624 9033 23630 9036
rect 23624 9027 23662 9033
rect 23650 8993 23662 9027
rect 23624 8987 23662 8993
rect 23624 8984 23630 8987
rect 16206 8916 16212 8968
rect 16264 8956 16270 8968
rect 17037 8959 17095 8965
rect 17037 8956 17049 8959
rect 16264 8928 17049 8956
rect 16264 8916 16270 8928
rect 17037 8925 17049 8928
rect 17083 8925 17095 8959
rect 20990 8956 20996 8968
rect 20951 8928 20996 8956
rect 17037 8919 17095 8925
rect 20990 8916 20996 8928
rect 21048 8916 21054 8968
rect 21266 8956 21272 8968
rect 21227 8928 21272 8956
rect 21266 8916 21272 8928
rect 21324 8956 21330 8968
rect 21913 8959 21971 8965
rect 21913 8956 21925 8959
rect 21324 8928 21925 8956
rect 21324 8916 21330 8928
rect 21913 8925 21925 8928
rect 21959 8925 21971 8959
rect 21913 8919 21971 8925
rect 17862 8888 17868 8900
rect 16132 8860 17868 8888
rect 17862 8848 17868 8860
rect 17920 8848 17926 8900
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 19797 8823 19855 8829
rect 19797 8820 19809 8823
rect 19576 8792 19809 8820
rect 19576 8780 19582 8792
rect 19797 8789 19809 8792
rect 19843 8789 19855 8823
rect 19797 8783 19855 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 4065 8619 4123 8625
rect 4065 8616 4077 8619
rect 2648 8588 4077 8616
rect 2648 8576 2654 8588
rect 4065 8585 4077 8588
rect 4111 8616 4123 8619
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 4111 8588 4445 8616
rect 4111 8585 4123 8588
rect 4065 8579 4123 8585
rect 4433 8585 4445 8588
rect 4479 8616 4491 8619
rect 4614 8616 4620 8628
rect 4479 8588 4620 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 8662 8616 8668 8628
rect 8623 8588 8668 8616
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 13538 8616 13544 8628
rect 13403 8588 13544 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 13722 8576 13728 8628
rect 13780 8616 13786 8628
rect 15378 8616 15384 8628
rect 13780 8588 15384 8616
rect 13780 8576 13786 8588
rect 4632 8480 4660 8576
rect 4982 8508 4988 8560
rect 5040 8548 5046 8560
rect 5077 8551 5135 8557
rect 5077 8548 5089 8551
rect 5040 8520 5089 8548
rect 5040 8508 5046 8520
rect 5077 8517 5089 8520
rect 5123 8548 5135 8551
rect 5997 8551 6055 8557
rect 5997 8548 6009 8551
rect 5123 8520 6009 8548
rect 5123 8517 5135 8520
rect 5077 8511 5135 8517
rect 5997 8517 6009 8520
rect 6043 8517 6055 8551
rect 10134 8548 10140 8560
rect 5997 8511 6055 8517
rect 9876 8520 10140 8548
rect 5721 8483 5779 8489
rect 4632 8452 5120 8480
rect 4154 8372 4160 8424
rect 4212 8412 4218 8424
rect 4801 8415 4859 8421
rect 4801 8412 4813 8415
rect 4212 8384 4813 8412
rect 4212 8372 4218 8384
rect 4801 8381 4813 8384
rect 4847 8412 4859 8415
rect 4890 8412 4896 8424
rect 4847 8384 4896 8412
rect 4847 8381 4859 8384
rect 4801 8375 4859 8381
rect 4890 8372 4896 8384
rect 4948 8412 4954 8424
rect 4985 8415 5043 8421
rect 4985 8412 4997 8415
rect 4948 8384 4997 8412
rect 4948 8372 4954 8384
rect 4985 8381 4997 8384
rect 5031 8381 5043 8415
rect 5092 8412 5120 8452
rect 5721 8449 5733 8483
rect 5767 8480 5779 8483
rect 6086 8480 6092 8492
rect 5767 8452 6092 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 6086 8440 6092 8452
rect 6144 8480 6150 8492
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 6144 8452 6377 8480
rect 6144 8440 6150 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 8110 8440 8116 8492
rect 8168 8480 8174 8492
rect 9876 8489 9904 8520
rect 10134 8508 10140 8520
rect 10192 8548 10198 8560
rect 10229 8551 10287 8557
rect 10229 8548 10241 8551
rect 10192 8520 10241 8548
rect 10192 8508 10198 8520
rect 10229 8517 10241 8520
rect 10275 8517 10287 8551
rect 10229 8511 10287 8517
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 8168 8452 9873 8480
rect 8168 8440 8174 8452
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 11609 8483 11667 8489
rect 11609 8480 11621 8483
rect 10100 8452 11621 8480
rect 10100 8440 10106 8452
rect 11609 8449 11621 8452
rect 11655 8449 11667 8483
rect 11609 8443 11667 8449
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8480 13875 8483
rect 14274 8480 14280 8492
rect 13863 8452 14280 8480
rect 13863 8449 13875 8452
rect 13817 8443 13875 8449
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 5215 8415 5273 8421
rect 5215 8412 5227 8415
rect 5092 8384 5227 8412
rect 4985 8375 5043 8381
rect 5215 8381 5227 8384
rect 5261 8381 5273 8415
rect 7374 8412 7380 8424
rect 7335 8384 7380 8412
rect 5215 8375 5273 8381
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 7558 8412 7564 8424
rect 7519 8384 7564 8412
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 8849 8415 8907 8421
rect 8849 8412 8861 8415
rect 8720 8384 8861 8412
rect 8720 8372 8726 8384
rect 8849 8381 8861 8384
rect 8895 8381 8907 8415
rect 9306 8412 9312 8424
rect 9267 8384 9312 8412
rect 8849 8375 8907 8381
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 10413 8415 10471 8421
rect 10413 8412 10425 8415
rect 9732 8384 10425 8412
rect 9732 8372 9738 8384
rect 10413 8381 10425 8384
rect 10459 8412 10471 8415
rect 10870 8412 10876 8424
rect 10459 8384 10876 8412
rect 10459 8381 10471 8384
rect 10413 8375 10471 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11330 8412 11336 8424
rect 11291 8384 11336 8412
rect 11330 8372 11336 8384
rect 11388 8412 11394 8424
rect 12158 8412 12164 8424
rect 11388 8384 12164 8412
rect 11388 8372 11394 8384
rect 12158 8372 12164 8384
rect 12216 8372 12222 8424
rect 12434 8372 12440 8424
rect 12492 8412 12498 8424
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12492 8384 12909 8412
rect 12492 8372 12498 8384
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 7834 8344 7840 8356
rect 7795 8316 7840 8344
rect 7834 8304 7840 8316
rect 7892 8304 7898 8356
rect 9398 8344 9404 8356
rect 8312 8316 9404 8344
rect 8110 8276 8116 8288
rect 8071 8248 8116 8276
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 8202 8236 8208 8288
rect 8260 8276 8266 8288
rect 8312 8276 8340 8316
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 9582 8344 9588 8356
rect 9543 8316 9588 8344
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 10134 8304 10140 8356
rect 10192 8344 10198 8356
rect 10734 8347 10792 8353
rect 10734 8344 10746 8347
rect 10192 8316 10746 8344
rect 10192 8304 10198 8316
rect 10734 8313 10746 8316
rect 10780 8313 10792 8347
rect 10734 8307 10792 8313
rect 14179 8347 14237 8353
rect 14179 8313 14191 8347
rect 14225 8344 14237 8347
rect 14384 8344 14412 8588
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 17126 8616 17132 8628
rect 17087 8588 17132 8616
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 18506 8576 18512 8628
rect 18564 8616 18570 8628
rect 18601 8619 18659 8625
rect 18601 8616 18613 8619
rect 18564 8588 18613 8616
rect 18564 8576 18570 8588
rect 18601 8585 18613 8588
rect 18647 8585 18659 8619
rect 18601 8579 18659 8585
rect 19058 8576 19064 8628
rect 19116 8616 19122 8628
rect 19245 8619 19303 8625
rect 19245 8616 19257 8619
rect 19116 8588 19257 8616
rect 19116 8576 19122 8588
rect 19245 8585 19257 8588
rect 19291 8585 19303 8619
rect 19245 8579 19303 8585
rect 19705 8619 19763 8625
rect 19705 8585 19717 8619
rect 19751 8616 19763 8619
rect 19978 8616 19984 8628
rect 19751 8588 19984 8616
rect 19751 8585 19763 8588
rect 19705 8579 19763 8585
rect 16666 8548 16672 8560
rect 16627 8520 16672 8548
rect 16666 8508 16672 8520
rect 16724 8508 16730 8560
rect 19260 8548 19288 8579
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 21542 8576 21548 8628
rect 21600 8616 21606 8628
rect 21637 8619 21695 8625
rect 21637 8616 21649 8619
rect 21600 8588 21649 8616
rect 21600 8576 21606 8588
rect 21637 8585 21649 8588
rect 21683 8585 21695 8619
rect 21637 8579 21695 8585
rect 23566 8576 23572 8628
rect 23624 8616 23630 8628
rect 23845 8619 23903 8625
rect 23845 8616 23857 8619
rect 23624 8588 23857 8616
rect 23624 8576 23630 8588
rect 23845 8585 23857 8588
rect 23891 8585 23903 8619
rect 23845 8579 23903 8585
rect 20901 8551 20959 8557
rect 20901 8548 20913 8551
rect 19260 8520 20913 8548
rect 20901 8517 20913 8520
rect 20947 8548 20959 8551
rect 21082 8548 21088 8560
rect 20947 8520 21088 8548
rect 20947 8517 20959 8520
rect 20901 8511 20959 8517
rect 21082 8508 21088 8520
rect 21140 8508 21146 8560
rect 15933 8483 15991 8489
rect 15933 8449 15945 8483
rect 15979 8480 15991 8483
rect 16206 8480 16212 8492
rect 15979 8452 16212 8480
rect 15979 8449 15991 8452
rect 15933 8443 15991 8449
rect 16206 8440 16212 8452
rect 16264 8440 16270 8492
rect 18782 8480 18788 8492
rect 18743 8452 18788 8480
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8480 19947 8483
rect 19978 8480 19984 8492
rect 19935 8452 19984 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 20533 8483 20591 8489
rect 20533 8449 20545 8483
rect 20579 8480 20591 8483
rect 21266 8480 21272 8492
rect 20579 8452 21272 8480
rect 20579 8449 20591 8452
rect 20533 8443 20591 8449
rect 21266 8440 21272 8452
rect 21324 8440 21330 8492
rect 14737 8415 14795 8421
rect 14737 8381 14749 8415
rect 14783 8412 14795 8415
rect 15194 8412 15200 8424
rect 14783 8384 15200 8412
rect 14783 8381 14795 8384
rect 14737 8375 14795 8381
rect 15194 8372 15200 8384
rect 15252 8372 15258 8424
rect 20806 8372 20812 8424
rect 20864 8412 20870 8424
rect 21453 8415 21511 8421
rect 21453 8412 21465 8415
rect 20864 8384 21465 8412
rect 20864 8372 20870 8384
rect 21453 8381 21465 8384
rect 21499 8412 21511 8415
rect 21634 8412 21640 8424
rect 21499 8384 21640 8412
rect 21499 8381 21511 8384
rect 21453 8375 21511 8381
rect 21634 8372 21640 8384
rect 21692 8372 21698 8424
rect 23474 8372 23480 8424
rect 23532 8412 23538 8424
rect 24397 8415 24455 8421
rect 24397 8412 24409 8415
rect 23532 8384 24409 8412
rect 23532 8372 23538 8384
rect 24397 8381 24409 8384
rect 24443 8412 24455 8415
rect 24949 8415 25007 8421
rect 24949 8412 24961 8415
rect 24443 8384 24961 8412
rect 24443 8381 24455 8384
rect 24397 8375 24455 8381
rect 24949 8381 24961 8384
rect 24995 8381 25007 8415
rect 24949 8375 25007 8381
rect 16114 8344 16120 8356
rect 14225 8316 14412 8344
rect 16075 8316 16120 8344
rect 14225 8313 14237 8316
rect 14179 8307 14237 8313
rect 16114 8304 16120 8316
rect 16172 8304 16178 8356
rect 16206 8304 16212 8356
rect 16264 8344 16270 8356
rect 19981 8347 20039 8353
rect 16264 8316 16309 8344
rect 16264 8304 16270 8316
rect 19981 8313 19993 8347
rect 20027 8344 20039 8347
rect 20070 8344 20076 8356
rect 20027 8316 20076 8344
rect 20027 8313 20039 8316
rect 19981 8307 20039 8313
rect 20070 8304 20076 8316
rect 20128 8304 20134 8356
rect 8260 8248 8340 8276
rect 8260 8236 8266 8248
rect 10962 8236 10968 8288
rect 11020 8276 11026 8288
rect 12621 8279 12679 8285
rect 12621 8276 12633 8279
rect 11020 8248 12633 8276
rect 11020 8236 11026 8248
rect 12621 8245 12633 8248
rect 12667 8245 12679 8279
rect 12621 8239 12679 8245
rect 24581 8279 24639 8285
rect 24581 8245 24593 8279
rect 24627 8276 24639 8279
rect 24670 8276 24676 8288
rect 24627 8248 24676 8276
rect 24627 8245 24639 8248
rect 24581 8239 24639 8245
rect 24670 8236 24676 8248
rect 24728 8236 24734 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 5997 8075 6055 8081
rect 5997 8041 6009 8075
rect 6043 8072 6055 8075
rect 7558 8072 7564 8084
rect 6043 8044 7564 8072
rect 6043 8041 6055 8044
rect 5997 8035 6055 8041
rect 5166 7936 5172 7948
rect 5127 7908 5172 7936
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 5353 7939 5411 7945
rect 5353 7905 5365 7939
rect 5399 7936 5411 7939
rect 5534 7936 5540 7948
rect 5399 7908 5540 7936
rect 5399 7905 5411 7908
rect 5353 7899 5411 7905
rect 5534 7896 5540 7908
rect 5592 7936 5598 7948
rect 6012 7936 6040 8035
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 7834 8072 7840 8084
rect 7795 8044 7840 8072
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 10042 8072 10048 8084
rect 10003 8044 10048 8072
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 10870 8072 10876 8084
rect 10831 8044 10876 8072
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 12894 8072 12900 8084
rect 12855 8044 12900 8072
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14645 8075 14703 8081
rect 14645 8072 14657 8075
rect 14332 8044 14657 8072
rect 14332 8032 14338 8044
rect 14645 8041 14657 8044
rect 14691 8041 14703 8075
rect 14645 8035 14703 8041
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 19518 8081 19524 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14884 8044 15025 8072
rect 14884 8032 14890 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 19475 8075 19524 8081
rect 19475 8041 19487 8075
rect 19521 8041 19524 8075
rect 19475 8035 19524 8041
rect 19518 8032 19524 8035
rect 19576 8032 19582 8084
rect 20990 8032 20996 8084
rect 21048 8072 21054 8084
rect 21361 8075 21419 8081
rect 21361 8072 21373 8075
rect 21048 8044 21373 8072
rect 21048 8032 21054 8044
rect 21361 8041 21373 8044
rect 21407 8041 21419 8075
rect 21361 8035 21419 8041
rect 21634 8032 21640 8084
rect 21692 8072 21698 8084
rect 21729 8075 21787 8081
rect 21729 8072 21741 8075
rect 21692 8044 21741 8072
rect 21692 8032 21698 8044
rect 21729 8041 21741 8044
rect 21775 8041 21787 8075
rect 24762 8072 24768 8084
rect 24723 8044 24768 8072
rect 21729 8035 21787 8041
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 11241 8007 11299 8013
rect 7024 7976 8616 8004
rect 6454 7936 6460 7948
rect 5592 7908 6040 7936
rect 6415 7908 6460 7936
rect 5592 7896 5598 7908
rect 6454 7896 6460 7908
rect 6512 7896 6518 7948
rect 6546 7896 6552 7948
rect 6604 7936 6610 7948
rect 7024 7945 7052 7976
rect 7009 7939 7067 7945
rect 7009 7936 7021 7939
rect 6604 7908 7021 7936
rect 6604 7896 6610 7908
rect 7009 7905 7021 7908
rect 7055 7905 7067 7939
rect 7009 7899 7067 7905
rect 7926 7896 7932 7948
rect 7984 7936 7990 7948
rect 8202 7936 8208 7948
rect 7984 7908 8208 7936
rect 7984 7896 7990 7908
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8588 7945 8616 7976
rect 9324 7976 10272 8004
rect 9324 7948 9352 7976
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7936 8631 7939
rect 8662 7936 8668 7948
rect 8619 7908 8668 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 8662 7896 8668 7908
rect 8720 7936 8726 7948
rect 9306 7936 9312 7948
rect 8720 7908 9312 7936
rect 8720 7896 8726 7908
rect 9306 7896 9312 7908
rect 9364 7896 9370 7948
rect 9766 7936 9772 7948
rect 9727 7908 9772 7936
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 10244 7945 10272 7976
rect 11241 7973 11253 8007
rect 11287 8004 11299 8007
rect 11422 8004 11428 8016
rect 11287 7976 11428 8004
rect 11287 7973 11299 7976
rect 11241 7967 11299 7973
rect 11422 7964 11428 7976
rect 11480 7964 11486 8016
rect 11517 8007 11575 8013
rect 11517 7973 11529 8007
rect 11563 8004 11575 8007
rect 11698 8004 11704 8016
rect 11563 7976 11704 8004
rect 11563 7973 11575 7976
rect 11517 7967 11575 7973
rect 11698 7964 11704 7976
rect 11756 7964 11762 8016
rect 13814 8004 13820 8016
rect 13775 7976 13820 8004
rect 13814 7964 13820 7976
rect 13872 7964 13878 8016
rect 15194 7964 15200 8016
rect 15252 8004 15258 8016
rect 15470 8004 15476 8016
rect 15252 7976 15476 8004
rect 15252 7964 15258 7976
rect 15470 7964 15476 7976
rect 15528 7964 15534 8016
rect 16022 8004 16028 8016
rect 15983 7976 16028 8004
rect 16022 7964 16028 7976
rect 16080 7964 16086 8016
rect 17862 7964 17868 8016
rect 17920 8013 17926 8016
rect 17920 8007 17968 8013
rect 17920 7973 17922 8007
rect 17956 7973 17968 8007
rect 17920 7967 17968 7973
rect 17920 7964 17926 7967
rect 10229 7939 10287 7945
rect 10229 7905 10241 7939
rect 10275 7936 10287 7939
rect 10870 7936 10876 7948
rect 10275 7908 10876 7936
rect 10275 7905 10287 7908
rect 10229 7899 10287 7905
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 17589 7939 17647 7945
rect 17589 7905 17601 7939
rect 17635 7936 17647 7939
rect 17678 7936 17684 7948
rect 17635 7908 17684 7936
rect 17635 7905 17647 7908
rect 17589 7899 17647 7905
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 19404 7939 19462 7945
rect 19404 7905 19416 7939
rect 19450 7936 19462 7939
rect 20968 7939 21026 7945
rect 19450 7908 20024 7936
rect 19450 7905 19462 7908
rect 19404 7899 19462 7905
rect 19996 7880 20024 7908
rect 20968 7905 20980 7939
rect 21014 7936 21026 7939
rect 21174 7936 21180 7948
rect 21014 7908 21180 7936
rect 21014 7905 21026 7908
rect 20968 7899 21026 7905
rect 21174 7896 21180 7908
rect 21232 7936 21238 7948
rect 21726 7936 21732 7948
rect 21232 7908 21732 7936
rect 21232 7896 21238 7908
rect 21726 7896 21732 7908
rect 21784 7896 21790 7948
rect 24578 7936 24584 7948
rect 24539 7908 24584 7936
rect 24578 7896 24584 7908
rect 24636 7936 24642 7948
rect 25406 7936 25412 7948
rect 24636 7908 25412 7936
rect 24636 7896 24642 7908
rect 25406 7896 25412 7908
rect 25464 7896 25470 7948
rect 5442 7868 5448 7880
rect 5403 7840 5448 7868
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 7190 7868 7196 7880
rect 7151 7840 7196 7868
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 8754 7868 8760 7880
rect 8715 7840 8760 7868
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 11514 7828 11520 7880
rect 11572 7868 11578 7880
rect 11701 7871 11759 7877
rect 11701 7868 11713 7871
rect 11572 7840 11713 7868
rect 11572 7828 11578 7840
rect 11701 7837 11713 7840
rect 11747 7837 11759 7871
rect 13722 7868 13728 7880
rect 13683 7840 13728 7868
rect 11701 7831 11759 7837
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 15378 7868 15384 7880
rect 15339 7840 15384 7868
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 19978 7828 19984 7880
rect 20036 7828 20042 7880
rect 12434 7760 12440 7812
rect 12492 7800 12498 7812
rect 14277 7803 14335 7809
rect 12492 7772 12537 7800
rect 12492 7760 12498 7772
rect 14277 7769 14289 7803
rect 14323 7800 14335 7803
rect 16114 7800 16120 7812
rect 14323 7772 16120 7800
rect 14323 7769 14335 7772
rect 14277 7763 14335 7769
rect 16114 7760 16120 7772
rect 16172 7800 16178 7812
rect 16301 7803 16359 7809
rect 16301 7800 16313 7803
rect 16172 7772 16313 7800
rect 16172 7760 16178 7772
rect 16301 7769 16313 7772
rect 16347 7769 16359 7803
rect 16301 7763 16359 7769
rect 18509 7803 18567 7809
rect 18509 7769 18521 7803
rect 18555 7800 18567 7803
rect 18966 7800 18972 7812
rect 18555 7772 18972 7800
rect 18555 7769 18567 7772
rect 18509 7763 18567 7769
rect 18966 7760 18972 7772
rect 19024 7760 19030 7812
rect 9214 7732 9220 7744
rect 9175 7704 9220 7732
rect 9214 7692 9220 7704
rect 9272 7692 9278 7744
rect 18874 7732 18880 7744
rect 18835 7704 18880 7732
rect 18874 7692 18880 7704
rect 18932 7692 18938 7744
rect 19886 7732 19892 7744
rect 19847 7704 19892 7732
rect 19886 7692 19892 7704
rect 19944 7692 19950 7744
rect 21039 7735 21097 7741
rect 21039 7701 21051 7735
rect 21085 7732 21097 7735
rect 21266 7732 21272 7744
rect 21085 7704 21272 7732
rect 21085 7701 21097 7704
rect 21039 7695 21097 7701
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 4709 7531 4767 7537
rect 4709 7497 4721 7531
rect 4755 7528 4767 7531
rect 5166 7528 5172 7540
rect 4755 7500 5172 7528
rect 4755 7497 4767 7500
rect 4709 7491 4767 7497
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 6546 7528 6552 7540
rect 6507 7500 6552 7528
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 8662 7528 8668 7540
rect 8623 7500 8668 7528
rect 8662 7488 8668 7500
rect 8720 7528 8726 7540
rect 8941 7531 8999 7537
rect 8941 7528 8953 7531
rect 8720 7500 8953 7528
rect 8720 7488 8726 7500
rect 8941 7497 8953 7500
rect 8987 7497 8999 7531
rect 8941 7491 8999 7497
rect 9766 7488 9772 7540
rect 9824 7528 9830 7540
rect 10137 7531 10195 7537
rect 10137 7528 10149 7531
rect 9824 7500 10149 7528
rect 9824 7488 9830 7500
rect 10137 7497 10149 7500
rect 10183 7497 10195 7531
rect 11698 7528 11704 7540
rect 11659 7500 11704 7528
rect 10137 7491 10195 7497
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 13078 7528 13084 7540
rect 12176 7500 13084 7528
rect 10502 7460 10508 7472
rect 10463 7432 10508 7460
rect 10502 7420 10508 7432
rect 10560 7420 10566 7472
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7392 5043 7395
rect 5031 7364 5488 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 5460 7336 5488 7364
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 9214 7392 9220 7404
rect 8352 7364 9220 7392
rect 8352 7352 8358 7364
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 9674 7392 9680 7404
rect 9635 7364 9680 7392
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 3694 7324 3700 7336
rect 3655 7296 3700 7324
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 4157 7327 4215 7333
rect 4157 7293 4169 7327
rect 4203 7324 4215 7327
rect 5074 7324 5080 7336
rect 4203 7296 5080 7324
rect 4203 7293 4215 7296
rect 4157 7287 4215 7293
rect 2774 7216 2780 7268
rect 2832 7256 2838 7268
rect 3513 7259 3571 7265
rect 3513 7256 3525 7259
rect 2832 7228 3525 7256
rect 2832 7216 2838 7228
rect 3513 7225 3525 7228
rect 3559 7256 3571 7259
rect 4172 7256 4200 7287
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 5442 7324 5448 7336
rect 5403 7296 5448 7324
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5592 7296 5641 7324
rect 5592 7284 5598 7296
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 7064 7296 7389 7324
rect 7064 7284 7070 7296
rect 7377 7293 7389 7296
rect 7423 7293 7435 7327
rect 10520 7324 10548 7420
rect 11238 7392 11244 7404
rect 11199 7364 11244 7392
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 10689 7327 10747 7333
rect 10689 7324 10701 7327
rect 10520 7296 10701 7324
rect 7377 7287 7435 7293
rect 10689 7293 10701 7296
rect 10735 7293 10747 7327
rect 10689 7287 10747 7293
rect 10870 7284 10876 7336
rect 10928 7324 10934 7336
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 10928 7296 11161 7324
rect 10928 7284 10934 7296
rect 11149 7293 11161 7296
rect 11195 7293 11207 7327
rect 11149 7287 11207 7293
rect 3559 7228 4200 7256
rect 5905 7259 5963 7265
rect 3559 7225 3571 7228
rect 3513 7219 3571 7225
rect 5905 7225 5917 7259
rect 5951 7256 5963 7259
rect 6178 7256 6184 7268
rect 5951 7228 6184 7256
rect 5951 7225 5963 7228
rect 5905 7219 5963 7225
rect 6178 7216 6184 7228
rect 6236 7216 6242 7268
rect 7698 7259 7756 7265
rect 7698 7256 7710 7259
rect 7208 7228 7710 7256
rect 3878 7188 3884 7200
rect 3839 7160 3884 7188
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 7098 7148 7104 7200
rect 7156 7188 7162 7200
rect 7208 7197 7236 7228
rect 7698 7225 7710 7228
rect 7744 7256 7756 7259
rect 8110 7256 8116 7268
rect 7744 7228 8116 7256
rect 7744 7225 7756 7228
rect 7698 7219 7756 7225
rect 8110 7216 8116 7228
rect 8168 7216 8174 7268
rect 9309 7259 9367 7265
rect 8312 7228 9168 7256
rect 8312 7197 8340 7228
rect 9140 7200 9168 7228
rect 9309 7225 9321 7259
rect 9355 7225 9367 7259
rect 9309 7219 9367 7225
rect 7193 7191 7251 7197
rect 7193 7188 7205 7191
rect 7156 7160 7205 7188
rect 7156 7148 7162 7160
rect 7193 7157 7205 7160
rect 7239 7157 7251 7191
rect 7193 7151 7251 7157
rect 8297 7191 8355 7197
rect 8297 7157 8309 7191
rect 8343 7157 8355 7191
rect 8297 7151 8355 7157
rect 9122 7148 9128 7200
rect 9180 7188 9186 7200
rect 9324 7188 9352 7219
rect 9180 7160 9352 7188
rect 9180 7148 9186 7160
rect 11606 7148 11612 7200
rect 11664 7188 11670 7200
rect 12176 7197 12204 7500
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 14507 7531 14565 7537
rect 14507 7497 14519 7531
rect 14553 7528 14565 7531
rect 15378 7528 15384 7540
rect 14553 7500 15384 7528
rect 14553 7497 14565 7500
rect 14507 7491 14565 7497
rect 15378 7488 15384 7500
rect 15436 7528 15442 7540
rect 16761 7531 16819 7537
rect 16761 7528 16773 7531
rect 15436 7500 16773 7528
rect 15436 7488 15442 7500
rect 16761 7497 16773 7500
rect 16807 7497 16819 7531
rect 16761 7491 16819 7497
rect 17678 7488 17684 7540
rect 17736 7528 17742 7540
rect 20530 7537 20536 7540
rect 18233 7531 18291 7537
rect 18233 7528 18245 7531
rect 17736 7500 18245 7528
rect 17736 7488 17742 7500
rect 18233 7497 18245 7500
rect 18279 7497 18291 7531
rect 18233 7491 18291 7497
rect 20487 7531 20536 7537
rect 20487 7497 20499 7531
rect 20533 7497 20536 7531
rect 20487 7491 20536 7497
rect 20530 7488 20536 7491
rect 20588 7488 20594 7540
rect 21174 7528 21180 7540
rect 21135 7500 21180 7528
rect 21174 7488 21180 7500
rect 21232 7488 21238 7540
rect 23474 7488 23480 7540
rect 23532 7528 23538 7540
rect 24719 7531 24777 7537
rect 24719 7528 24731 7531
rect 23532 7500 24731 7528
rect 23532 7488 23538 7500
rect 24719 7497 24731 7500
rect 24765 7497 24777 7531
rect 25406 7528 25412 7540
rect 25367 7500 25412 7528
rect 24719 7491 24777 7497
rect 25406 7488 25412 7500
rect 25464 7488 25470 7540
rect 13722 7420 13728 7472
rect 13780 7460 13786 7472
rect 14093 7463 14151 7469
rect 14093 7460 14105 7463
rect 13780 7432 14105 7460
rect 13780 7420 13786 7432
rect 14093 7429 14105 7432
rect 14139 7460 14151 7463
rect 14139 7432 16988 7460
rect 14139 7429 14151 7432
rect 14093 7423 14151 7429
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 14918 7392 14924 7404
rect 12492 7364 12537 7392
rect 14879 7364 14924 7392
rect 12492 7352 12498 7364
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15194 7352 15200 7404
rect 15252 7392 15258 7404
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15252 7364 15485 7392
rect 15252 7352 15258 7364
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15930 7392 15936 7404
rect 15891 7364 15936 7392
rect 15473 7355 15531 7361
rect 15930 7352 15936 7364
rect 15988 7352 15994 7404
rect 16960 7401 16988 7432
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 17862 7392 17868 7404
rect 17727 7364 17868 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 18874 7392 18880 7404
rect 18835 7364 18880 7392
rect 18874 7352 18880 7364
rect 18932 7352 18938 7404
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7324 13415 7327
rect 13722 7324 13728 7336
rect 13403 7296 13728 7324
rect 13403 7293 13415 7296
rect 13357 7287 13415 7293
rect 13722 7284 13728 7296
rect 13780 7284 13786 7336
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 14436 7327 14494 7333
rect 14436 7324 14448 7327
rect 13964 7296 14448 7324
rect 13964 7284 13970 7296
rect 14436 7293 14448 7296
rect 14482 7324 14494 7327
rect 14936 7324 14964 7352
rect 24670 7333 24676 7336
rect 20384 7327 20442 7333
rect 20384 7324 20396 7327
rect 14482 7296 14964 7324
rect 19536 7296 20396 7324
rect 14482 7293 14494 7296
rect 14436 7287 14494 7293
rect 19536 7268 19564 7296
rect 20384 7293 20396 7296
rect 20430 7324 20442 7327
rect 20809 7327 20867 7333
rect 20809 7324 20821 7327
rect 20430 7296 20821 7324
rect 20430 7293 20442 7296
rect 20384 7287 20442 7293
rect 20809 7293 20821 7296
rect 20855 7293 20867 7327
rect 24648 7327 24676 7333
rect 24648 7324 24660 7327
rect 24583 7296 24660 7324
rect 20809 7287 20867 7293
rect 24648 7293 24660 7296
rect 24728 7324 24734 7336
rect 25041 7327 25099 7333
rect 25041 7324 25053 7327
rect 24728 7296 25053 7324
rect 24648 7287 24676 7293
rect 24670 7284 24676 7287
rect 24728 7284 24734 7296
rect 25041 7293 25053 7296
rect 25087 7293 25099 7327
rect 25041 7287 25099 7293
rect 12799 7259 12857 7265
rect 12799 7225 12811 7259
rect 12845 7256 12857 7259
rect 13078 7256 13084 7268
rect 12845 7228 13084 7256
rect 12845 7225 12857 7228
rect 12799 7219 12857 7225
rect 13078 7216 13084 7228
rect 13136 7216 13142 7268
rect 13633 7259 13691 7265
rect 13633 7225 13645 7259
rect 13679 7256 13691 7259
rect 13814 7256 13820 7268
rect 13679 7228 13820 7256
rect 13679 7225 13691 7228
rect 13633 7219 13691 7225
rect 13814 7216 13820 7228
rect 13872 7256 13878 7268
rect 15565 7259 15623 7265
rect 15565 7256 15577 7259
rect 13872 7228 15577 7256
rect 13872 7216 13878 7228
rect 15304 7200 15332 7228
rect 15565 7225 15577 7228
rect 15611 7225 15623 7259
rect 15565 7219 15623 7225
rect 18693 7259 18751 7265
rect 18693 7225 18705 7259
rect 18739 7256 18751 7259
rect 18966 7256 18972 7268
rect 18739 7228 18972 7256
rect 18739 7225 18751 7228
rect 18693 7219 18751 7225
rect 18966 7216 18972 7228
rect 19024 7216 19030 7268
rect 19518 7256 19524 7268
rect 19479 7228 19524 7256
rect 19518 7216 19524 7228
rect 19576 7216 19582 7268
rect 12161 7191 12219 7197
rect 12161 7188 12173 7191
rect 11664 7160 12173 7188
rect 11664 7148 11670 7160
rect 12161 7157 12173 7160
rect 12207 7157 12219 7191
rect 15286 7188 15292 7200
rect 15247 7160 15292 7188
rect 12161 7151 12219 7157
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15470 7148 15476 7200
rect 15528 7188 15534 7200
rect 16393 7191 16451 7197
rect 16393 7188 16405 7191
rect 15528 7160 16405 7188
rect 15528 7148 15534 7160
rect 16393 7157 16405 7160
rect 16439 7157 16451 7191
rect 16393 7151 16451 7157
rect 19889 7191 19947 7197
rect 19889 7157 19901 7191
rect 19935 7188 19947 7191
rect 19978 7188 19984 7200
rect 19935 7160 19984 7188
rect 19935 7157 19947 7160
rect 19889 7151 19947 7157
rect 19978 7148 19984 7160
rect 20036 7148 20042 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 3694 6984 3700 6996
rect 3655 6956 3700 6984
rect 3694 6944 3700 6956
rect 3752 6984 3758 6996
rect 6454 6984 6460 6996
rect 3752 6956 6460 6984
rect 3752 6944 3758 6956
rect 6454 6944 6460 6956
rect 6512 6944 6518 6996
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7064 6956 7420 6984
rect 7064 6944 7070 6956
rect 4985 6919 5043 6925
rect 4985 6885 4997 6919
rect 5031 6916 5043 6919
rect 5074 6916 5080 6928
rect 5031 6888 5080 6916
rect 5031 6885 5043 6888
rect 4985 6879 5043 6885
rect 5074 6876 5080 6888
rect 5132 6916 5138 6928
rect 5132 6888 5580 6916
rect 5132 6876 5138 6888
rect 5552 6860 5580 6888
rect 7098 6876 7104 6928
rect 7156 6916 7162 6928
rect 7238 6919 7296 6925
rect 7238 6916 7250 6919
rect 7156 6888 7250 6916
rect 7156 6876 7162 6888
rect 7238 6885 7250 6888
rect 7284 6885 7296 6919
rect 7392 6916 7420 6956
rect 7926 6944 7932 6996
rect 7984 6984 7990 6996
rect 8113 6987 8171 6993
rect 8113 6984 8125 6987
rect 7984 6956 8125 6984
rect 7984 6944 7990 6956
rect 8113 6953 8125 6956
rect 8159 6953 8171 6987
rect 9122 6984 9128 6996
rect 9083 6956 9128 6984
rect 8113 6947 8171 6953
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 10781 6987 10839 6993
rect 10781 6953 10793 6987
rect 10827 6984 10839 6987
rect 10870 6984 10876 6996
rect 10827 6956 10876 6984
rect 10827 6953 10839 6956
rect 10781 6947 10839 6953
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 11149 6987 11207 6993
rect 11149 6953 11161 6987
rect 11195 6984 11207 6987
rect 11238 6984 11244 6996
rect 11195 6956 11244 6984
rect 11195 6953 11207 6956
rect 11149 6947 11207 6953
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 9858 6916 9864 6928
rect 7392 6888 8248 6916
rect 9819 6888 9864 6916
rect 7238 6879 7296 6885
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 5460 6780 5488 6811
rect 5534 6808 5540 6860
rect 5592 6848 5598 6860
rect 5813 6851 5871 6857
rect 5813 6848 5825 6851
rect 5592 6820 5825 6848
rect 5592 6808 5598 6820
rect 5813 6817 5825 6820
rect 5859 6817 5871 6851
rect 5994 6848 6000 6860
rect 5813 6811 5871 6817
rect 5920 6820 6000 6848
rect 5920 6780 5948 6820
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 6914 6848 6920 6860
rect 6875 6820 6920 6848
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 8220 6848 8248 6888
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 11606 6925 11612 6928
rect 11603 6916 11612 6925
rect 11567 6888 11612 6916
rect 11603 6879 11612 6888
rect 11606 6876 11612 6879
rect 11664 6876 11670 6928
rect 13170 6916 13176 6928
rect 13131 6888 13176 6916
rect 13170 6876 13176 6888
rect 13228 6876 13234 6928
rect 15470 6916 15476 6928
rect 15431 6888 15476 6916
rect 15470 6876 15476 6888
rect 15528 6876 15534 6928
rect 16025 6919 16083 6925
rect 16025 6885 16037 6919
rect 16071 6916 16083 6919
rect 16114 6916 16120 6928
rect 16071 6888 16120 6916
rect 16071 6885 16083 6888
rect 16025 6879 16083 6885
rect 16114 6876 16120 6888
rect 16172 6876 16178 6928
rect 17215 6919 17273 6925
rect 17215 6885 17227 6919
rect 17261 6916 17273 6919
rect 17402 6916 17408 6928
rect 17261 6888 17408 6916
rect 17261 6885 17273 6888
rect 17215 6879 17273 6885
rect 17402 6876 17408 6888
rect 17460 6916 17466 6928
rect 17862 6916 17868 6928
rect 17460 6888 17868 6916
rect 17460 6876 17466 6888
rect 17862 6876 17868 6888
rect 17920 6876 17926 6928
rect 18782 6916 18788 6928
rect 18743 6888 18788 6916
rect 18782 6876 18788 6888
rect 18840 6876 18846 6928
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 8220 6820 8493 6848
rect 8481 6817 8493 6820
rect 8527 6817 8539 6851
rect 8481 6811 8539 6817
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 11241 6851 11299 6857
rect 11241 6848 11253 6851
rect 11204 6820 11253 6848
rect 11204 6808 11210 6820
rect 11241 6817 11253 6820
rect 11287 6817 11299 6851
rect 12526 6848 12532 6860
rect 12487 6820 12532 6848
rect 11241 6811 11299 6817
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 16850 6848 16856 6860
rect 16811 6820 16856 6848
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 20990 6848 20996 6860
rect 20951 6820 20996 6848
rect 20990 6808 20996 6820
rect 21048 6808 21054 6860
rect 6086 6780 6092 6792
rect 5460 6752 5948 6780
rect 6047 6752 6092 6780
rect 6086 6740 6092 6752
rect 6144 6740 6150 6792
rect 9030 6740 9036 6792
rect 9088 6780 9094 6792
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 9088 6752 9781 6780
rect 9088 6740 9094 6752
rect 9769 6749 9781 6752
rect 9815 6749 9827 6783
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 9769 6743 9827 6749
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6780 13139 6783
rect 13262 6780 13268 6792
rect 13127 6752 13268 6780
rect 13127 6749 13139 6752
rect 13081 6743 13139 6749
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6749 13415 6783
rect 15378 6780 15384 6792
rect 15339 6752 15384 6780
rect 13357 6743 13415 6749
rect 12986 6672 12992 6724
rect 13044 6712 13050 6724
rect 13372 6712 13400 6743
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 18690 6780 18696 6792
rect 18651 6752 18696 6780
rect 18690 6740 18696 6752
rect 18748 6740 18754 6792
rect 18874 6740 18880 6792
rect 18932 6780 18938 6792
rect 18969 6783 19027 6789
rect 18969 6780 18981 6783
rect 18932 6752 18981 6780
rect 18932 6740 18938 6752
rect 18969 6749 18981 6752
rect 19015 6749 19027 6783
rect 20898 6780 20904 6792
rect 20859 6752 20904 6780
rect 18969 6743 19027 6749
rect 20898 6740 20904 6752
rect 20956 6740 20962 6792
rect 13998 6712 14004 6724
rect 13044 6684 14004 6712
rect 13044 6672 13050 6684
rect 13998 6672 14004 6684
rect 14056 6672 14062 6724
rect 15102 6672 15108 6724
rect 15160 6672 15166 6724
rect 7834 6644 7840 6656
rect 7795 6616 7840 6644
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 12158 6644 12164 6656
rect 12119 6616 12164 6644
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 14274 6644 14280 6656
rect 14235 6616 14280 6644
rect 14274 6604 14280 6616
rect 14332 6604 14338 6656
rect 14826 6604 14832 6656
rect 14884 6644 14890 6656
rect 15013 6647 15071 6653
rect 15013 6644 15025 6647
rect 14884 6616 15025 6644
rect 14884 6604 14890 6616
rect 15013 6613 15025 6616
rect 15059 6644 15071 6647
rect 15120 6644 15148 6672
rect 17770 6644 17776 6656
rect 15059 6616 15148 6644
rect 17731 6616 17776 6644
rect 15059 6613 15071 6616
rect 15013 6607 15071 6613
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 18049 6647 18107 6653
rect 18049 6644 18061 6647
rect 18012 6616 18061 6644
rect 18012 6604 18018 6616
rect 18049 6613 18061 6616
rect 18095 6613 18107 6647
rect 18049 6607 18107 6613
rect 19426 6604 19432 6656
rect 19484 6644 19490 6656
rect 19613 6647 19671 6653
rect 19613 6644 19625 6647
rect 19484 6616 19625 6644
rect 19484 6604 19490 6616
rect 19613 6613 19625 6616
rect 19659 6613 19671 6647
rect 19613 6607 19671 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 5074 6440 5080 6452
rect 5035 6412 5080 6440
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 5994 6400 6000 6452
rect 6052 6440 6058 6452
rect 6181 6443 6239 6449
rect 6181 6440 6193 6443
rect 6052 6412 6193 6440
rect 6052 6400 6058 6412
rect 6181 6409 6193 6412
rect 6227 6409 6239 6443
rect 6181 6403 6239 6409
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 6914 6440 6920 6452
rect 6687 6412 6920 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 9030 6440 9036 6452
rect 8991 6412 9036 6440
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 9398 6440 9404 6452
rect 9311 6412 9404 6440
rect 9398 6400 9404 6412
rect 9456 6440 9462 6452
rect 9858 6440 9864 6452
rect 9456 6412 9864 6440
rect 9456 6400 9462 6412
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 10284 6412 10425 6440
rect 10284 6400 10290 6412
rect 10413 6409 10425 6412
rect 10459 6409 10471 6443
rect 10413 6403 10471 6409
rect 11517 6443 11575 6449
rect 11517 6409 11529 6443
rect 11563 6440 11575 6443
rect 11790 6440 11796 6452
rect 11563 6412 11796 6440
rect 11563 6409 11575 6412
rect 11517 6403 11575 6409
rect 6086 6264 6092 6316
rect 6144 6304 6150 6316
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 6144 6276 7757 6304
rect 6144 6264 6150 6276
rect 7745 6273 7757 6276
rect 7791 6304 7803 6307
rect 8294 6304 8300 6316
rect 7791 6276 8300 6304
rect 7791 6273 7803 6276
rect 7745 6267 7803 6273
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 5442 6236 5448 6248
rect 4755 6208 5448 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 5534 6196 5540 6248
rect 5592 6236 5598 6248
rect 5629 6239 5687 6245
rect 5629 6236 5641 6239
rect 5592 6208 5641 6236
rect 5592 6196 5598 6208
rect 5629 6205 5641 6208
rect 5675 6205 5687 6239
rect 5629 6199 5687 6205
rect 5905 6239 5963 6245
rect 5905 6205 5917 6239
rect 5951 6236 5963 6239
rect 7006 6236 7012 6248
rect 5951 6208 7012 6236
rect 5951 6205 5963 6208
rect 5905 6199 5963 6205
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6236 8723 6239
rect 9122 6236 9128 6248
rect 8711 6208 9128 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 9560 6239 9618 6245
rect 9560 6205 9572 6239
rect 9606 6236 9618 6239
rect 9606 6208 10088 6236
rect 9606 6205 9618 6208
rect 9560 6199 9618 6205
rect 8066 6171 8124 6177
rect 8066 6168 8078 6171
rect 7576 6140 8078 6168
rect 7098 6100 7104 6112
rect 7059 6072 7104 6100
rect 7098 6060 7104 6072
rect 7156 6100 7162 6112
rect 7576 6109 7604 6140
rect 8066 6137 8078 6140
rect 8112 6137 8124 6171
rect 8066 6131 8124 6137
rect 10060 6112 10088 6208
rect 10428 6168 10456 6403
rect 11790 6400 11796 6412
rect 11848 6440 11854 6452
rect 13170 6440 13176 6452
rect 11848 6412 13176 6440
rect 11848 6400 11854 6412
rect 13170 6400 13176 6412
rect 13228 6440 13234 6452
rect 13633 6443 13691 6449
rect 13633 6440 13645 6443
rect 13228 6412 13645 6440
rect 13228 6400 13234 6412
rect 13633 6409 13645 6412
rect 13679 6409 13691 6443
rect 13633 6403 13691 6409
rect 15381 6443 15439 6449
rect 15381 6409 15393 6443
rect 15427 6440 15439 6443
rect 15470 6440 15476 6452
rect 15427 6412 15476 6440
rect 15427 6409 15439 6412
rect 15381 6403 15439 6409
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 17402 6440 17408 6452
rect 17363 6412 17408 6440
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 18782 6400 18788 6452
rect 18840 6400 18846 6452
rect 20990 6440 20996 6452
rect 20951 6412 20996 6440
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 18800 6372 18828 6400
rect 19061 6375 19119 6381
rect 19061 6372 19073 6375
rect 17144 6344 19073 6372
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6304 10655 6307
rect 11238 6304 11244 6316
rect 10643 6276 11244 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12526 6304 12532 6316
rect 12483 6276 12532 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 12526 6264 12532 6276
rect 12584 6264 12590 6316
rect 14274 6304 14280 6316
rect 14235 6276 14280 6304
rect 14274 6264 14280 6276
rect 14332 6264 14338 6316
rect 14366 6264 14372 6316
rect 14424 6304 14430 6316
rect 14553 6307 14611 6313
rect 14553 6304 14565 6307
rect 14424 6276 14565 6304
rect 14424 6264 14430 6276
rect 14553 6273 14565 6276
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 14734 6264 14740 6316
rect 14792 6304 14798 6316
rect 15378 6304 15384 6316
rect 14792 6276 15384 6304
rect 14792 6264 14798 6276
rect 15378 6264 15384 6276
rect 15436 6304 15442 6316
rect 17144 6313 17172 6344
rect 19061 6341 19073 6344
rect 19107 6372 19119 6375
rect 19429 6375 19487 6381
rect 19429 6372 19441 6375
rect 19107 6344 19441 6372
rect 19107 6341 19119 6344
rect 19061 6335 19119 6341
rect 19429 6341 19441 6344
rect 19475 6372 19487 6375
rect 19794 6372 19800 6384
rect 19475 6344 19800 6372
rect 19475 6341 19487 6344
rect 19429 6335 19487 6341
rect 19794 6332 19800 6344
rect 19852 6332 19858 6384
rect 24762 6372 24768 6384
rect 24723 6344 24768 6372
rect 24762 6332 24768 6344
rect 24820 6332 24826 6384
rect 15657 6307 15715 6313
rect 15657 6304 15669 6307
rect 15436 6276 15669 6304
rect 15436 6264 15442 6276
rect 15657 6273 15669 6276
rect 15703 6273 15715 6307
rect 15657 6267 15715 6273
rect 17129 6307 17187 6313
rect 17129 6273 17141 6307
rect 17175 6273 17187 6307
rect 17129 6267 17187 6273
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6304 18843 6307
rect 18874 6304 18880 6316
rect 18831 6276 18880 6304
rect 18831 6273 18843 6276
rect 18785 6267 18843 6273
rect 18874 6264 18880 6276
rect 18932 6264 18938 6316
rect 19334 6264 19340 6316
rect 19392 6304 19398 6316
rect 19981 6307 20039 6313
rect 19981 6304 19993 6307
rect 19392 6276 19993 6304
rect 19392 6264 19398 6276
rect 19981 6273 19993 6276
rect 20027 6273 20039 6307
rect 19981 6267 20039 6273
rect 13357 6239 13415 6245
rect 13357 6205 13369 6239
rect 13403 6236 13415 6239
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13403 6208 14013 6236
rect 13403 6205 13415 6208
rect 13357 6199 13415 6205
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 16301 6239 16359 6245
rect 16301 6205 16313 6239
rect 16347 6236 16359 6239
rect 16485 6239 16543 6245
rect 16485 6236 16497 6239
rect 16347 6208 16497 6236
rect 16347 6205 16359 6208
rect 16301 6199 16359 6205
rect 16485 6205 16497 6208
rect 16531 6236 16543 6239
rect 17770 6236 17776 6248
rect 16531 6208 17776 6236
rect 16531 6205 16543 6208
rect 16485 6199 16543 6205
rect 10918 6171 10976 6177
rect 10918 6168 10930 6171
rect 10428 6140 10930 6168
rect 10918 6137 10930 6140
rect 10964 6168 10976 6171
rect 11606 6168 11612 6180
rect 10964 6140 11612 6168
rect 10964 6137 10976 6140
rect 10918 6131 10976 6137
rect 11606 6128 11612 6140
rect 11664 6168 11670 6180
rect 11793 6171 11851 6177
rect 11793 6168 11805 6171
rect 11664 6140 11805 6168
rect 11664 6128 11670 6140
rect 11793 6137 11805 6140
rect 11839 6168 11851 6171
rect 12161 6171 12219 6177
rect 12161 6168 12173 6171
rect 11839 6140 12173 6168
rect 11839 6137 11851 6140
rect 11793 6131 11851 6137
rect 12161 6137 12173 6140
rect 12207 6168 12219 6171
rect 12758 6171 12816 6177
rect 12758 6168 12770 6171
rect 12207 6140 12770 6168
rect 12207 6137 12219 6140
rect 12161 6131 12219 6137
rect 12758 6137 12770 6140
rect 12804 6137 12816 6171
rect 12758 6131 12816 6137
rect 7561 6103 7619 6109
rect 7561 6100 7573 6103
rect 7156 6072 7573 6100
rect 7156 6060 7162 6072
rect 7561 6069 7573 6072
rect 7607 6069 7619 6103
rect 7561 6063 7619 6069
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 9631 6103 9689 6109
rect 9631 6100 9643 6103
rect 9548 6072 9643 6100
rect 9548 6060 9554 6072
rect 9631 6069 9643 6072
rect 9677 6069 9689 6103
rect 10042 6100 10048 6112
rect 10003 6072 10048 6100
rect 9631 6063 9689 6069
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 14016 6100 14044 6199
rect 17770 6196 17776 6208
rect 17828 6196 17834 6248
rect 19426 6196 19432 6248
rect 19484 6196 19490 6248
rect 24578 6236 24584 6248
rect 24539 6208 24584 6236
rect 24578 6196 24584 6208
rect 24636 6236 24642 6248
rect 25133 6239 25191 6245
rect 25133 6236 25145 6239
rect 24636 6208 25145 6236
rect 24636 6196 24642 6208
rect 25133 6205 25145 6208
rect 25179 6205 25191 6239
rect 25133 6199 25191 6205
rect 14369 6171 14427 6177
rect 14369 6137 14381 6171
rect 14415 6137 14427 6171
rect 14369 6131 14427 6137
rect 14384 6100 14412 6131
rect 17954 6128 17960 6180
rect 18012 6168 18018 6180
rect 18141 6171 18199 6177
rect 18141 6168 18153 6171
rect 18012 6140 18153 6168
rect 18012 6128 18018 6140
rect 18141 6137 18153 6140
rect 18187 6137 18199 6171
rect 18141 6131 18199 6137
rect 18233 6171 18291 6177
rect 18233 6137 18245 6171
rect 18279 6137 18291 6171
rect 19444 6168 19472 6196
rect 19705 6171 19763 6177
rect 19705 6168 19717 6171
rect 19444 6140 19717 6168
rect 18233 6131 18291 6137
rect 19705 6137 19717 6140
rect 19751 6137 19763 6171
rect 19705 6131 19763 6137
rect 14016 6072 14412 6100
rect 17770 6060 17776 6112
rect 17828 6100 17834 6112
rect 18248 6100 18276 6131
rect 19794 6128 19800 6180
rect 19852 6168 19858 6180
rect 19852 6140 19897 6168
rect 19852 6128 19858 6140
rect 17828 6072 18276 6100
rect 17828 6060 17834 6072
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 5261 5899 5319 5905
rect 5261 5865 5273 5899
rect 5307 5896 5319 5899
rect 5534 5896 5540 5908
rect 5307 5868 5540 5896
rect 5307 5865 5319 5868
rect 5261 5859 5319 5865
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 8294 5896 8300 5908
rect 8255 5868 8300 5896
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8711 5899 8769 5905
rect 8711 5865 8723 5899
rect 8757 5896 8769 5899
rect 9030 5896 9036 5908
rect 8757 5868 9036 5896
rect 8757 5865 8769 5868
rect 8711 5859 8769 5865
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5896 9183 5899
rect 9214 5896 9220 5908
rect 9171 5868 9220 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9214 5856 9220 5868
rect 9272 5896 9278 5908
rect 10134 5896 10140 5908
rect 9272 5868 10140 5896
rect 9272 5856 9278 5868
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 11146 5856 11152 5908
rect 11204 5896 11210 5908
rect 11241 5899 11299 5905
rect 11241 5896 11253 5899
rect 11204 5868 11253 5896
rect 11204 5856 11210 5868
rect 11241 5865 11253 5868
rect 11287 5865 11299 5899
rect 12894 5896 12900 5908
rect 11241 5859 11299 5865
rect 12636 5868 12900 5896
rect 12636 5840 12664 5868
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 13170 5856 13176 5908
rect 13228 5856 13234 5908
rect 13998 5896 14004 5908
rect 13959 5868 14004 5896
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 14323 5899 14381 5905
rect 14323 5865 14335 5899
rect 14369 5896 14381 5899
rect 14826 5896 14832 5908
rect 14369 5868 14832 5896
rect 14369 5865 14381 5868
rect 14323 5859 14381 5865
rect 14826 5856 14832 5868
rect 14884 5856 14890 5908
rect 16850 5896 16856 5908
rect 16811 5868 16856 5896
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 7098 5837 7104 5840
rect 7095 5828 7104 5837
rect 7059 5800 7104 5828
rect 7095 5791 7104 5800
rect 7098 5788 7104 5791
rect 7156 5788 7162 5840
rect 8021 5831 8079 5837
rect 8021 5797 8033 5831
rect 8067 5828 8079 5831
rect 9398 5828 9404 5840
rect 8067 5800 9404 5828
rect 8067 5797 8079 5800
rect 8021 5791 8079 5797
rect 6178 5720 6184 5772
rect 6236 5760 6242 5772
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 6236 5732 6745 5760
rect 6236 5720 6242 5732
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 6733 5723 6791 5729
rect 7558 5720 7564 5772
rect 7616 5760 7622 5772
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 7616 5732 7665 5760
rect 7616 5720 7622 5732
rect 7653 5729 7665 5732
rect 7699 5760 7711 5763
rect 8036 5760 8064 5791
rect 9398 5788 9404 5800
rect 9456 5788 9462 5840
rect 9858 5828 9864 5840
rect 9819 5800 9864 5828
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 12618 5828 12624 5840
rect 12579 5800 12624 5828
rect 12618 5788 12624 5800
rect 12676 5788 12682 5840
rect 12713 5831 12771 5837
rect 12713 5797 12725 5831
rect 12759 5828 12771 5831
rect 13188 5828 13216 5856
rect 15286 5828 15292 5840
rect 12759 5800 13216 5828
rect 15247 5800 15292 5828
rect 12759 5797 12771 5800
rect 12713 5791 12771 5797
rect 15286 5788 15292 5800
rect 15344 5788 15350 5840
rect 17770 5828 17776 5840
rect 17731 5800 17776 5828
rect 17770 5788 17776 5800
rect 17828 5788 17834 5840
rect 19242 5788 19248 5840
rect 19300 5828 19306 5840
rect 19337 5831 19395 5837
rect 19337 5828 19349 5831
rect 19300 5800 19349 5828
rect 19300 5788 19306 5800
rect 19337 5797 19349 5800
rect 19383 5828 19395 5831
rect 20898 5828 20904 5840
rect 19383 5800 20904 5828
rect 19383 5797 19395 5800
rect 19337 5791 19395 5797
rect 20898 5788 20904 5800
rect 20956 5788 20962 5840
rect 8662 5769 8668 5772
rect 7699 5732 8064 5760
rect 8640 5763 8668 5769
rect 7699 5729 7711 5732
rect 7653 5723 7711 5729
rect 8640 5729 8652 5763
rect 8640 5723 8668 5729
rect 8662 5720 8668 5723
rect 8720 5720 8726 5772
rect 14252 5763 14310 5769
rect 14252 5729 14264 5763
rect 14298 5760 14310 5763
rect 14550 5760 14556 5772
rect 14298 5732 14556 5760
rect 14298 5729 14310 5732
rect 14252 5723 14310 5729
rect 14550 5720 14556 5732
rect 14608 5720 14614 5772
rect 15470 5760 15476 5772
rect 15431 5732 15476 5760
rect 15470 5720 15476 5732
rect 15528 5720 15534 5772
rect 9766 5692 9772 5704
rect 9727 5664 9772 5692
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 10045 5695 10103 5701
rect 10045 5661 10057 5695
rect 10091 5661 10103 5695
rect 10045 5655 10103 5661
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 10060 5624 10088 5655
rect 10962 5652 10968 5704
rect 11020 5692 11026 5704
rect 11425 5695 11483 5701
rect 11425 5692 11437 5695
rect 11020 5664 11437 5692
rect 11020 5652 11026 5664
rect 11425 5661 11437 5664
rect 11471 5661 11483 5695
rect 11425 5655 11483 5661
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 13630 5692 13636 5704
rect 13320 5664 13636 5692
rect 13320 5652 13326 5664
rect 13630 5652 13636 5664
rect 13688 5652 13694 5704
rect 16758 5652 16764 5704
rect 16816 5692 16822 5704
rect 17681 5695 17739 5701
rect 17681 5692 17693 5695
rect 16816 5664 17693 5692
rect 16816 5652 16822 5664
rect 17681 5661 17693 5664
rect 17727 5661 17739 5695
rect 17681 5655 17739 5661
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5692 18383 5695
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 18371 5664 19257 5692
rect 18371 5661 18383 5664
rect 18325 5655 18383 5661
rect 19245 5661 19257 5664
rect 19291 5692 19303 5695
rect 19334 5692 19340 5704
rect 19291 5664 19340 5692
rect 19291 5661 19303 5664
rect 19245 5655 19303 5661
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 19518 5692 19524 5704
rect 19479 5664 19524 5692
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 9732 5596 10088 5624
rect 10873 5627 10931 5633
rect 9732 5584 9738 5596
rect 10873 5593 10885 5627
rect 10919 5624 10931 5627
rect 11054 5624 11060 5636
rect 10919 5596 11060 5624
rect 10919 5593 10931 5596
rect 10873 5587 10931 5593
rect 11054 5584 11060 5596
rect 11112 5624 11118 5636
rect 11790 5624 11796 5636
rect 11112 5596 11796 5624
rect 11112 5584 11118 5596
rect 11790 5584 11796 5596
rect 11848 5584 11854 5636
rect 13078 5584 13084 5636
rect 13136 5624 13142 5636
rect 13173 5627 13231 5633
rect 13173 5624 13185 5627
rect 13136 5596 13185 5624
rect 13136 5584 13142 5596
rect 13173 5593 13185 5596
rect 13219 5624 13231 5627
rect 14274 5624 14280 5636
rect 13219 5596 14280 5624
rect 13219 5593 13231 5596
rect 13173 5587 13231 5593
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 17770 5516 17776 5568
rect 17828 5556 17834 5568
rect 18601 5559 18659 5565
rect 18601 5556 18613 5559
rect 17828 5528 18613 5556
rect 17828 5516 17834 5528
rect 18601 5525 18613 5528
rect 18647 5556 18659 5559
rect 18690 5556 18696 5568
rect 18647 5528 18696 5556
rect 18647 5525 18659 5528
rect 18601 5519 18659 5525
rect 18690 5516 18696 5528
rect 18748 5516 18754 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 6178 5352 6184 5364
rect 6139 5324 6184 5352
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 7098 5352 7104 5364
rect 7059 5324 7104 5352
rect 7098 5312 7104 5324
rect 7156 5312 7162 5364
rect 8662 5352 8668 5364
rect 8623 5324 8668 5352
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 9953 5355 10011 5361
rect 9953 5352 9965 5355
rect 9916 5324 9965 5352
rect 9916 5312 9922 5324
rect 9953 5321 9965 5324
rect 9999 5321 10011 5355
rect 11790 5352 11796 5364
rect 11751 5324 11796 5352
rect 9953 5315 10011 5321
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 13814 5352 13820 5364
rect 13775 5324 13820 5352
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 14550 5312 14556 5364
rect 14608 5352 14614 5364
rect 15013 5355 15071 5361
rect 15013 5352 15025 5355
rect 14608 5324 15025 5352
rect 14608 5312 14614 5324
rect 15013 5321 15025 5324
rect 15059 5321 15071 5355
rect 15470 5352 15476 5364
rect 15431 5324 15476 5352
rect 15013 5315 15071 5321
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 17083 5355 17141 5361
rect 17083 5321 17095 5355
rect 17129 5352 17141 5355
rect 17770 5352 17776 5364
rect 17129 5324 17776 5352
rect 17129 5321 17141 5324
rect 17083 5315 17141 5321
rect 17770 5312 17776 5324
rect 17828 5312 17834 5364
rect 19242 5352 19248 5364
rect 19203 5324 19248 5352
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19521 5355 19579 5361
rect 19521 5352 19533 5355
rect 19392 5324 19533 5352
rect 19392 5312 19398 5324
rect 19521 5321 19533 5324
rect 19567 5321 19579 5355
rect 19521 5315 19579 5321
rect 23474 5312 23480 5364
rect 23532 5352 23538 5364
rect 24719 5355 24777 5361
rect 24719 5352 24731 5355
rect 23532 5324 24731 5352
rect 23532 5312 23538 5324
rect 24719 5321 24731 5324
rect 24765 5321 24777 5355
rect 24719 5315 24777 5321
rect 9398 5244 9404 5296
rect 9456 5284 9462 5296
rect 9582 5284 9588 5296
rect 9456 5256 9588 5284
rect 9456 5244 9462 5256
rect 9582 5244 9588 5256
rect 9640 5244 9646 5296
rect 12069 5287 12127 5293
rect 12069 5253 12081 5287
rect 12115 5284 12127 5287
rect 12618 5284 12624 5296
rect 12115 5256 12624 5284
rect 12115 5253 12127 5256
rect 12069 5247 12127 5253
rect 12618 5244 12624 5256
rect 12676 5244 12682 5296
rect 13078 5284 13084 5296
rect 13039 5256 13084 5284
rect 13078 5244 13084 5256
rect 13136 5244 13142 5296
rect 13998 5244 14004 5296
rect 14056 5244 14062 5296
rect 9033 5219 9091 5225
rect 9033 5185 9045 5219
rect 9079 5216 9091 5219
rect 9214 5216 9220 5228
rect 9079 5188 9220 5216
rect 9079 5185 9091 5188
rect 9033 5179 9091 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5216 10747 5219
rect 10873 5219 10931 5225
rect 10873 5216 10885 5219
rect 10735 5188 10885 5216
rect 10735 5185 10747 5188
rect 10689 5179 10747 5185
rect 10873 5185 10885 5188
rect 10919 5216 10931 5219
rect 10962 5216 10968 5228
rect 10919 5188 10968 5216
rect 10919 5185 10931 5188
rect 10873 5179 10931 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 12526 5216 12532 5228
rect 12439 5188 12532 5216
rect 12526 5176 12532 5188
rect 12584 5216 12590 5228
rect 13449 5219 13507 5225
rect 13449 5216 13461 5219
rect 12584 5188 13461 5216
rect 12584 5176 12590 5188
rect 13449 5185 13461 5188
rect 13495 5185 13507 5219
rect 14016 5216 14044 5244
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 14016 5188 14105 5216
rect 13449 5179 13507 5185
rect 14093 5185 14105 5188
rect 14139 5185 14151 5219
rect 14366 5216 14372 5228
rect 14327 5188 14372 5216
rect 14093 5179 14151 5185
rect 14366 5176 14372 5188
rect 14424 5216 14430 5228
rect 14424 5188 14964 5216
rect 14424 5176 14430 5188
rect 14936 5148 14964 5188
rect 17126 5176 17132 5228
rect 17184 5216 17190 5228
rect 17405 5219 17463 5225
rect 17405 5216 17417 5219
rect 17184 5188 17417 5216
rect 17184 5176 17190 5188
rect 17405 5185 17417 5188
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 17773 5219 17831 5225
rect 17773 5216 17785 5219
rect 17736 5188 17785 5216
rect 17736 5176 17742 5188
rect 17773 5185 17785 5188
rect 17819 5185 17831 5219
rect 17773 5179 17831 5185
rect 18049 5219 18107 5225
rect 18049 5185 18061 5219
rect 18095 5216 18107 5219
rect 19426 5216 19432 5228
rect 18095 5188 19432 5216
rect 18095 5185 18107 5188
rect 18049 5179 18107 5185
rect 19426 5176 19432 5188
rect 19484 5176 19490 5228
rect 15600 5151 15658 5157
rect 15600 5148 15612 5151
rect 14936 5120 15612 5148
rect 15600 5117 15612 5120
rect 15646 5148 15658 5151
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 15646 5120 16037 5148
rect 15646 5117 15658 5120
rect 15600 5111 15658 5117
rect 16025 5117 16037 5120
rect 16071 5117 16083 5151
rect 16025 5111 16083 5117
rect 17012 5151 17070 5157
rect 17012 5117 17024 5151
rect 17058 5148 17070 5151
rect 17144 5148 17172 5176
rect 17058 5120 17172 5148
rect 24648 5151 24706 5157
rect 17058 5117 17070 5120
rect 17012 5111 17070 5117
rect 24648 5117 24660 5151
rect 24694 5148 24706 5151
rect 24694 5120 25176 5148
rect 24694 5117 24706 5120
rect 24648 5111 24706 5117
rect 6362 5040 6368 5092
rect 6420 5080 6426 5092
rect 6641 5083 6699 5089
rect 6641 5080 6653 5083
rect 6420 5052 6653 5080
rect 6420 5040 6426 5052
rect 6641 5049 6653 5052
rect 6687 5080 6699 5083
rect 7469 5083 7527 5089
rect 7469 5080 7481 5083
rect 6687 5052 7481 5080
rect 6687 5049 6699 5052
rect 6641 5043 6699 5049
rect 7469 5049 7481 5052
rect 7515 5049 7527 5083
rect 7469 5043 7527 5049
rect 7558 5040 7564 5092
rect 7616 5080 7622 5092
rect 8110 5080 8116 5092
rect 7616 5052 7661 5080
rect 8071 5052 8116 5080
rect 7616 5040 7622 5052
rect 8110 5040 8116 5052
rect 8168 5040 8174 5092
rect 9122 5040 9128 5092
rect 9180 5080 9186 5092
rect 10965 5083 11023 5089
rect 9180 5052 9225 5080
rect 9180 5040 9186 5052
rect 10965 5049 10977 5083
rect 11011 5080 11023 5083
rect 11054 5080 11060 5092
rect 11011 5052 11060 5080
rect 11011 5049 11023 5052
rect 10965 5043 11023 5049
rect 11054 5040 11060 5052
rect 11112 5040 11118 5092
rect 11514 5080 11520 5092
rect 11475 5052 11520 5080
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 11974 5040 11980 5092
rect 12032 5080 12038 5092
rect 12526 5080 12532 5092
rect 12032 5052 12532 5080
rect 12032 5040 12038 5052
rect 12526 5040 12532 5052
rect 12584 5040 12590 5092
rect 12618 5040 12624 5092
rect 12676 5080 12682 5092
rect 14185 5083 14243 5089
rect 12676 5052 12721 5080
rect 12676 5040 12682 5052
rect 14185 5049 14197 5083
rect 14231 5049 14243 5083
rect 14185 5043 14243 5049
rect 10870 4972 10876 5024
rect 10928 5012 10934 5024
rect 11330 5012 11336 5024
rect 10928 4984 11336 5012
rect 10928 4972 10934 4984
rect 11330 4972 11336 4984
rect 11388 5012 11394 5024
rect 12069 5015 12127 5021
rect 12069 5012 12081 5015
rect 11388 4984 12081 5012
rect 11388 4972 11394 4984
rect 12069 4981 12081 4984
rect 12115 5012 12127 5015
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 12115 4984 12173 5012
rect 12115 4981 12127 4984
rect 12069 4975 12127 4981
rect 12161 4981 12173 4984
rect 12207 4981 12219 5015
rect 12161 4975 12219 4981
rect 13814 4972 13820 5024
rect 13872 5012 13878 5024
rect 14200 5012 14228 5043
rect 25148 5024 25176 5120
rect 15746 5021 15752 5024
rect 13872 4984 14228 5012
rect 15703 5015 15752 5021
rect 13872 4972 13878 4984
rect 15703 4981 15715 5015
rect 15749 4981 15752 5015
rect 15703 4975 15752 4981
rect 15746 4972 15752 4975
rect 15804 4972 15810 5024
rect 16758 5012 16764 5024
rect 16719 4984 16764 5012
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 25130 5012 25136 5024
rect 25091 4984 25136 5012
rect 25130 4972 25136 4984
rect 25188 4972 25194 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 6362 4808 6368 4820
rect 6323 4780 6368 4808
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 9033 4811 9091 4817
rect 9033 4777 9045 4811
rect 9079 4808 9091 4811
rect 9122 4808 9128 4820
rect 9079 4780 9128 4808
rect 9079 4777 9091 4780
rect 9033 4771 9091 4777
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 10137 4811 10195 4817
rect 10137 4808 10149 4811
rect 9824 4780 10149 4808
rect 9824 4768 9830 4780
rect 10137 4777 10149 4780
rect 10183 4777 10195 4811
rect 10137 4771 10195 4777
rect 12894 4768 12900 4820
rect 12952 4808 12958 4820
rect 17862 4817 17868 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 12952 4780 13277 4808
rect 12952 4768 12958 4780
rect 13265 4777 13277 4780
rect 13311 4777 13323 4811
rect 13265 4771 13323 4777
rect 17819 4811 17868 4817
rect 17819 4777 17831 4811
rect 17865 4777 17868 4811
rect 17819 4771 17868 4777
rect 17862 4768 17868 4771
rect 17920 4768 17926 4820
rect 24762 4808 24768 4820
rect 24723 4780 24768 4808
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 7558 4740 7564 4752
rect 7519 4712 7564 4740
rect 7558 4700 7564 4712
rect 7616 4700 7622 4752
rect 8113 4743 8171 4749
rect 8113 4709 8125 4743
rect 8159 4740 8171 4743
rect 8202 4740 8208 4752
rect 8159 4712 8208 4740
rect 8159 4709 8171 4712
rect 8113 4703 8171 4709
rect 8202 4700 8208 4712
rect 8260 4700 8266 4752
rect 10870 4740 10876 4752
rect 10831 4712 10876 4740
rect 10870 4700 10876 4712
rect 10928 4700 10934 4752
rect 11425 4743 11483 4749
rect 11425 4709 11437 4743
rect 11471 4740 11483 4743
rect 11514 4740 11520 4752
rect 11471 4712 11520 4740
rect 11471 4709 11483 4712
rect 11425 4703 11483 4709
rect 11514 4700 11520 4712
rect 11572 4700 11578 4752
rect 12066 4700 12072 4752
rect 12124 4740 12130 4752
rect 12342 4740 12348 4752
rect 12124 4712 12348 4740
rect 12124 4700 12130 4712
rect 12342 4700 12348 4712
rect 12400 4740 12406 4752
rect 12437 4743 12495 4749
rect 12437 4740 12449 4743
rect 12400 4712 12449 4740
rect 12400 4700 12406 4712
rect 12437 4709 12449 4712
rect 12483 4709 12495 4743
rect 12437 4703 12495 4709
rect 12989 4743 13047 4749
rect 12989 4709 13001 4743
rect 13035 4740 13047 4743
rect 13078 4740 13084 4752
rect 13035 4712 13084 4740
rect 13035 4709 13047 4712
rect 12989 4703 13047 4709
rect 13078 4700 13084 4712
rect 13136 4700 13142 4752
rect 9744 4675 9802 4681
rect 9744 4641 9756 4675
rect 9790 4672 9802 4675
rect 9858 4672 9864 4684
rect 9790 4644 9864 4672
rect 9790 4641 9802 4644
rect 9744 4635 9802 4641
rect 9858 4632 9864 4644
rect 9916 4672 9922 4684
rect 10594 4672 10600 4684
rect 9916 4644 10600 4672
rect 9916 4632 9922 4644
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 13868 4675 13926 4681
rect 13868 4641 13880 4675
rect 13914 4672 13926 4675
rect 14182 4672 14188 4684
rect 13914 4644 14188 4672
rect 13914 4641 13926 4644
rect 13868 4635 13926 4641
rect 14182 4632 14188 4644
rect 14240 4632 14246 4684
rect 15746 4672 15752 4684
rect 15707 4644 15752 4672
rect 15746 4632 15752 4644
rect 15804 4632 15810 4684
rect 17586 4632 17592 4684
rect 17644 4672 17650 4684
rect 17716 4675 17774 4681
rect 17716 4672 17728 4675
rect 17644 4644 17728 4672
rect 17644 4632 17650 4644
rect 17716 4641 17728 4644
rect 17762 4641 17774 4675
rect 17716 4635 17774 4641
rect 24210 4632 24216 4684
rect 24268 4672 24274 4684
rect 24581 4675 24639 4681
rect 24581 4672 24593 4675
rect 24268 4644 24593 4672
rect 24268 4632 24274 4644
rect 24581 4641 24593 4644
rect 24627 4641 24639 4675
rect 24581 4635 24639 4641
rect 7190 4564 7196 4616
rect 7248 4604 7254 4616
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 7248 4576 7481 4604
rect 7248 4564 7254 4576
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 10134 4564 10140 4616
rect 10192 4604 10198 4616
rect 10781 4607 10839 4613
rect 10781 4604 10793 4607
rect 10192 4576 10793 4604
rect 10192 4564 10198 4576
rect 10781 4573 10793 4576
rect 10827 4573 10839 4607
rect 12342 4604 12348 4616
rect 12303 4576 12348 4604
rect 10781 4567 10839 4573
rect 12342 4564 12348 4576
rect 12400 4604 12406 4616
rect 13955 4607 14013 4613
rect 13955 4604 13967 4607
rect 12400 4576 13967 4604
rect 12400 4564 12406 4576
rect 13955 4573 13967 4576
rect 14001 4573 14013 4607
rect 13955 4567 14013 4573
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 9815 4471 9873 4477
rect 9815 4468 9827 4471
rect 9732 4440 9827 4468
rect 9732 4428 9738 4440
rect 9815 4437 9827 4440
rect 9861 4437 9873 4471
rect 15930 4468 15936 4480
rect 15891 4440 15936 4468
rect 9815 4431 9873 4437
rect 15930 4428 15936 4440
rect 15988 4428 15994 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 7558 4264 7564 4276
rect 7116 4236 7564 4264
rect 7116 4196 7144 4236
rect 7558 4224 7564 4236
rect 7616 4224 7622 4276
rect 9858 4264 9864 4276
rect 9819 4236 9864 4264
rect 9858 4224 9864 4236
rect 9916 4224 9922 4276
rect 10689 4267 10747 4273
rect 10689 4233 10701 4267
rect 10735 4264 10747 4267
rect 10870 4264 10876 4276
rect 10735 4236 10876 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 11885 4267 11943 4273
rect 11885 4233 11897 4267
rect 11931 4264 11943 4267
rect 12342 4264 12348 4276
rect 11931 4236 12348 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 12342 4224 12348 4236
rect 12400 4224 12406 4276
rect 13909 4267 13967 4273
rect 13909 4233 13921 4267
rect 13955 4264 13967 4267
rect 14182 4264 14188 4276
rect 13955 4236 14188 4264
rect 13955 4233 13967 4236
rect 13909 4227 13967 4233
rect 14182 4224 14188 4236
rect 14240 4264 14246 4276
rect 15746 4264 15752 4276
rect 14240 4236 15056 4264
rect 15707 4236 15752 4264
rect 14240 4224 14246 4236
rect 6932 4168 7144 4196
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6932 4128 6960 4168
rect 7190 4156 7196 4208
rect 7248 4196 7254 4208
rect 7248 4168 8248 4196
rect 7248 4156 7254 4168
rect 6687 4100 6960 4128
rect 8021 4131 8079 4137
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8110 4128 8116 4140
rect 8067 4100 8116 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8220 4128 8248 4168
rect 9214 4156 9220 4208
rect 9272 4196 9278 4208
rect 9493 4199 9551 4205
rect 9493 4196 9505 4199
rect 9272 4168 9505 4196
rect 9272 4156 9278 4168
rect 9493 4165 9505 4168
rect 9539 4165 9551 4199
rect 14366 4196 14372 4208
rect 9493 4159 9551 4165
rect 13740 4168 14372 4196
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8220 4100 8309 4128
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8570 4088 8576 4140
rect 8628 4128 8634 4140
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 8628 4100 8677 4128
rect 8628 4088 8634 4100
rect 8665 4097 8677 4100
rect 8711 4097 8723 4131
rect 8938 4128 8944 4140
rect 8851 4100 8944 4128
rect 8665 4091 8723 4097
rect 7374 3992 7380 4004
rect 7335 3964 7380 3992
rect 7374 3952 7380 3964
rect 7432 3952 7438 4004
rect 7469 3995 7527 4001
rect 7469 3961 7481 3995
rect 7515 3992 7527 3995
rect 8680 3992 8708 4091
rect 8938 4088 8944 4100
rect 8996 4128 9002 4140
rect 9582 4128 9588 4140
rect 8996 4100 9588 4128
rect 8996 4088 9002 4100
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 11514 4128 11520 4140
rect 11475 4100 11520 4128
rect 11514 4088 11520 4100
rect 11572 4128 11578 4140
rect 12526 4128 12532 4140
rect 11572 4100 12532 4128
rect 11572 4088 11578 4100
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 13173 4131 13231 4137
rect 13173 4097 13185 4131
rect 13219 4128 13231 4131
rect 13740 4128 13768 4168
rect 14366 4156 14372 4168
rect 14424 4156 14430 4208
rect 15028 4196 15056 4236
rect 15746 4224 15752 4236
rect 15804 4224 15810 4276
rect 17586 4224 17592 4276
rect 17644 4264 17650 4276
rect 17681 4267 17739 4273
rect 17681 4264 17693 4267
rect 17644 4236 17693 4264
rect 17644 4224 17650 4236
rect 17681 4233 17693 4236
rect 17727 4233 17739 4267
rect 17681 4227 17739 4233
rect 24210 4224 24216 4276
rect 24268 4264 24274 4276
rect 24581 4267 24639 4273
rect 24581 4264 24593 4267
rect 24268 4236 24593 4264
rect 24268 4224 24274 4236
rect 24581 4233 24593 4236
rect 24627 4233 24639 4267
rect 24581 4227 24639 4233
rect 16114 4196 16120 4208
rect 15028 4168 16120 4196
rect 16114 4156 16120 4168
rect 16172 4156 16178 4208
rect 13219 4100 13768 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 12066 4020 12072 4072
rect 12124 4060 12130 4072
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 12124 4032 12173 4060
rect 12124 4020 12130 4032
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 14436 4063 14494 4069
rect 14436 4029 14448 4063
rect 14482 4060 14494 4063
rect 14482 4032 14964 4060
rect 14482 4029 14494 4032
rect 14436 4023 14494 4029
rect 9033 3995 9091 4001
rect 9033 3992 9045 3995
rect 7515 3964 9045 3992
rect 7515 3961 7527 3964
rect 7469 3955 7527 3961
rect 9033 3961 9045 3964
rect 9079 3961 9091 3995
rect 9033 3955 9091 3961
rect 7193 3927 7251 3933
rect 7193 3893 7205 3927
rect 7239 3924 7251 3927
rect 7484 3924 7512 3955
rect 10042 3952 10048 4004
rect 10100 3992 10106 4004
rect 10870 3992 10876 4004
rect 10100 3964 10876 3992
rect 10100 3952 10106 3964
rect 10870 3952 10876 3964
rect 10928 3952 10934 4004
rect 10962 3952 10968 4004
rect 11020 3992 11026 4004
rect 12084 3992 12112 4020
rect 12526 3992 12532 4004
rect 11020 3964 12112 3992
rect 12487 3964 12532 3992
rect 11020 3952 11026 3964
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 12621 3995 12679 4001
rect 12621 3961 12633 3995
rect 12667 3961 12679 3995
rect 12621 3955 12679 3961
rect 7239 3896 7512 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 10192 3896 10241 3924
rect 10192 3884 10198 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 10229 3887 10287 3893
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12636 3924 12664 3955
rect 14936 3936 14964 4032
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 20257 4063 20315 4069
rect 20257 4060 20269 4063
rect 19484 4032 20269 4060
rect 19484 4020 19490 4032
rect 20257 4029 20269 4032
rect 20303 4060 20315 4063
rect 20809 4063 20867 4069
rect 20809 4060 20821 4063
rect 20303 4032 20821 4060
rect 20303 4029 20315 4032
rect 20257 4023 20315 4029
rect 20809 4029 20821 4032
rect 20855 4029 20867 4063
rect 20809 4023 20867 4029
rect 12492 3896 12664 3924
rect 14507 3927 14565 3933
rect 12492 3884 12498 3896
rect 14507 3893 14519 3927
rect 14553 3924 14565 3927
rect 14734 3924 14740 3936
rect 14553 3896 14740 3924
rect 14553 3893 14565 3896
rect 14507 3887 14565 3893
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 14918 3924 14924 3936
rect 14879 3896 14924 3924
rect 14918 3884 14924 3896
rect 14976 3884 14982 3936
rect 20438 3924 20444 3936
rect 20399 3896 20444 3924
rect 20438 3884 20444 3896
rect 20496 3884 20502 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 2363 3723 2421 3729
rect 2363 3689 2375 3723
rect 2409 3720 2421 3723
rect 2682 3720 2688 3732
rect 2409 3692 2688 3720
rect 2409 3689 2421 3692
rect 2363 3683 2421 3689
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 5442 3680 5448 3732
rect 5500 3729 5506 3732
rect 5500 3723 5549 3729
rect 5500 3689 5503 3723
rect 5537 3689 5549 3723
rect 5500 3683 5549 3689
rect 6503 3723 6561 3729
rect 6503 3689 6515 3723
rect 6549 3720 6561 3723
rect 7285 3723 7343 3729
rect 7285 3720 7297 3723
rect 6549 3692 7297 3720
rect 6549 3689 6561 3692
rect 6503 3683 6561 3689
rect 7285 3689 7297 3692
rect 7331 3720 7343 3723
rect 7374 3720 7380 3732
rect 7331 3692 7380 3720
rect 7331 3689 7343 3692
rect 7285 3683 7343 3689
rect 5500 3680 5506 3683
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 8938 3720 8944 3732
rect 8899 3692 8944 3720
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 11149 3723 11207 3729
rect 11149 3720 11161 3723
rect 10928 3692 11161 3720
rect 10928 3680 10934 3692
rect 11149 3689 11161 3692
rect 11195 3689 11207 3723
rect 11149 3683 11207 3689
rect 11839 3723 11897 3729
rect 11839 3689 11851 3723
rect 11885 3720 11897 3723
rect 11974 3720 11980 3732
rect 11885 3692 11980 3720
rect 11885 3689 11897 3692
rect 11839 3683 11897 3689
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 12492 3692 12537 3720
rect 12492 3680 12498 3692
rect 7561 3655 7619 3661
rect 7561 3621 7573 3655
rect 7607 3652 7619 3655
rect 7742 3652 7748 3664
rect 7607 3624 7748 3652
rect 7607 3621 7619 3624
rect 7561 3615 7619 3621
rect 7742 3612 7748 3624
rect 7800 3612 7806 3664
rect 8110 3652 8116 3664
rect 8071 3624 8116 3652
rect 8110 3612 8116 3624
rect 8168 3612 8174 3664
rect 9490 3612 9496 3664
rect 9548 3652 9554 3664
rect 9766 3652 9772 3664
rect 9548 3624 9772 3652
rect 9548 3612 9554 3624
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 9858 3612 9864 3664
rect 9916 3652 9922 3664
rect 9916 3624 9961 3652
rect 9916 3612 9922 3624
rect 12526 3612 12532 3664
rect 12584 3652 12590 3664
rect 12805 3655 12863 3661
rect 12805 3652 12817 3655
rect 12584 3624 12817 3652
rect 12584 3612 12590 3624
rect 12805 3621 12817 3624
rect 12851 3621 12863 3655
rect 12805 3615 12863 3621
rect 2292 3587 2350 3593
rect 2292 3553 2304 3587
rect 2338 3584 2350 3587
rect 2498 3584 2504 3596
rect 2338 3556 2504 3584
rect 2338 3553 2350 3556
rect 2292 3547 2350 3553
rect 2498 3544 2504 3556
rect 2556 3544 2562 3596
rect 5442 3593 5448 3596
rect 5420 3587 5448 3593
rect 5420 3553 5432 3587
rect 5420 3547 5448 3553
rect 5442 3544 5448 3547
rect 5500 3544 5506 3596
rect 6362 3544 6368 3596
rect 6420 3593 6426 3596
rect 6420 3587 6458 3593
rect 6446 3553 6458 3587
rect 6420 3547 6458 3553
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3584 10931 3587
rect 10962 3584 10968 3596
rect 10919 3556 10968 3584
rect 10919 3553 10931 3556
rect 10873 3547 10931 3553
rect 6420 3544 6426 3547
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11790 3593 11796 3596
rect 11768 3587 11796 3593
rect 11768 3553 11780 3587
rect 11768 3547 11796 3553
rect 11790 3544 11796 3547
rect 11848 3544 11854 3596
rect 21266 3544 21272 3596
rect 21324 3584 21330 3596
rect 21637 3587 21695 3593
rect 21637 3584 21649 3587
rect 21324 3556 21649 3584
rect 21324 3544 21330 3556
rect 21637 3553 21649 3556
rect 21683 3584 21695 3587
rect 22094 3584 22100 3596
rect 21683 3556 22100 3584
rect 21683 3553 21695 3556
rect 21637 3547 21695 3553
rect 22094 3544 22100 3556
rect 22152 3544 22158 3596
rect 7466 3516 7472 3528
rect 7427 3488 7472 3516
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 9214 3476 9220 3528
rect 9272 3516 9278 3528
rect 10045 3519 10103 3525
rect 10045 3516 10057 3519
rect 9272 3488 10057 3516
rect 9272 3476 9278 3488
rect 10045 3485 10057 3488
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 21818 3448 21824 3460
rect 21779 3420 21824 3448
rect 21818 3408 21824 3420
rect 21876 3408 21882 3460
rect 12894 3340 12900 3392
rect 12952 3380 12958 3392
rect 15378 3380 15384 3392
rect 12952 3352 15384 3380
rect 12952 3340 12958 3352
rect 15378 3340 15384 3352
rect 15436 3340 15442 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 6963 3179 7021 3185
rect 6963 3145 6975 3179
rect 7009 3176 7021 3179
rect 7466 3176 7472 3188
rect 7009 3148 7472 3176
rect 7009 3145 7021 3148
rect 6963 3139 7021 3145
rect 7466 3136 7472 3148
rect 7524 3176 7530 3188
rect 8021 3179 8079 3185
rect 8021 3176 8033 3179
rect 7524 3148 8033 3176
rect 7524 3136 7530 3148
rect 8021 3145 8033 3148
rect 8067 3145 8079 3179
rect 8021 3139 8079 3145
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 9493 3179 9551 3185
rect 9493 3176 9505 3179
rect 9456 3148 9505 3176
rect 9456 3136 9462 3148
rect 9493 3145 9505 3148
rect 9539 3145 9551 3179
rect 9493 3139 9551 3145
rect 7742 3108 7748 3120
rect 7703 3080 7748 3108
rect 7742 3068 7748 3080
rect 7800 3068 7806 3120
rect 6638 2932 6644 2984
rect 6696 2972 6702 2984
rect 6892 2975 6950 2981
rect 6892 2972 6904 2975
rect 6696 2944 6904 2972
rect 6696 2932 6702 2944
rect 6892 2941 6904 2944
rect 6938 2972 6950 2975
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 6938 2944 7297 2972
rect 6938 2941 6950 2944
rect 6892 2935 6950 2941
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 9508 2972 9536 3139
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 10505 3179 10563 3185
rect 10505 3176 10517 3179
rect 9824 3148 10517 3176
rect 9824 3136 9830 3148
rect 10505 3145 10517 3148
rect 10551 3145 10563 3179
rect 11790 3176 11796 3188
rect 11751 3148 11796 3176
rect 10505 3139 10563 3145
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 21726 3176 21732 3188
rect 21687 3148 21732 3176
rect 21726 3136 21732 3148
rect 21784 3136 21790 3188
rect 22094 3176 22100 3188
rect 22055 3148 22100 3176
rect 22094 3136 22100 3148
rect 22152 3136 22158 3188
rect 9858 3068 9864 3120
rect 9916 3108 9922 3120
rect 10137 3111 10195 3117
rect 10137 3108 10149 3111
rect 9916 3080 10149 3108
rect 9916 3068 9922 3080
rect 10137 3077 10149 3080
rect 10183 3077 10195 3111
rect 10137 3071 10195 3077
rect 18233 3111 18291 3117
rect 18233 3077 18245 3111
rect 18279 3108 18291 3111
rect 20070 3108 20076 3120
rect 18279 3080 20076 3108
rect 18279 3077 18291 3080
rect 18233 3071 18291 3077
rect 20070 3068 20076 3080
rect 20128 3068 20134 3120
rect 9712 2975 9770 2981
rect 9712 2972 9724 2975
rect 9508 2944 9724 2972
rect 7285 2935 7343 2941
rect 9712 2941 9724 2944
rect 9758 2941 9770 2975
rect 9712 2935 9770 2941
rect 12710 2932 12716 2984
rect 12768 2972 12774 2984
rect 13576 2975 13634 2981
rect 13576 2972 13588 2975
rect 12768 2944 13588 2972
rect 12768 2932 12774 2944
rect 13576 2941 13588 2944
rect 13622 2972 13634 2975
rect 14001 2975 14059 2981
rect 14001 2972 14013 2975
rect 13622 2944 14013 2972
rect 13622 2941 13634 2944
rect 13576 2935 13634 2941
rect 14001 2941 14013 2944
rect 14047 2941 14059 2975
rect 14001 2935 14059 2941
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 18012 2944 18061 2972
rect 18012 2932 18018 2944
rect 18049 2941 18061 2944
rect 18095 2972 18107 2975
rect 18601 2975 18659 2981
rect 18601 2972 18613 2975
rect 18095 2944 18613 2972
rect 18095 2941 18107 2944
rect 18049 2935 18107 2941
rect 18601 2941 18613 2944
rect 18647 2941 18659 2975
rect 18601 2935 18659 2941
rect 21177 2975 21235 2981
rect 21177 2941 21189 2975
rect 21223 2972 21235 2975
rect 21726 2972 21732 2984
rect 21223 2944 21732 2972
rect 21223 2941 21235 2944
rect 21177 2935 21235 2941
rect 21726 2932 21732 2944
rect 21784 2932 21790 2984
rect 24302 2972 24308 2984
rect 24263 2944 24308 2972
rect 24302 2932 24308 2944
rect 24360 2972 24366 2984
rect 24857 2975 24915 2981
rect 24857 2972 24869 2975
rect 24360 2944 24869 2972
rect 24360 2932 24366 2944
rect 24857 2941 24869 2944
rect 24903 2941 24915 2975
rect 24857 2935 24915 2941
rect 9815 2907 9873 2913
rect 9815 2873 9827 2907
rect 9861 2904 9873 2907
rect 10962 2904 10968 2916
rect 9861 2876 10968 2904
rect 9861 2873 9873 2876
rect 9815 2867 9873 2873
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 13722 2913 13728 2916
rect 13679 2907 13728 2913
rect 13679 2873 13691 2907
rect 13725 2873 13728 2907
rect 13679 2867 13728 2873
rect 13722 2864 13728 2867
rect 13780 2864 13786 2916
rect 2317 2839 2375 2845
rect 2317 2805 2329 2839
rect 2363 2836 2375 2839
rect 2498 2836 2504 2848
rect 2363 2808 2504 2836
rect 2363 2805 2375 2808
rect 2317 2799 2375 2805
rect 2498 2796 2504 2808
rect 2556 2796 2562 2848
rect 5442 2836 5448 2848
rect 5403 2808 5448 2836
rect 5442 2796 5448 2808
rect 5500 2796 5506 2848
rect 6362 2836 6368 2848
rect 6323 2808 6368 2836
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 21361 2839 21419 2845
rect 21361 2805 21373 2839
rect 21407 2836 21419 2839
rect 23198 2836 23204 2848
rect 21407 2808 23204 2836
rect 21407 2805 21419 2808
rect 21361 2799 21419 2805
rect 23198 2796 23204 2808
rect 23256 2796 23262 2848
rect 24486 2836 24492 2848
rect 24447 2808 24492 2836
rect 24486 2796 24492 2808
rect 24544 2796 24550 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1578 2641 1584 2644
rect 1535 2635 1584 2641
rect 1535 2601 1547 2635
rect 1581 2601 1584 2635
rect 1535 2595 1584 2601
rect 1578 2592 1584 2595
rect 1636 2592 1642 2644
rect 4614 2641 4620 2644
rect 4571 2635 4620 2641
rect 4571 2601 4583 2635
rect 4617 2601 4620 2635
rect 4571 2595 4620 2601
rect 4614 2592 4620 2595
rect 4672 2592 4678 2644
rect 7147 2635 7205 2641
rect 7147 2601 7159 2635
rect 7193 2632 7205 2635
rect 7374 2632 7380 2644
rect 7193 2604 7380 2632
rect 7193 2601 7205 2604
rect 7147 2595 7205 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 9950 2592 9956 2644
rect 10008 2641 10014 2644
rect 10008 2635 10057 2641
rect 10008 2601 10011 2635
rect 10045 2601 10057 2635
rect 10008 2595 10057 2601
rect 10008 2592 10014 2595
rect 10778 2592 10784 2644
rect 10836 2632 10842 2644
rect 16758 2641 16764 2644
rect 11011 2635 11069 2641
rect 11011 2632 11023 2635
rect 10836 2604 11023 2632
rect 10836 2592 10842 2604
rect 11011 2601 11023 2604
rect 11057 2601 11069 2635
rect 11011 2595 11069 2601
rect 16715 2635 16764 2641
rect 16715 2601 16727 2635
rect 16761 2601 16764 2635
rect 16715 2595 16764 2601
rect 16758 2592 16764 2595
rect 16816 2592 16822 2644
rect 18966 2632 18972 2644
rect 18927 2604 18972 2632
rect 18966 2592 18972 2604
rect 19024 2592 19030 2644
rect 20073 2635 20131 2641
rect 20073 2601 20085 2635
rect 20119 2632 20131 2635
rect 20254 2632 20260 2644
rect 20119 2604 20260 2632
rect 20119 2601 20131 2604
rect 20073 2595 20131 2601
rect 1394 2456 1400 2508
rect 1452 2505 1458 2508
rect 1452 2499 1490 2505
rect 1478 2496 1490 2499
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1478 2468 1869 2496
rect 1478 2465 1490 2468
rect 1452 2459 1490 2465
rect 1857 2465 1869 2468
rect 1903 2465 1915 2499
rect 1857 2459 1915 2465
rect 4500 2499 4558 2505
rect 4500 2465 4512 2499
rect 4546 2496 4558 2499
rect 7076 2499 7134 2505
rect 4546 2468 4660 2496
rect 4546 2465 4558 2468
rect 4500 2459 4558 2465
rect 1452 2456 1458 2459
rect 4632 2440 4660 2468
rect 7076 2465 7088 2499
rect 7122 2496 7134 2499
rect 7122 2468 7604 2496
rect 7122 2465 7134 2468
rect 7076 2459 7134 2465
rect 4614 2388 4620 2440
rect 4672 2428 4678 2440
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 4672 2400 4905 2428
rect 4672 2388 4678 2400
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 7576 2301 7604 2468
rect 9858 2456 9864 2508
rect 9916 2505 9922 2508
rect 9916 2499 9954 2505
rect 9942 2496 9954 2499
rect 10321 2499 10379 2505
rect 10321 2496 10333 2499
rect 9942 2468 10333 2496
rect 9942 2465 9954 2468
rect 9916 2459 9954 2465
rect 10321 2465 10333 2468
rect 10367 2465 10379 2499
rect 10321 2459 10379 2465
rect 10940 2499 10998 2505
rect 10940 2465 10952 2499
rect 10986 2496 10998 2499
rect 16644 2499 16702 2505
rect 10986 2468 11468 2496
rect 10986 2465 10998 2468
rect 10940 2459 10998 2465
rect 9916 2456 9922 2459
rect 7561 2295 7619 2301
rect 7561 2261 7573 2295
rect 7607 2292 7619 2295
rect 7650 2292 7656 2304
rect 7607 2264 7656 2292
rect 7607 2261 7619 2264
rect 7561 2255 7619 2261
rect 7650 2252 7656 2264
rect 7708 2252 7714 2304
rect 11440 2301 11468 2468
rect 16644 2465 16656 2499
rect 16690 2496 16702 2499
rect 17034 2496 17040 2508
rect 16690 2468 17040 2496
rect 16690 2465 16702 2468
rect 16644 2459 16702 2465
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2496 18383 2499
rect 18984 2496 19012 2592
rect 18371 2468 19012 2496
rect 19429 2499 19487 2505
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 19429 2465 19441 2499
rect 19475 2496 19487 2499
rect 20088 2496 20116 2595
rect 20254 2592 20260 2604
rect 20312 2592 20318 2644
rect 21910 2632 21916 2644
rect 21871 2604 21916 2632
rect 21910 2592 21916 2604
rect 21968 2592 21974 2644
rect 21726 2496 21732 2508
rect 19475 2468 20116 2496
rect 21687 2468 21732 2496
rect 19475 2465 19487 2468
rect 19429 2459 19487 2465
rect 21726 2456 21732 2468
rect 21784 2496 21790 2508
rect 22281 2499 22339 2505
rect 22281 2496 22293 2499
rect 21784 2468 22293 2496
rect 21784 2456 21790 2468
rect 22281 2465 22293 2468
rect 22327 2465 22339 2499
rect 22830 2496 22836 2508
rect 22791 2468 22836 2496
rect 22281 2459 22339 2465
rect 22830 2456 22836 2468
rect 22888 2496 22894 2508
rect 23385 2499 23443 2505
rect 23385 2496 23397 2499
rect 22888 2468 23397 2496
rect 22888 2456 22894 2468
rect 23385 2465 23397 2468
rect 23431 2465 23443 2499
rect 23385 2459 23443 2465
rect 23658 2456 23664 2508
rect 23716 2496 23722 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 23716 2468 24593 2496
rect 23716 2456 23722 2468
rect 24581 2465 24593 2468
rect 24627 2496 24639 2499
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24627 2468 25145 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 18509 2363 18567 2369
rect 18509 2329 18521 2363
rect 18555 2360 18567 2363
rect 19058 2360 19064 2372
rect 18555 2332 19064 2360
rect 18555 2329 18567 2332
rect 18509 2323 18567 2329
rect 19058 2320 19064 2332
rect 19116 2320 19122 2372
rect 19613 2363 19671 2369
rect 19613 2329 19625 2363
rect 19659 2360 19671 2363
rect 21174 2360 21180 2372
rect 19659 2332 21180 2360
rect 19659 2329 19671 2332
rect 19613 2323 19671 2329
rect 21174 2320 21180 2332
rect 21232 2320 21238 2372
rect 23017 2363 23075 2369
rect 23017 2329 23029 2363
rect 23063 2360 23075 2363
rect 25314 2360 25320 2372
rect 23063 2332 25320 2360
rect 23063 2329 23075 2332
rect 23017 2323 23075 2329
rect 25314 2320 25320 2332
rect 25372 2320 25378 2372
rect 11425 2295 11483 2301
rect 11425 2261 11437 2295
rect 11471 2292 11483 2295
rect 11790 2292 11796 2304
rect 11471 2264 11796 2292
rect 11471 2261 11483 2264
rect 11425 2255 11483 2261
rect 11790 2252 11796 2264
rect 11848 2252 11854 2304
rect 17034 2292 17040 2304
rect 16995 2264 17040 2292
rect 17034 2252 17040 2264
rect 17092 2252 17098 2304
rect 24762 2292 24768 2304
rect 24723 2264 24768 2292
rect 24762 2252 24768 2264
rect 24820 2252 24826 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 4068 26256 4120 26308
rect 6184 26256 6236 26308
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 10876 25372 10928 25424
rect 12716 25347 12768 25356
rect 12716 25313 12734 25347
rect 12734 25313 12768 25347
rect 12716 25304 12768 25313
rect 9680 25236 9732 25288
rect 10140 25279 10192 25288
rect 10140 25245 10149 25279
rect 10149 25245 10183 25279
rect 10183 25245 10192 25279
rect 10140 25236 10192 25245
rect 10692 25100 10744 25152
rect 12532 25100 12584 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 12716 24939 12768 24948
rect 12716 24905 12725 24939
rect 12725 24905 12759 24939
rect 12759 24905 12768 24939
rect 12716 24896 12768 24905
rect 5540 24760 5592 24812
rect 8576 24803 8628 24812
rect 8576 24769 8585 24803
rect 8585 24769 8619 24803
rect 8619 24769 8628 24803
rect 8576 24760 8628 24769
rect 10140 24760 10192 24812
rect 15936 24803 15988 24812
rect 15936 24769 15945 24803
rect 15945 24769 15979 24803
rect 15979 24769 15988 24803
rect 15936 24760 15988 24769
rect 9956 24692 10008 24744
rect 13268 24735 13320 24744
rect 13268 24701 13277 24735
rect 13277 24701 13311 24735
rect 13311 24701 13320 24735
rect 13268 24692 13320 24701
rect 9128 24667 9180 24676
rect 9128 24633 9137 24667
rect 9137 24633 9171 24667
rect 9171 24633 9180 24667
rect 9128 24624 9180 24633
rect 9220 24667 9272 24676
rect 9220 24633 9229 24667
rect 9229 24633 9263 24667
rect 9263 24633 9272 24667
rect 9220 24624 9272 24633
rect 10140 24624 10192 24676
rect 10692 24667 10744 24676
rect 10692 24633 10701 24667
rect 10701 24633 10735 24667
rect 10735 24633 10744 24667
rect 10692 24624 10744 24633
rect 5448 24556 5500 24608
rect 6828 24599 6880 24608
rect 6828 24565 6837 24599
rect 6837 24565 6871 24599
rect 6871 24565 6880 24599
rect 6828 24556 6880 24565
rect 7656 24556 7708 24608
rect 10876 24624 10928 24676
rect 11428 24624 11480 24676
rect 13452 24599 13504 24608
rect 13452 24565 13461 24599
rect 13461 24565 13495 24599
rect 13495 24565 13504 24599
rect 13452 24556 13504 24565
rect 16212 24556 16264 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 9128 24395 9180 24404
rect 9128 24361 9137 24395
rect 9137 24361 9171 24395
rect 9171 24361 9180 24395
rect 9128 24352 9180 24361
rect 18236 24395 18288 24404
rect 18236 24361 18245 24395
rect 18245 24361 18279 24395
rect 18279 24361 18288 24395
rect 18236 24352 18288 24361
rect 6552 24327 6604 24336
rect 6552 24293 6561 24327
rect 6561 24293 6595 24327
rect 6595 24293 6604 24327
rect 6552 24284 6604 24293
rect 8116 24327 8168 24336
rect 8116 24293 8125 24327
rect 8125 24293 8159 24327
rect 8159 24293 8168 24327
rect 8116 24284 8168 24293
rect 8484 24284 8536 24336
rect 9220 24284 9272 24336
rect 10968 24284 11020 24336
rect 11428 24327 11480 24336
rect 11428 24293 11437 24327
rect 11437 24293 11471 24327
rect 11471 24293 11480 24327
rect 11428 24284 11480 24293
rect 12992 24327 13044 24336
rect 12992 24293 13001 24327
rect 13001 24293 13035 24327
rect 13035 24293 13044 24327
rect 12992 24284 13044 24293
rect 1492 24259 1544 24268
rect 1492 24225 1510 24259
rect 1510 24225 1544 24259
rect 1492 24216 1544 24225
rect 4620 24216 4672 24268
rect 2688 24080 2740 24132
rect 9956 24216 10008 24268
rect 15384 24259 15436 24268
rect 15384 24225 15402 24259
rect 15402 24225 15436 24259
rect 15384 24216 15436 24225
rect 16304 24259 16356 24268
rect 16304 24225 16313 24259
rect 16313 24225 16347 24259
rect 16347 24225 16356 24259
rect 16304 24216 16356 24225
rect 18420 24216 18472 24268
rect 6460 24191 6512 24200
rect 6460 24157 6469 24191
rect 6469 24157 6503 24191
rect 6503 24157 6512 24191
rect 6460 24148 6512 24157
rect 6736 24191 6788 24200
rect 6736 24157 6745 24191
rect 6745 24157 6779 24191
rect 6779 24157 6788 24191
rect 6736 24148 6788 24157
rect 11520 24148 11572 24200
rect 12716 24148 12768 24200
rect 13544 24191 13596 24200
rect 13544 24157 13553 24191
rect 13553 24157 13587 24191
rect 13587 24157 13596 24191
rect 13544 24148 13596 24157
rect 6644 24080 6696 24132
rect 9864 24080 9916 24132
rect 16488 24123 16540 24132
rect 16488 24089 16497 24123
rect 16497 24089 16531 24123
rect 16531 24089 16540 24123
rect 16488 24080 16540 24089
rect 5264 24055 5316 24064
rect 5264 24021 5273 24055
rect 5273 24021 5307 24055
rect 5307 24021 5316 24055
rect 5264 24012 5316 24021
rect 5540 24012 5592 24064
rect 7564 24055 7616 24064
rect 7564 24021 7573 24055
rect 7573 24021 7607 24055
rect 7607 24021 7616 24055
rect 7564 24012 7616 24021
rect 10692 24012 10744 24064
rect 14096 24055 14148 24064
rect 14096 24021 14105 24055
rect 14105 24021 14139 24055
rect 14139 24021 14148 24055
rect 14096 24012 14148 24021
rect 15292 24012 15344 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1492 23808 1544 23860
rect 4620 23808 4672 23860
rect 6644 23808 6696 23860
rect 8116 23808 8168 23860
rect 9128 23808 9180 23860
rect 9956 23851 10008 23860
rect 9956 23817 9965 23851
rect 9965 23817 9999 23851
rect 9999 23817 10008 23851
rect 11520 23851 11572 23860
rect 9956 23808 10008 23817
rect 6552 23783 6604 23792
rect 6552 23749 6561 23783
rect 6561 23749 6595 23783
rect 6595 23749 6604 23783
rect 6552 23740 6604 23749
rect 8484 23783 8536 23792
rect 8484 23749 8493 23783
rect 8493 23749 8527 23783
rect 8527 23749 8536 23783
rect 8484 23740 8536 23749
rect 5264 23715 5316 23724
rect 5264 23681 5273 23715
rect 5273 23681 5307 23715
rect 5307 23681 5316 23715
rect 5264 23672 5316 23681
rect 7840 23715 7892 23724
rect 7840 23681 7849 23715
rect 7849 23681 7883 23715
rect 7883 23681 7892 23715
rect 7840 23672 7892 23681
rect 11520 23817 11529 23851
rect 11529 23817 11563 23851
rect 11563 23817 11572 23851
rect 11520 23808 11572 23817
rect 12164 23851 12216 23860
rect 12164 23817 12173 23851
rect 12173 23817 12207 23851
rect 12207 23817 12216 23851
rect 12164 23808 12216 23817
rect 15936 23851 15988 23860
rect 15936 23817 15945 23851
rect 15945 23817 15979 23851
rect 15979 23817 15988 23851
rect 15936 23808 15988 23817
rect 16304 23808 16356 23860
rect 16488 23808 16540 23860
rect 17132 23808 17184 23860
rect 19248 23851 19300 23860
rect 19248 23817 19257 23851
rect 19257 23817 19291 23851
rect 19291 23817 19300 23851
rect 19248 23808 19300 23817
rect 21272 23851 21324 23860
rect 21272 23817 21281 23851
rect 21281 23817 21315 23851
rect 21315 23817 21324 23851
rect 21272 23808 21324 23817
rect 22376 23851 22428 23860
rect 22376 23817 22385 23851
rect 22385 23817 22419 23851
rect 22419 23817 22428 23851
rect 22376 23808 22428 23817
rect 11244 23740 11296 23792
rect 12532 23715 12584 23724
rect 12532 23681 12541 23715
rect 12541 23681 12575 23715
rect 12575 23681 12584 23715
rect 12532 23672 12584 23681
rect 13544 23672 13596 23724
rect 14188 23672 14240 23724
rect 17132 23672 17184 23724
rect 480 23604 532 23656
rect 2504 23647 2556 23656
rect 2504 23613 2522 23647
rect 2522 23613 2556 23647
rect 2504 23604 2556 23613
rect 3516 23604 3568 23656
rect 5356 23579 5408 23588
rect 5356 23545 5365 23579
rect 5365 23545 5399 23579
rect 5399 23545 5408 23579
rect 5356 23536 5408 23545
rect 5908 23579 5960 23588
rect 5908 23545 5917 23579
rect 5917 23545 5951 23579
rect 5951 23545 5960 23579
rect 5908 23536 5960 23545
rect 7564 23579 7616 23588
rect 7564 23545 7573 23579
rect 7573 23545 7607 23579
rect 7607 23545 7616 23579
rect 7564 23536 7616 23545
rect 2688 23468 2740 23520
rect 6460 23468 6512 23520
rect 7104 23468 7156 23520
rect 7748 23536 7800 23588
rect 15384 23647 15436 23656
rect 15384 23613 15393 23647
rect 15393 23613 15427 23647
rect 15427 23613 15436 23647
rect 15384 23604 15436 23613
rect 16856 23647 16908 23656
rect 10692 23579 10744 23588
rect 10692 23545 10701 23579
rect 10701 23545 10735 23579
rect 10735 23545 10744 23579
rect 10692 23536 10744 23545
rect 11428 23536 11480 23588
rect 12164 23536 12216 23588
rect 14096 23579 14148 23588
rect 14096 23545 14105 23579
rect 14105 23545 14139 23579
rect 14139 23545 14148 23579
rect 14096 23536 14148 23545
rect 10968 23468 11020 23520
rect 12992 23468 13044 23520
rect 15108 23536 15160 23588
rect 16856 23613 16865 23647
rect 16865 23613 16899 23647
rect 16899 23613 16908 23647
rect 16856 23604 16908 23613
rect 18052 23647 18104 23656
rect 18052 23613 18096 23647
rect 18096 23613 18104 23647
rect 18052 23604 18104 23613
rect 18512 23604 18564 23656
rect 19432 23672 19484 23724
rect 22192 23647 22244 23656
rect 22192 23613 22201 23647
rect 22201 23613 22235 23647
rect 22235 23613 22244 23647
rect 22192 23604 22244 23613
rect 16396 23511 16448 23520
rect 16396 23477 16405 23511
rect 16405 23477 16439 23511
rect 16439 23477 16448 23511
rect 16396 23468 16448 23477
rect 18420 23468 18472 23520
rect 21640 23511 21692 23520
rect 21640 23477 21649 23511
rect 21649 23477 21683 23511
rect 21683 23477 21692 23511
rect 21640 23468 21692 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 5356 23264 5408 23316
rect 5540 23264 5592 23316
rect 6460 23264 6512 23316
rect 10140 23264 10192 23316
rect 12532 23307 12584 23316
rect 12532 23273 12541 23307
rect 12541 23273 12575 23307
rect 12575 23273 12584 23307
rect 12532 23264 12584 23273
rect 12716 23264 12768 23316
rect 16396 23264 16448 23316
rect 6000 23196 6052 23248
rect 7288 23239 7340 23248
rect 7288 23205 7297 23239
rect 7297 23205 7331 23239
rect 7331 23205 7340 23239
rect 7840 23239 7892 23248
rect 7288 23196 7340 23205
rect 7840 23205 7849 23239
rect 7849 23205 7883 23239
rect 7883 23205 7892 23239
rect 7840 23196 7892 23205
rect 11336 23239 11388 23248
rect 11336 23205 11345 23239
rect 11345 23205 11379 23239
rect 11379 23205 11388 23239
rect 11336 23196 11388 23205
rect 13820 23239 13872 23248
rect 13820 23205 13829 23239
rect 13829 23205 13863 23239
rect 13863 23205 13872 23239
rect 13820 23196 13872 23205
rect 10968 23128 11020 23180
rect 15292 23171 15344 23180
rect 15292 23137 15336 23171
rect 15336 23137 15344 23171
rect 15292 23128 15344 23137
rect 16304 23171 16356 23180
rect 16304 23137 16348 23171
rect 16348 23137 16356 23171
rect 16304 23128 16356 23137
rect 17040 23128 17092 23180
rect 5908 23060 5960 23112
rect 6828 23060 6880 23112
rect 6920 23060 6972 23112
rect 11244 23103 11296 23112
rect 11244 23069 11253 23103
rect 11253 23069 11287 23103
rect 11287 23069 11296 23103
rect 11244 23060 11296 23069
rect 11428 23060 11480 23112
rect 12624 23060 12676 23112
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 14188 23103 14240 23112
rect 14188 23069 14197 23103
rect 14197 23069 14231 23103
rect 14231 23069 14240 23103
rect 14188 23060 14240 23069
rect 15384 22924 15436 22976
rect 17868 22924 17920 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 5540 22720 5592 22772
rect 6920 22720 6972 22772
rect 10692 22720 10744 22772
rect 11336 22763 11388 22772
rect 11336 22729 11345 22763
rect 11345 22729 11379 22763
rect 11379 22729 11388 22763
rect 11336 22720 11388 22729
rect 13268 22720 13320 22772
rect 13728 22720 13780 22772
rect 16488 22720 16540 22772
rect 17040 22720 17092 22772
rect 11244 22652 11296 22704
rect 7656 22627 7708 22636
rect 7656 22593 7665 22627
rect 7665 22593 7699 22627
rect 7699 22593 7708 22627
rect 7656 22584 7708 22593
rect 7840 22584 7892 22636
rect 14188 22584 14240 22636
rect 15292 22627 15344 22636
rect 15292 22593 15301 22627
rect 15301 22593 15335 22627
rect 15335 22593 15344 22627
rect 15292 22584 15344 22593
rect 17224 22584 17276 22636
rect 6552 22448 6604 22500
rect 7472 22448 7524 22500
rect 10968 22559 11020 22568
rect 10968 22525 10977 22559
rect 10977 22525 11011 22559
rect 11011 22525 11020 22559
rect 10968 22516 11020 22525
rect 12624 22516 12676 22568
rect 9956 22448 10008 22500
rect 14004 22491 14056 22500
rect 14004 22457 14013 22491
rect 14013 22457 14047 22491
rect 14047 22457 14056 22491
rect 14004 22448 14056 22457
rect 14740 22448 14792 22500
rect 16304 22448 16356 22500
rect 6000 22380 6052 22432
rect 7288 22380 7340 22432
rect 9128 22423 9180 22432
rect 9128 22389 9137 22423
rect 9137 22389 9171 22423
rect 9171 22389 9180 22423
rect 9128 22380 9180 22389
rect 13820 22380 13872 22432
rect 14648 22380 14700 22432
rect 15384 22380 15436 22432
rect 17132 22380 17184 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5080 22219 5132 22228
rect 5080 22185 5089 22219
rect 5089 22185 5123 22219
rect 5123 22185 5132 22219
rect 5080 22176 5132 22185
rect 7472 22176 7524 22228
rect 7840 22176 7892 22228
rect 6184 22108 6236 22160
rect 7656 22108 7708 22160
rect 11336 22176 11388 22228
rect 5080 22083 5132 22092
rect 5080 22049 5089 22083
rect 5089 22049 5123 22083
rect 5123 22049 5132 22083
rect 5080 22040 5132 22049
rect 5448 22040 5500 22092
rect 8116 22083 8168 22092
rect 8116 22049 8160 22083
rect 8160 22049 8168 22083
rect 9956 22108 10008 22160
rect 8116 22040 8168 22049
rect 8668 22040 8720 22092
rect 12256 22040 12308 22092
rect 14004 22176 14056 22228
rect 14188 22219 14240 22228
rect 14188 22185 14197 22219
rect 14197 22185 14231 22219
rect 14231 22185 14240 22219
rect 14188 22176 14240 22185
rect 15568 22083 15620 22092
rect 6368 22015 6420 22024
rect 6368 21981 6377 22015
rect 6377 21981 6411 22015
rect 6411 21981 6420 22015
rect 6368 21972 6420 21981
rect 7564 21972 7616 22024
rect 10140 21972 10192 22024
rect 11888 21972 11940 22024
rect 15568 22049 15577 22083
rect 15577 22049 15611 22083
rect 15611 22049 15620 22083
rect 15568 22040 15620 22049
rect 15752 22083 15804 22092
rect 15752 22049 15761 22083
rect 15761 22049 15795 22083
rect 15795 22049 15804 22083
rect 15752 22040 15804 22049
rect 17224 22108 17276 22160
rect 17040 21947 17092 21956
rect 17040 21913 17049 21947
rect 17049 21913 17083 21947
rect 17083 21913 17092 21947
rect 17040 21904 17092 21913
rect 6000 21836 6052 21888
rect 7288 21879 7340 21888
rect 7288 21845 7297 21879
rect 7297 21845 7331 21879
rect 7331 21845 7340 21879
rect 7288 21836 7340 21845
rect 14280 21836 14332 21888
rect 14648 21836 14700 21888
rect 16304 21879 16356 21888
rect 16304 21845 16313 21879
rect 16313 21845 16347 21879
rect 16347 21845 16356 21879
rect 16304 21836 16356 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 6184 21675 6236 21684
rect 6184 21641 6193 21675
rect 6193 21641 6227 21675
rect 6227 21641 6236 21675
rect 6184 21632 6236 21641
rect 11888 21675 11940 21684
rect 11888 21641 11897 21675
rect 11897 21641 11931 21675
rect 11931 21641 11940 21675
rect 11888 21632 11940 21641
rect 13728 21675 13780 21684
rect 13728 21641 13737 21675
rect 13737 21641 13771 21675
rect 13771 21641 13780 21675
rect 13728 21632 13780 21641
rect 6000 21496 6052 21548
rect 6552 21496 6604 21548
rect 8668 21539 8720 21548
rect 5632 21471 5684 21480
rect 5632 21437 5641 21471
rect 5641 21437 5675 21471
rect 5675 21437 5684 21471
rect 5632 21428 5684 21437
rect 7012 21428 7064 21480
rect 8668 21505 8677 21539
rect 8677 21505 8711 21539
rect 8711 21505 8720 21539
rect 8668 21496 8720 21505
rect 9312 21539 9364 21548
rect 9312 21505 9321 21539
rect 9321 21505 9355 21539
rect 9355 21505 9364 21539
rect 9312 21496 9364 21505
rect 14280 21564 14332 21616
rect 16028 21564 16080 21616
rect 14740 21539 14792 21548
rect 14740 21505 14749 21539
rect 14749 21505 14783 21539
rect 14783 21505 14792 21539
rect 14740 21496 14792 21505
rect 10692 21428 10744 21480
rect 4528 21335 4580 21344
rect 4528 21301 4537 21335
rect 4537 21301 4571 21335
rect 4571 21301 4580 21335
rect 4528 21292 4580 21301
rect 5080 21292 5132 21344
rect 6184 21292 6236 21344
rect 8668 21360 8720 21412
rect 11336 21360 11388 21412
rect 12440 21360 12492 21412
rect 12992 21360 13044 21412
rect 14280 21403 14332 21412
rect 14280 21369 14289 21403
rect 14289 21369 14323 21403
rect 14323 21369 14332 21403
rect 14280 21360 14332 21369
rect 15844 21403 15896 21412
rect 8208 21335 8260 21344
rect 8208 21301 8217 21335
rect 8217 21301 8251 21335
rect 8251 21301 8260 21335
rect 8208 21292 8260 21301
rect 9956 21292 10008 21344
rect 12256 21335 12308 21344
rect 12256 21301 12265 21335
rect 12265 21301 12299 21335
rect 12299 21301 12308 21335
rect 12256 21292 12308 21301
rect 14004 21335 14056 21344
rect 14004 21301 14013 21335
rect 14013 21301 14047 21335
rect 14047 21301 14056 21335
rect 15844 21369 15853 21403
rect 15853 21369 15887 21403
rect 15887 21369 15896 21403
rect 15844 21360 15896 21369
rect 16304 21360 16356 21412
rect 15292 21335 15344 21344
rect 14004 21292 14056 21301
rect 15292 21301 15301 21335
rect 15301 21301 15335 21335
rect 15335 21301 15344 21335
rect 15292 21292 15344 21301
rect 15568 21292 15620 21344
rect 17224 21292 17276 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 7012 21131 7064 21140
rect 7012 21097 7021 21131
rect 7021 21097 7055 21131
rect 7055 21097 7064 21131
rect 7012 21088 7064 21097
rect 8668 21131 8720 21140
rect 8668 21097 8677 21131
rect 8677 21097 8711 21131
rect 8711 21097 8720 21131
rect 8668 21088 8720 21097
rect 11060 21088 11112 21140
rect 6368 21063 6420 21072
rect 6368 21029 6377 21063
rect 6377 21029 6411 21063
rect 6411 21029 6420 21063
rect 6368 21020 6420 21029
rect 7288 21020 7340 21072
rect 8208 21020 8260 21072
rect 9312 21020 9364 21072
rect 12992 21088 13044 21140
rect 14004 21088 14056 21140
rect 15016 21131 15068 21140
rect 15016 21097 15025 21131
rect 15025 21097 15059 21131
rect 15059 21097 15068 21131
rect 15016 21088 15068 21097
rect 15844 21088 15896 21140
rect 12256 21020 12308 21072
rect 15384 21063 15436 21072
rect 15384 21029 15393 21063
rect 15393 21029 15427 21063
rect 15427 21029 15436 21063
rect 15384 21020 15436 21029
rect 15476 21063 15528 21072
rect 15476 21029 15485 21063
rect 15485 21029 15519 21063
rect 15519 21029 15528 21063
rect 16028 21063 16080 21072
rect 15476 21020 15528 21029
rect 16028 21029 16037 21063
rect 16037 21029 16071 21063
rect 16071 21029 16080 21063
rect 16028 21020 16080 21029
rect 5632 20995 5684 21004
rect 5632 20961 5641 20995
rect 5641 20961 5675 20995
rect 5675 20961 5684 20995
rect 5632 20952 5684 20961
rect 6184 20995 6236 21004
rect 6184 20961 6193 20995
rect 6193 20961 6227 20995
rect 6227 20961 6236 20995
rect 6184 20952 6236 20961
rect 10416 20952 10468 21004
rect 6920 20884 6972 20936
rect 9864 20884 9916 20936
rect 10692 20884 10744 20936
rect 11152 20927 11204 20936
rect 11152 20893 11161 20927
rect 11161 20893 11195 20927
rect 11195 20893 11204 20927
rect 11152 20884 11204 20893
rect 11612 20927 11664 20936
rect 11612 20893 11621 20927
rect 11621 20893 11655 20927
rect 11655 20893 11664 20927
rect 11612 20884 11664 20893
rect 12808 20927 12860 20936
rect 12808 20893 12817 20927
rect 12817 20893 12851 20927
rect 12851 20893 12860 20927
rect 12808 20884 12860 20893
rect 13728 20884 13780 20936
rect 9680 20816 9732 20868
rect 10140 20816 10192 20868
rect 4528 20748 4580 20800
rect 5448 20748 5500 20800
rect 9772 20748 9824 20800
rect 14464 20791 14516 20800
rect 14464 20757 14473 20791
rect 14473 20757 14507 20791
rect 14507 20757 14516 20791
rect 14464 20748 14516 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 6184 20587 6236 20596
rect 6184 20553 6193 20587
rect 6193 20553 6227 20587
rect 6227 20553 6236 20587
rect 6184 20544 6236 20553
rect 6828 20544 6880 20596
rect 7288 20587 7340 20596
rect 7288 20553 7297 20587
rect 7297 20553 7331 20587
rect 7331 20553 7340 20587
rect 7288 20544 7340 20553
rect 11060 20587 11112 20596
rect 11060 20553 11069 20587
rect 11069 20553 11103 20587
rect 11103 20553 11112 20587
rect 11060 20544 11112 20553
rect 13728 20544 13780 20596
rect 15384 20544 15436 20596
rect 8208 20519 8260 20528
rect 8208 20485 8217 20519
rect 8217 20485 8251 20519
rect 8251 20485 8260 20519
rect 8208 20476 8260 20485
rect 9956 20476 10008 20528
rect 12256 20476 12308 20528
rect 15476 20519 15528 20528
rect 15476 20485 15485 20519
rect 15485 20485 15519 20519
rect 15519 20485 15528 20519
rect 15476 20476 15528 20485
rect 9128 20451 9180 20460
rect 9128 20417 9137 20451
rect 9137 20417 9171 20451
rect 9171 20417 9180 20451
rect 9128 20408 9180 20417
rect 11152 20408 11204 20460
rect 14096 20408 14148 20460
rect 14740 20451 14792 20460
rect 14740 20417 14749 20451
rect 14749 20417 14783 20451
rect 14783 20417 14792 20451
rect 14740 20408 14792 20417
rect 15844 20408 15896 20460
rect 5356 20383 5408 20392
rect 5356 20349 5365 20383
rect 5365 20349 5399 20383
rect 5399 20349 5408 20383
rect 5356 20340 5408 20349
rect 5448 20340 5500 20392
rect 5724 20383 5776 20392
rect 5724 20349 5733 20383
rect 5733 20349 5767 20383
rect 5767 20349 5776 20383
rect 5724 20340 5776 20349
rect 10416 20383 10468 20392
rect 10416 20349 10425 20383
rect 10425 20349 10459 20383
rect 10459 20349 10468 20383
rect 10416 20340 10468 20349
rect 7748 20315 7800 20324
rect 7748 20281 7757 20315
rect 7757 20281 7791 20315
rect 7791 20281 7800 20315
rect 7748 20272 7800 20281
rect 8576 20247 8628 20256
rect 8576 20213 8585 20247
rect 8585 20213 8619 20247
rect 8619 20213 8628 20247
rect 8576 20204 8628 20213
rect 8760 20204 8812 20256
rect 9956 20272 10008 20324
rect 12256 20340 12308 20392
rect 12440 20340 12492 20392
rect 13268 20340 13320 20392
rect 13820 20340 13872 20392
rect 14464 20315 14516 20324
rect 14464 20281 14473 20315
rect 14473 20281 14507 20315
rect 14507 20281 14516 20315
rect 14464 20272 14516 20281
rect 11980 20204 12032 20256
rect 14188 20247 14240 20256
rect 14188 20213 14197 20247
rect 14197 20213 14231 20247
rect 14231 20213 14240 20247
rect 14188 20204 14240 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 5540 20000 5592 20052
rect 7196 20000 7248 20052
rect 7748 20000 7800 20052
rect 9128 20043 9180 20052
rect 9128 20009 9137 20043
rect 9137 20009 9171 20043
rect 9171 20009 9180 20043
rect 9128 20000 9180 20009
rect 11888 20000 11940 20052
rect 13268 20043 13320 20052
rect 6552 19975 6604 19984
rect 6552 19941 6555 19975
rect 6555 19941 6589 19975
rect 6589 19941 6604 19975
rect 6552 19932 6604 19941
rect 8024 19932 8076 19984
rect 9956 19932 10008 19984
rect 13268 20009 13277 20043
rect 13277 20009 13311 20043
rect 13311 20009 13320 20043
rect 13268 20000 13320 20009
rect 12624 19975 12676 19984
rect 12624 19941 12633 19975
rect 12633 19941 12667 19975
rect 12667 19941 12676 19975
rect 12624 19932 12676 19941
rect 13820 19975 13872 19984
rect 13820 19941 13829 19975
rect 13829 19941 13863 19975
rect 13863 19941 13872 19975
rect 13820 19932 13872 19941
rect 14096 19932 14148 19984
rect 5080 19864 5132 19916
rect 16028 19864 16080 19916
rect 8300 19796 8352 19848
rect 8208 19728 8260 19780
rect 8576 19771 8628 19780
rect 8576 19737 8585 19771
rect 8585 19737 8619 19771
rect 8619 19737 8628 19771
rect 8576 19728 8628 19737
rect 6000 19703 6052 19712
rect 6000 19669 6009 19703
rect 6009 19669 6043 19703
rect 6043 19669 6052 19703
rect 6000 19660 6052 19669
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 11612 19660 11664 19712
rect 12256 19796 12308 19848
rect 12992 19796 13044 19848
rect 14372 19839 14424 19848
rect 14372 19805 14381 19839
rect 14381 19805 14415 19839
rect 14415 19805 14424 19839
rect 14372 19796 14424 19805
rect 13912 19728 13964 19780
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 6552 19499 6604 19508
rect 6552 19465 6561 19499
rect 6561 19465 6595 19499
rect 6595 19465 6604 19499
rect 6552 19456 6604 19465
rect 7748 19499 7800 19508
rect 7748 19465 7757 19499
rect 7757 19465 7791 19499
rect 7791 19465 7800 19499
rect 7748 19456 7800 19465
rect 8024 19499 8076 19508
rect 8024 19465 8033 19499
rect 8033 19465 8067 19499
rect 8067 19465 8076 19499
rect 8024 19456 8076 19465
rect 11888 19499 11940 19508
rect 11888 19465 11897 19499
rect 11897 19465 11931 19499
rect 11931 19465 11940 19499
rect 11888 19456 11940 19465
rect 12992 19499 13044 19508
rect 12992 19465 13001 19499
rect 13001 19465 13035 19499
rect 13035 19465 13044 19499
rect 12992 19456 13044 19465
rect 14188 19456 14240 19508
rect 13820 19388 13872 19440
rect 16028 19431 16080 19440
rect 16028 19397 16037 19431
rect 16037 19397 16071 19431
rect 16071 19397 16080 19431
rect 16028 19388 16080 19397
rect 6000 19320 6052 19372
rect 9588 19363 9640 19372
rect 9588 19329 9597 19363
rect 9597 19329 9631 19363
rect 9631 19329 9640 19363
rect 9588 19320 9640 19329
rect 5540 19252 5592 19304
rect 5724 19295 5776 19304
rect 5724 19261 5733 19295
rect 5733 19261 5767 19295
rect 5767 19261 5776 19295
rect 5724 19252 5776 19261
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 8300 19252 8352 19304
rect 9036 19295 9088 19304
rect 9036 19261 9045 19295
rect 9045 19261 9079 19295
rect 9079 19261 9088 19295
rect 9036 19252 9088 19261
rect 10692 19295 10744 19304
rect 5356 19184 5408 19236
rect 6552 19184 6604 19236
rect 10692 19261 10701 19295
rect 10701 19261 10735 19295
rect 10735 19261 10744 19295
rect 10692 19252 10744 19261
rect 11060 19295 11112 19304
rect 11060 19261 11069 19295
rect 11069 19261 11103 19295
rect 11103 19261 11112 19295
rect 11060 19252 11112 19261
rect 11336 19252 11388 19304
rect 13084 19252 13136 19304
rect 21364 19320 21416 19372
rect 21640 19320 21692 19372
rect 14924 19295 14976 19304
rect 12440 19184 12492 19236
rect 12992 19184 13044 19236
rect 14924 19261 14933 19295
rect 14933 19261 14967 19295
rect 14967 19261 14976 19295
rect 14924 19252 14976 19261
rect 5080 19159 5132 19168
rect 5080 19125 5089 19159
rect 5089 19125 5123 19159
rect 5123 19125 5132 19159
rect 5080 19116 5132 19125
rect 8852 19159 8904 19168
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 8852 19116 8904 19125
rect 10140 19159 10192 19168
rect 10140 19125 10149 19159
rect 10149 19125 10183 19159
rect 10183 19125 10192 19159
rect 10140 19116 10192 19125
rect 15200 19159 15252 19168
rect 15200 19125 15209 19159
rect 15209 19125 15243 19159
rect 15243 19125 15252 19159
rect 15200 19116 15252 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 7472 18912 7524 18964
rect 6828 18844 6880 18896
rect 9680 18912 9732 18964
rect 10692 18955 10744 18964
rect 10692 18921 10701 18955
rect 10701 18921 10735 18955
rect 10735 18921 10744 18955
rect 10692 18912 10744 18921
rect 11060 18912 11112 18964
rect 10968 18844 11020 18896
rect 11152 18844 11204 18896
rect 12164 18844 12216 18896
rect 12440 18955 12492 18964
rect 12440 18921 12449 18955
rect 12449 18921 12483 18955
rect 12483 18921 12492 18955
rect 13084 18955 13136 18964
rect 12440 18912 12492 18921
rect 13084 18921 13093 18955
rect 13093 18921 13127 18955
rect 13127 18921 13136 18955
rect 13084 18912 13136 18921
rect 13912 18955 13964 18964
rect 13912 18921 13921 18955
rect 13921 18921 13955 18955
rect 13955 18921 13964 18955
rect 13912 18912 13964 18921
rect 14924 18955 14976 18964
rect 14924 18921 14933 18955
rect 14933 18921 14967 18955
rect 14967 18921 14976 18955
rect 14924 18912 14976 18921
rect 5540 18776 5592 18828
rect 6460 18819 6512 18828
rect 6460 18785 6469 18819
rect 6469 18785 6503 18819
rect 6503 18785 6512 18819
rect 6460 18776 6512 18785
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 8208 18751 8260 18760
rect 8208 18717 8217 18751
rect 8217 18717 8251 18751
rect 8251 18717 8260 18751
rect 8208 18708 8260 18717
rect 9036 18751 9088 18760
rect 9036 18717 9045 18751
rect 9045 18717 9079 18751
rect 9079 18717 9088 18751
rect 10692 18776 10744 18828
rect 11060 18776 11112 18828
rect 13360 18819 13412 18828
rect 9036 18708 9088 18717
rect 10968 18708 11020 18760
rect 11336 18751 11388 18760
rect 11336 18717 11345 18751
rect 11345 18717 11379 18751
rect 11379 18717 11388 18751
rect 11336 18708 11388 18717
rect 11612 18751 11664 18760
rect 11612 18717 11621 18751
rect 11621 18717 11655 18751
rect 11655 18717 11664 18751
rect 11612 18708 11664 18717
rect 13360 18785 13369 18819
rect 13369 18785 13403 18819
rect 13403 18785 13412 18819
rect 13360 18776 13412 18785
rect 15384 18819 15436 18828
rect 15384 18785 15402 18819
rect 15402 18785 15436 18819
rect 15384 18776 15436 18785
rect 13176 18708 13228 18760
rect 14924 18708 14976 18760
rect 5724 18640 5776 18692
rect 6368 18572 6420 18624
rect 6920 18615 6972 18624
rect 6920 18581 6929 18615
rect 6929 18581 6963 18615
rect 6963 18581 6972 18615
rect 6920 18572 6972 18581
rect 14280 18615 14332 18624
rect 14280 18581 14289 18615
rect 14289 18581 14323 18615
rect 14323 18581 14332 18615
rect 14280 18572 14332 18581
rect 15936 18572 15988 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 5172 18368 5224 18420
rect 5540 18368 5592 18420
rect 6552 18411 6604 18420
rect 6552 18377 6561 18411
rect 6561 18377 6595 18411
rect 6595 18377 6604 18411
rect 6552 18368 6604 18377
rect 7472 18368 7524 18420
rect 11152 18411 11204 18420
rect 11152 18377 11161 18411
rect 11161 18377 11195 18411
rect 11195 18377 11204 18411
rect 11152 18368 11204 18377
rect 11336 18368 11388 18420
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 13360 18368 13412 18420
rect 15384 18411 15436 18420
rect 15384 18377 15393 18411
rect 15393 18377 15427 18411
rect 15427 18377 15436 18411
rect 15384 18368 15436 18377
rect 6460 18232 6512 18284
rect 12440 18275 12492 18284
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 14372 18232 14424 18284
rect 5540 18164 5592 18216
rect 6920 18164 6972 18216
rect 9220 18164 9272 18216
rect 10692 18164 10744 18216
rect 11888 18164 11940 18216
rect 6552 18096 6604 18148
rect 7840 18096 7892 18148
rect 8760 18096 8812 18148
rect 10140 18096 10192 18148
rect 13268 18164 13320 18216
rect 10968 18028 11020 18080
rect 12164 18071 12216 18080
rect 12164 18037 12173 18071
rect 12173 18037 12207 18071
rect 12207 18037 12216 18071
rect 12164 18028 12216 18037
rect 16580 18207 16632 18216
rect 16580 18173 16589 18207
rect 16589 18173 16623 18207
rect 16623 18173 16632 18207
rect 16580 18164 16632 18173
rect 13820 18096 13872 18148
rect 14280 18139 14332 18148
rect 14280 18105 14289 18139
rect 14289 18105 14323 18139
rect 14323 18105 14332 18139
rect 14280 18096 14332 18105
rect 16764 18028 16816 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 7104 17824 7156 17876
rect 7564 17824 7616 17876
rect 10876 17824 10928 17876
rect 11336 17867 11388 17876
rect 11336 17833 11345 17867
rect 11345 17833 11379 17867
rect 11379 17833 11388 17867
rect 11336 17824 11388 17833
rect 13176 17867 13228 17876
rect 6552 17756 6604 17808
rect 10140 17756 10192 17808
rect 12164 17756 12216 17808
rect 13176 17833 13185 17867
rect 13185 17833 13219 17867
rect 13219 17833 13228 17867
rect 13176 17824 13228 17833
rect 13452 17756 13504 17808
rect 15476 17824 15528 17876
rect 16212 17867 16264 17876
rect 16212 17833 16221 17867
rect 16221 17833 16255 17867
rect 16255 17833 16264 17867
rect 16212 17824 16264 17833
rect 14372 17799 14424 17808
rect 14372 17765 14381 17799
rect 14381 17765 14415 17799
rect 14415 17765 14424 17799
rect 14372 17756 14424 17765
rect 16580 17756 16632 17808
rect 5172 17731 5224 17740
rect 5172 17697 5181 17731
rect 5181 17697 5215 17731
rect 5215 17697 5224 17731
rect 5172 17688 5224 17697
rect 5356 17731 5408 17740
rect 5356 17697 5365 17731
rect 5365 17697 5399 17731
rect 5399 17697 5408 17731
rect 5356 17688 5408 17697
rect 8668 17688 8720 17740
rect 15384 17731 15436 17740
rect 15384 17697 15402 17731
rect 15402 17697 15436 17731
rect 15384 17688 15436 17697
rect 5448 17663 5500 17672
rect 5448 17629 5457 17663
rect 5457 17629 5491 17663
rect 5491 17629 5500 17663
rect 5448 17620 5500 17629
rect 6460 17663 6512 17672
rect 6460 17629 6469 17663
rect 6469 17629 6503 17663
rect 6503 17629 6512 17663
rect 6460 17620 6512 17629
rect 9680 17663 9732 17672
rect 9680 17629 9689 17663
rect 9689 17629 9723 17663
rect 9723 17629 9732 17663
rect 9680 17620 9732 17629
rect 11796 17620 11848 17672
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 15752 17620 15804 17672
rect 16672 17620 16724 17672
rect 16948 17552 17000 17604
rect 9220 17527 9272 17536
rect 9220 17493 9229 17527
rect 9229 17493 9263 17527
rect 9263 17493 9272 17527
rect 9220 17484 9272 17493
rect 10968 17527 11020 17536
rect 10968 17493 10977 17527
rect 10977 17493 11011 17527
rect 11011 17493 11020 17527
rect 10968 17484 11020 17493
rect 16120 17484 16172 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 5172 17280 5224 17332
rect 6276 17323 6328 17332
rect 6276 17289 6285 17323
rect 6285 17289 6319 17323
rect 6319 17289 6328 17323
rect 6276 17280 6328 17289
rect 6644 17323 6696 17332
rect 6644 17289 6653 17323
rect 6653 17289 6687 17323
rect 6687 17289 6696 17323
rect 6644 17280 6696 17289
rect 7104 17280 7156 17332
rect 7748 17280 7800 17332
rect 10140 17323 10192 17332
rect 10140 17289 10149 17323
rect 10149 17289 10183 17323
rect 10183 17289 10192 17323
rect 10140 17280 10192 17289
rect 10876 17280 10928 17332
rect 5356 17212 5408 17264
rect 8208 17255 8260 17264
rect 8208 17221 8217 17255
rect 8217 17221 8251 17255
rect 8251 17221 8260 17255
rect 8208 17212 8260 17221
rect 8668 17255 8720 17264
rect 8668 17221 8677 17255
rect 8677 17221 8711 17255
rect 8711 17221 8720 17255
rect 8668 17212 8720 17221
rect 12164 17280 12216 17332
rect 13452 17323 13504 17332
rect 13452 17289 13461 17323
rect 13461 17289 13495 17323
rect 13495 17289 13504 17323
rect 13452 17280 13504 17289
rect 13820 17280 13872 17332
rect 14648 17280 14700 17332
rect 15384 17323 15436 17332
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 11612 17212 11664 17264
rect 16212 17212 16264 17264
rect 10968 17144 11020 17196
rect 6736 17076 6788 17128
rect 9496 17076 9548 17128
rect 9588 17119 9640 17128
rect 9588 17085 9597 17119
rect 9597 17085 9631 17119
rect 9631 17085 9640 17119
rect 9588 17076 9640 17085
rect 13636 17119 13688 17128
rect 6460 17008 6512 17060
rect 7656 17051 7708 17060
rect 7656 17017 7665 17051
rect 7665 17017 7699 17051
rect 7699 17017 7708 17051
rect 7656 17008 7708 17017
rect 7748 17051 7800 17060
rect 7748 17017 7757 17051
rect 7757 17017 7791 17051
rect 7791 17017 7800 17051
rect 7748 17008 7800 17017
rect 10876 17008 10928 17060
rect 13636 17085 13638 17119
rect 13638 17085 13688 17119
rect 14096 17119 14148 17128
rect 13636 17076 13688 17085
rect 14096 17085 14105 17119
rect 14105 17085 14139 17119
rect 14139 17085 14148 17119
rect 14096 17076 14148 17085
rect 14648 17119 14700 17128
rect 14648 17085 14666 17119
rect 14666 17085 14700 17119
rect 14648 17076 14700 17085
rect 17040 17076 17092 17128
rect 16764 17008 16816 17060
rect 16948 17051 17000 17060
rect 16948 17017 16957 17051
rect 16957 17017 16991 17051
rect 16991 17017 17000 17051
rect 16948 17008 17000 17017
rect 18052 17051 18104 17060
rect 18052 17017 18061 17051
rect 18061 17017 18095 17051
rect 18095 17017 18104 17051
rect 18052 17008 18104 17017
rect 9220 16983 9272 16992
rect 9220 16949 9229 16983
rect 9229 16949 9263 16983
rect 9263 16949 9272 16983
rect 9220 16940 9272 16949
rect 12992 16983 13044 16992
rect 12992 16949 13001 16983
rect 13001 16949 13035 16983
rect 13035 16949 13044 16983
rect 12992 16940 13044 16949
rect 14464 16940 14516 16992
rect 15752 16983 15804 16992
rect 15752 16949 15761 16983
rect 15761 16949 15795 16983
rect 15795 16949 15804 16983
rect 15752 16940 15804 16949
rect 16488 16940 16540 16992
rect 18328 16940 18380 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 4344 16779 4396 16788
rect 4344 16745 4353 16779
rect 4353 16745 4387 16779
rect 4387 16745 4396 16779
rect 4344 16736 4396 16745
rect 5172 16736 5224 16788
rect 6184 16736 6236 16788
rect 6460 16779 6512 16788
rect 6460 16745 6469 16779
rect 6469 16745 6503 16779
rect 6503 16745 6512 16779
rect 6460 16736 6512 16745
rect 7656 16668 7708 16720
rect 4252 16600 4304 16652
rect 5172 16643 5224 16652
rect 5172 16609 5216 16643
rect 5216 16609 5224 16643
rect 6184 16643 6236 16652
rect 5172 16600 5224 16609
rect 6184 16609 6193 16643
rect 6193 16609 6227 16643
rect 6227 16609 6236 16643
rect 6184 16600 6236 16609
rect 7932 16600 7984 16652
rect 8484 16600 8536 16652
rect 8852 16736 8904 16788
rect 9588 16736 9640 16788
rect 11152 16736 11204 16788
rect 13728 16736 13780 16788
rect 9680 16668 9732 16720
rect 11796 16668 11848 16720
rect 11980 16711 12032 16720
rect 11980 16677 11989 16711
rect 11989 16677 12023 16711
rect 12023 16677 12032 16711
rect 11980 16668 12032 16677
rect 12348 16668 12400 16720
rect 15200 16668 15252 16720
rect 16672 16711 16724 16720
rect 16672 16677 16681 16711
rect 16681 16677 16715 16711
rect 16715 16677 16724 16711
rect 16672 16668 16724 16677
rect 16764 16711 16816 16720
rect 16764 16677 16773 16711
rect 16773 16677 16807 16711
rect 16807 16677 16816 16711
rect 16764 16668 16816 16677
rect 17316 16668 17368 16720
rect 18788 16736 18840 16788
rect 18328 16711 18380 16720
rect 18328 16677 18337 16711
rect 18337 16677 18371 16711
rect 18371 16677 18380 16711
rect 18328 16668 18380 16677
rect 10140 16600 10192 16652
rect 10692 16600 10744 16652
rect 13452 16643 13504 16652
rect 13452 16609 13496 16643
rect 13496 16609 13504 16643
rect 13452 16600 13504 16609
rect 15292 16643 15344 16652
rect 15292 16609 15336 16643
rect 15336 16609 15344 16643
rect 15292 16600 15344 16609
rect 19432 16600 19484 16652
rect 11336 16532 11388 16584
rect 10784 16464 10836 16516
rect 13728 16464 13780 16516
rect 18144 16464 18196 16516
rect 12624 16396 12676 16448
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 15660 16396 15712 16448
rect 16212 16439 16264 16448
rect 16212 16405 16221 16439
rect 16221 16405 16255 16439
rect 16255 16405 16264 16439
rect 16212 16396 16264 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 6184 16192 6236 16244
rect 8484 16235 8536 16244
rect 8484 16201 8493 16235
rect 8493 16201 8527 16235
rect 8527 16201 8536 16235
rect 8484 16192 8536 16201
rect 10232 16192 10284 16244
rect 7932 16124 7984 16176
rect 10140 16124 10192 16176
rect 13360 16192 13412 16244
rect 15568 16235 15620 16244
rect 15568 16201 15577 16235
rect 15577 16201 15611 16235
rect 15611 16201 15620 16235
rect 15568 16192 15620 16201
rect 17040 16235 17092 16244
rect 17040 16201 17049 16235
rect 17049 16201 17083 16235
rect 17083 16201 17092 16235
rect 17040 16192 17092 16201
rect 17316 16235 17368 16244
rect 17316 16201 17325 16235
rect 17325 16201 17359 16235
rect 17359 16201 17368 16235
rect 17316 16192 17368 16201
rect 18052 16192 18104 16244
rect 5264 16031 5316 16040
rect 5264 15997 5273 16031
rect 5273 15997 5307 16031
rect 5307 15997 5316 16031
rect 5264 15988 5316 15997
rect 7564 16031 7616 16040
rect 4252 15895 4304 15904
rect 4252 15861 4261 15895
rect 4261 15861 4295 15895
rect 4295 15861 4304 15895
rect 4252 15852 4304 15861
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 5632 15852 5684 15861
rect 7564 15997 7573 16031
rect 7573 15997 7607 16031
rect 7607 15997 7616 16031
rect 7564 15988 7616 15997
rect 7748 15963 7800 15972
rect 7748 15929 7757 15963
rect 7757 15929 7791 15963
rect 7791 15929 7800 15963
rect 7748 15920 7800 15929
rect 8760 15988 8812 16040
rect 9036 15988 9088 16040
rect 14188 16124 14240 16176
rect 15292 16124 15344 16176
rect 9680 15963 9732 15972
rect 9680 15929 9689 15963
rect 9689 15929 9723 15963
rect 9723 15929 9732 15963
rect 9680 15920 9732 15929
rect 10140 15920 10192 15972
rect 13912 15988 13964 16040
rect 18144 16099 18196 16108
rect 18144 16065 18153 16099
rect 18153 16065 18187 16099
rect 18187 16065 18196 16099
rect 18144 16056 18196 16065
rect 15568 15988 15620 16040
rect 15660 15988 15712 16040
rect 12624 15963 12676 15972
rect 12624 15929 12633 15963
rect 12633 15929 12667 15963
rect 12667 15929 12676 15963
rect 13176 15963 13228 15972
rect 12624 15920 12676 15929
rect 13176 15929 13185 15963
rect 13185 15929 13219 15963
rect 13219 15929 13228 15963
rect 13176 15920 13228 15929
rect 16212 15920 16264 15972
rect 18144 15920 18196 15972
rect 18880 15920 18932 15972
rect 19156 15920 19208 15972
rect 7932 15852 7984 15904
rect 8760 15895 8812 15904
rect 8760 15861 8769 15895
rect 8769 15861 8803 15895
rect 8803 15861 8812 15895
rect 8760 15852 8812 15861
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 12348 15852 12400 15904
rect 13452 15895 13504 15904
rect 13452 15861 13461 15895
rect 13461 15861 13495 15895
rect 13495 15861 13504 15895
rect 13452 15852 13504 15861
rect 13544 15852 13596 15904
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 19064 15852 19116 15861
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 5632 15648 5684 15700
rect 7104 15691 7156 15700
rect 7104 15657 7113 15691
rect 7113 15657 7147 15691
rect 7147 15657 7156 15691
rect 7104 15648 7156 15657
rect 7564 15648 7616 15700
rect 9036 15691 9088 15700
rect 9036 15657 9045 15691
rect 9045 15657 9079 15691
rect 9079 15657 9088 15691
rect 9036 15648 9088 15657
rect 9680 15648 9732 15700
rect 10692 15648 10744 15700
rect 11980 15648 12032 15700
rect 13544 15648 13596 15700
rect 16488 15691 16540 15700
rect 16488 15657 16497 15691
rect 16497 15657 16531 15691
rect 16531 15657 16540 15691
rect 16488 15648 16540 15657
rect 16672 15648 16724 15700
rect 17960 15648 18012 15700
rect 18328 15691 18380 15700
rect 18328 15657 18337 15691
rect 18337 15657 18371 15691
rect 18371 15657 18380 15691
rect 18328 15648 18380 15657
rect 18788 15691 18840 15700
rect 18788 15657 18797 15691
rect 18797 15657 18831 15691
rect 18831 15657 18840 15691
rect 18788 15648 18840 15657
rect 7840 15623 7892 15632
rect 7840 15589 7843 15623
rect 7843 15589 7877 15623
rect 7877 15589 7892 15623
rect 7840 15580 7892 15589
rect 10876 15580 10928 15632
rect 11336 15623 11388 15632
rect 11336 15589 11345 15623
rect 11345 15589 11379 15623
rect 11379 15589 11388 15623
rect 11336 15580 11388 15589
rect 12348 15623 12400 15632
rect 12348 15589 12357 15623
rect 12357 15589 12391 15623
rect 12391 15589 12400 15623
rect 12348 15580 12400 15589
rect 16212 15580 16264 15632
rect 17040 15580 17092 15632
rect 17500 15623 17552 15632
rect 17500 15589 17509 15623
rect 17509 15589 17543 15623
rect 17543 15589 17552 15623
rect 17500 15580 17552 15589
rect 18972 15623 19024 15632
rect 18972 15589 18981 15623
rect 18981 15589 19015 15623
rect 19015 15589 19024 15623
rect 18972 15580 19024 15589
rect 19156 15580 19208 15632
rect 6000 15512 6052 15564
rect 8392 15555 8444 15564
rect 5448 15444 5500 15496
rect 8392 15521 8401 15555
rect 8401 15521 8435 15555
rect 8435 15521 8444 15555
rect 8392 15512 8444 15521
rect 13728 15555 13780 15564
rect 13728 15521 13772 15555
rect 13772 15521 13780 15555
rect 13728 15512 13780 15521
rect 7012 15444 7064 15496
rect 8208 15444 8260 15496
rect 10692 15487 10744 15496
rect 10692 15453 10701 15487
rect 10701 15453 10735 15487
rect 10735 15453 10744 15487
rect 10692 15444 10744 15453
rect 15568 15487 15620 15496
rect 15568 15453 15577 15487
rect 15577 15453 15611 15487
rect 15611 15453 15620 15487
rect 15568 15444 15620 15453
rect 16948 15444 17000 15496
rect 17868 15444 17920 15496
rect 5540 15376 5592 15428
rect 12440 15376 12492 15428
rect 18880 15376 18932 15428
rect 19524 15419 19576 15428
rect 19524 15385 19533 15419
rect 19533 15385 19567 15419
rect 19567 15385 19576 15419
rect 19524 15376 19576 15385
rect 15292 15308 15344 15360
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 7840 15104 7892 15156
rect 8300 15104 8352 15156
rect 10508 15147 10560 15156
rect 10508 15113 10517 15147
rect 10517 15113 10551 15147
rect 10551 15113 10560 15147
rect 10508 15104 10560 15113
rect 11244 15147 11296 15156
rect 11244 15113 11253 15147
rect 11253 15113 11287 15147
rect 11287 15113 11296 15147
rect 11244 15104 11296 15113
rect 13728 15147 13780 15156
rect 13728 15113 13737 15147
rect 13737 15113 13771 15147
rect 13771 15113 13780 15147
rect 13728 15104 13780 15113
rect 14832 15147 14884 15156
rect 14832 15113 14841 15147
rect 14841 15113 14875 15147
rect 14875 15113 14884 15147
rect 14832 15104 14884 15113
rect 16212 15104 16264 15156
rect 17500 15147 17552 15156
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 17960 15104 18012 15156
rect 19156 15104 19208 15156
rect 19984 15104 20036 15156
rect 7104 15036 7156 15088
rect 10232 15036 10284 15088
rect 11060 15036 11112 15088
rect 11152 15036 11204 15088
rect 12440 15036 12492 15088
rect 13176 15036 13228 15088
rect 5540 14968 5592 15020
rect 7748 14968 7800 15020
rect 9588 15011 9640 15020
rect 9588 14977 9597 15011
rect 9597 14977 9631 15011
rect 9631 14977 9640 15011
rect 9588 14968 9640 14977
rect 12348 14968 12400 15020
rect 13544 14968 13596 15020
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 11336 14943 11388 14952
rect 7840 14832 7892 14884
rect 5448 14764 5500 14816
rect 6644 14807 6696 14816
rect 6644 14773 6653 14807
rect 6653 14773 6687 14807
rect 6687 14773 6696 14807
rect 6644 14764 6696 14773
rect 7564 14764 7616 14816
rect 11336 14909 11345 14943
rect 11345 14909 11379 14943
rect 11379 14909 11388 14943
rect 11336 14900 11388 14909
rect 14832 14900 14884 14952
rect 15476 14943 15528 14952
rect 15476 14909 15485 14943
rect 15485 14909 15519 14943
rect 15519 14909 15528 14943
rect 15476 14900 15528 14909
rect 15844 14943 15896 14952
rect 15844 14909 15853 14943
rect 15853 14909 15887 14943
rect 15887 14909 15896 14943
rect 15844 14900 15896 14909
rect 16212 14943 16264 14952
rect 16212 14909 16221 14943
rect 16221 14909 16255 14943
rect 16255 14909 16264 14943
rect 16212 14900 16264 14909
rect 10232 14832 10284 14884
rect 10876 14875 10928 14884
rect 10876 14841 10885 14875
rect 10885 14841 10919 14875
rect 10919 14841 10928 14875
rect 10876 14832 10928 14841
rect 12716 14764 12768 14816
rect 14096 14764 14148 14816
rect 15660 14807 15712 14816
rect 15660 14773 15669 14807
rect 15669 14773 15703 14807
rect 15703 14773 15712 14807
rect 15660 14764 15712 14773
rect 20720 14900 20772 14952
rect 23572 14900 23624 14952
rect 19064 14832 19116 14884
rect 21180 14832 21232 14884
rect 24216 14832 24268 14884
rect 17592 14764 17644 14816
rect 18420 14807 18472 14816
rect 18420 14773 18429 14807
rect 18429 14773 18463 14807
rect 18463 14773 18472 14807
rect 18420 14764 18472 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 7840 14560 7892 14612
rect 10692 14560 10744 14612
rect 12716 14603 12768 14612
rect 12716 14569 12725 14603
rect 12725 14569 12759 14603
rect 12759 14569 12768 14603
rect 12716 14560 12768 14569
rect 15752 14560 15804 14612
rect 18972 14603 19024 14612
rect 18972 14569 18981 14603
rect 18981 14569 19015 14603
rect 19015 14569 19024 14603
rect 18972 14560 19024 14569
rect 19156 14560 19208 14612
rect 7012 14535 7064 14544
rect 7012 14501 7021 14535
rect 7021 14501 7055 14535
rect 7055 14501 7064 14535
rect 7012 14492 7064 14501
rect 8392 14492 8444 14544
rect 11060 14492 11112 14544
rect 11704 14535 11756 14544
rect 11704 14501 11707 14535
rect 11707 14501 11741 14535
rect 11741 14501 11756 14535
rect 11704 14492 11756 14501
rect 13452 14535 13504 14544
rect 13452 14501 13455 14535
rect 13455 14501 13489 14535
rect 13489 14501 13504 14535
rect 13452 14492 13504 14501
rect 18420 14492 18472 14544
rect 19340 14535 19392 14544
rect 19340 14501 19349 14535
rect 19349 14501 19383 14535
rect 19383 14501 19392 14535
rect 19340 14492 19392 14501
rect 19984 14535 20036 14544
rect 19984 14501 19993 14535
rect 19993 14501 20027 14535
rect 20027 14501 20036 14535
rect 19984 14492 20036 14501
rect 21180 14492 21232 14544
rect 5356 14424 5408 14476
rect 6552 14467 6604 14476
rect 6552 14433 6561 14467
rect 6561 14433 6595 14467
rect 6595 14433 6604 14467
rect 6552 14424 6604 14433
rect 7104 14424 7156 14476
rect 13084 14467 13136 14476
rect 13084 14433 13093 14467
rect 13093 14433 13127 14467
rect 13127 14433 13136 14467
rect 13084 14424 13136 14433
rect 14648 14424 14700 14476
rect 16580 14467 16632 14476
rect 16580 14433 16589 14467
rect 16589 14433 16623 14467
rect 16623 14433 16632 14467
rect 16580 14424 16632 14433
rect 16672 14424 16724 14476
rect 17040 14424 17092 14476
rect 17592 14467 17644 14476
rect 17592 14433 17601 14467
rect 17601 14433 17635 14467
rect 17635 14433 17644 14467
rect 17592 14424 17644 14433
rect 7472 14356 7524 14408
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 8392 14288 8444 14340
rect 10692 14356 10744 14408
rect 11980 14356 12032 14408
rect 17960 14356 18012 14408
rect 20996 14399 21048 14408
rect 20996 14365 21005 14399
rect 21005 14365 21039 14399
rect 21039 14365 21048 14399
rect 20996 14356 21048 14365
rect 21272 14399 21324 14408
rect 21272 14365 21281 14399
rect 21281 14365 21315 14399
rect 21315 14365 21324 14399
rect 21272 14356 21324 14365
rect 6000 14263 6052 14272
rect 6000 14229 6009 14263
rect 6009 14229 6043 14263
rect 6043 14229 6052 14263
rect 6000 14220 6052 14229
rect 6828 14220 6880 14272
rect 9128 14220 9180 14272
rect 11152 14263 11204 14272
rect 11152 14229 11161 14263
rect 11161 14229 11195 14263
rect 11195 14229 11204 14263
rect 11152 14220 11204 14229
rect 12256 14263 12308 14272
rect 12256 14229 12265 14263
rect 12265 14229 12299 14263
rect 12299 14229 12308 14263
rect 12256 14220 12308 14229
rect 12808 14220 12860 14272
rect 14740 14263 14792 14272
rect 14740 14229 14749 14263
rect 14749 14229 14783 14263
rect 14783 14229 14792 14263
rect 14740 14220 14792 14229
rect 15476 14220 15528 14272
rect 15844 14220 15896 14272
rect 16672 14220 16724 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 4160 14059 4212 14068
rect 4160 14025 4169 14059
rect 4169 14025 4203 14059
rect 4203 14025 4212 14059
rect 4160 14016 4212 14025
rect 6276 14016 6328 14068
rect 6552 14016 6604 14068
rect 7104 14059 7156 14068
rect 7104 14025 7113 14059
rect 7113 14025 7147 14059
rect 7147 14025 7156 14059
rect 7104 14016 7156 14025
rect 8484 14016 8536 14068
rect 9036 14059 9088 14068
rect 9036 14025 9045 14059
rect 9045 14025 9079 14059
rect 9079 14025 9088 14059
rect 9036 14016 9088 14025
rect 9864 14016 9916 14068
rect 10600 14059 10652 14068
rect 10600 14025 10609 14059
rect 10609 14025 10643 14059
rect 10643 14025 10652 14059
rect 10600 14016 10652 14025
rect 14648 14016 14700 14068
rect 16304 14016 16356 14068
rect 11428 13991 11480 14000
rect 11428 13957 11437 13991
rect 11437 13957 11471 13991
rect 11471 13957 11480 13991
rect 11428 13948 11480 13957
rect 15844 13948 15896 14000
rect 6368 13880 6420 13932
rect 6552 13880 6604 13932
rect 8024 13880 8076 13932
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 9680 13923 9732 13932
rect 9680 13889 9689 13923
rect 9689 13889 9723 13923
rect 9723 13889 9732 13923
rect 9680 13880 9732 13889
rect 9956 13880 10008 13932
rect 11152 13880 11204 13932
rect 12808 13880 12860 13932
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 14004 13880 14056 13932
rect 14648 13880 14700 13932
rect 15292 13880 15344 13932
rect 4160 13812 4212 13864
rect 4896 13812 4948 13864
rect 5356 13855 5408 13864
rect 5356 13821 5365 13855
rect 5365 13821 5399 13855
rect 5399 13821 5408 13855
rect 5356 13812 5408 13821
rect 7564 13855 7616 13864
rect 7564 13821 7573 13855
rect 7573 13821 7607 13855
rect 7607 13821 7616 13855
rect 7564 13812 7616 13821
rect 9220 13855 9272 13864
rect 9220 13821 9229 13855
rect 9229 13821 9263 13855
rect 9263 13821 9272 13855
rect 9220 13812 9272 13821
rect 4344 13787 4396 13796
rect 4344 13753 4353 13787
rect 4353 13753 4387 13787
rect 4387 13753 4396 13787
rect 4344 13744 4396 13753
rect 9128 13744 9180 13796
rect 10600 13812 10652 13864
rect 14740 13812 14792 13864
rect 15476 13855 15528 13864
rect 12440 13744 12492 13796
rect 12808 13787 12860 13796
rect 12808 13753 12817 13787
rect 12817 13753 12851 13787
rect 12851 13753 12860 13787
rect 15476 13821 15485 13855
rect 15485 13821 15519 13855
rect 15519 13821 15528 13855
rect 15476 13812 15528 13821
rect 15844 13855 15896 13864
rect 15844 13821 15853 13855
rect 15853 13821 15887 13855
rect 15887 13821 15896 13855
rect 15844 13812 15896 13821
rect 16212 13880 16264 13932
rect 12808 13744 12860 13753
rect 11244 13676 11296 13728
rect 11704 13676 11756 13728
rect 13452 13676 13504 13728
rect 14372 13719 14424 13728
rect 14372 13685 14381 13719
rect 14381 13685 14415 13719
rect 14415 13685 14424 13719
rect 14372 13676 14424 13685
rect 15568 13744 15620 13796
rect 16672 13812 16724 13864
rect 16856 13744 16908 13796
rect 19064 14016 19116 14068
rect 19156 14016 19208 14068
rect 19340 14016 19392 14068
rect 21180 14059 21232 14068
rect 21180 14025 21189 14059
rect 21189 14025 21223 14059
rect 21223 14025 21232 14059
rect 21180 14016 21232 14025
rect 19984 13880 20036 13932
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 18880 13744 18932 13796
rect 20904 13855 20956 13864
rect 20904 13821 20913 13855
rect 20913 13821 20947 13855
rect 20947 13821 20956 13855
rect 21548 13855 21600 13864
rect 20904 13812 20956 13821
rect 21548 13821 21557 13855
rect 21557 13821 21591 13855
rect 21591 13821 21600 13855
rect 21548 13812 21600 13821
rect 20720 13744 20772 13796
rect 17040 13719 17092 13728
rect 17040 13685 17049 13719
rect 17049 13685 17083 13719
rect 17083 13685 17092 13719
rect 17040 13676 17092 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 9864 13472 9916 13524
rect 10048 13472 10100 13524
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 13084 13472 13136 13524
rect 14372 13515 14424 13524
rect 14372 13481 14381 13515
rect 14381 13481 14415 13515
rect 14415 13481 14424 13515
rect 14372 13472 14424 13481
rect 15476 13472 15528 13524
rect 19524 13472 19576 13524
rect 19984 13472 20036 13524
rect 4160 13404 4212 13456
rect 4620 13336 4672 13388
rect 11244 13404 11296 13456
rect 12256 13404 12308 13456
rect 18052 13447 18104 13456
rect 18052 13413 18061 13447
rect 18061 13413 18095 13447
rect 18095 13413 18104 13447
rect 18052 13404 18104 13413
rect 18880 13404 18932 13456
rect 20720 13404 20772 13456
rect 7288 13379 7340 13388
rect 7288 13345 7297 13379
rect 7297 13345 7331 13379
rect 7331 13345 7340 13379
rect 7288 13336 7340 13345
rect 8760 13336 8812 13388
rect 14372 13336 14424 13388
rect 15476 13336 15528 13388
rect 16580 13379 16632 13388
rect 16580 13345 16589 13379
rect 16589 13345 16623 13379
rect 16623 13345 16632 13379
rect 16580 13336 16632 13345
rect 16672 13336 16724 13388
rect 16856 13336 16908 13388
rect 17040 13336 17092 13388
rect 4344 13268 4396 13320
rect 5264 13268 5316 13320
rect 5540 13268 5592 13320
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 11428 13268 11480 13320
rect 12072 13268 12124 13320
rect 12716 13268 12768 13320
rect 12992 13268 13044 13320
rect 14004 13268 14056 13320
rect 15292 13268 15344 13320
rect 16948 13268 17000 13320
rect 17960 13336 18012 13388
rect 20996 13379 21048 13388
rect 20996 13345 21005 13379
rect 21005 13345 21039 13379
rect 21039 13345 21048 13379
rect 20996 13336 21048 13345
rect 8024 13200 8076 13252
rect 8576 13200 8628 13252
rect 9220 13243 9272 13252
rect 9220 13209 9229 13243
rect 9229 13209 9263 13243
rect 9263 13209 9272 13243
rect 9220 13200 9272 13209
rect 12532 13200 12584 13252
rect 8116 13175 8168 13184
rect 8116 13141 8125 13175
rect 8125 13141 8159 13175
rect 8159 13141 8168 13175
rect 8116 13132 8168 13141
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 9128 13132 9180 13184
rect 11704 13175 11756 13184
rect 11704 13141 11713 13175
rect 11713 13141 11747 13175
rect 11747 13141 11756 13175
rect 11704 13132 11756 13141
rect 11980 13175 12032 13184
rect 11980 13141 11989 13175
rect 11989 13141 12023 13175
rect 12023 13141 12032 13175
rect 11980 13132 12032 13141
rect 14464 13132 14516 13184
rect 15568 13200 15620 13252
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 4160 12928 4212 12980
rect 5264 12928 5316 12980
rect 7288 12928 7340 12980
rect 8760 12971 8812 12980
rect 8760 12937 8769 12971
rect 8769 12937 8803 12971
rect 8803 12937 8812 12971
rect 8760 12928 8812 12937
rect 10140 12971 10192 12980
rect 10140 12937 10149 12971
rect 10149 12937 10183 12971
rect 10183 12937 10192 12971
rect 10140 12928 10192 12937
rect 11704 12928 11756 12980
rect 12624 12928 12676 12980
rect 16028 12928 16080 12980
rect 16580 12928 16632 12980
rect 17960 12928 18012 12980
rect 18788 12928 18840 12980
rect 19248 12928 19300 12980
rect 20996 12971 21048 12980
rect 20996 12937 21005 12971
rect 21005 12937 21039 12971
rect 21039 12937 21048 12971
rect 20996 12928 21048 12937
rect 6920 12860 6972 12912
rect 2872 12699 2924 12708
rect 2872 12665 2881 12699
rect 2881 12665 2915 12699
rect 2915 12665 2924 12699
rect 2872 12656 2924 12665
rect 2596 12631 2648 12640
rect 2596 12597 2605 12631
rect 2605 12597 2639 12631
rect 2639 12597 2648 12631
rect 2596 12588 2648 12597
rect 3608 12631 3660 12640
rect 3608 12597 3617 12631
rect 3617 12597 3651 12631
rect 3651 12597 3660 12631
rect 3608 12588 3660 12597
rect 4436 12724 4488 12776
rect 8484 12860 8536 12912
rect 8300 12835 8352 12844
rect 8300 12801 8309 12835
rect 8309 12801 8343 12835
rect 8343 12801 8352 12835
rect 8300 12792 8352 12801
rect 5172 12699 5224 12708
rect 5172 12665 5181 12699
rect 5181 12665 5215 12699
rect 5215 12665 5224 12699
rect 5172 12656 5224 12665
rect 7564 12699 7616 12708
rect 7564 12665 7573 12699
rect 7573 12665 7607 12699
rect 7607 12665 7616 12699
rect 8116 12724 8168 12776
rect 9036 12724 9088 12776
rect 12256 12903 12308 12912
rect 12256 12869 12265 12903
rect 12265 12869 12299 12903
rect 12299 12869 12308 12903
rect 12256 12860 12308 12869
rect 13728 12860 13780 12912
rect 9404 12724 9456 12776
rect 10048 12724 10100 12776
rect 11980 12792 12032 12844
rect 12532 12835 12584 12844
rect 12532 12801 12541 12835
rect 12541 12801 12575 12835
rect 12575 12801 12584 12835
rect 12532 12792 12584 12801
rect 12716 12792 12768 12844
rect 13452 12835 13504 12844
rect 13452 12801 13461 12835
rect 13461 12801 13495 12835
rect 13495 12801 13504 12835
rect 20260 12860 20312 12912
rect 13452 12792 13504 12801
rect 14372 12767 14424 12776
rect 14372 12733 14381 12767
rect 14381 12733 14415 12767
rect 14415 12733 14424 12767
rect 14372 12724 14424 12733
rect 15292 12767 15344 12776
rect 7564 12656 7616 12665
rect 12624 12699 12676 12708
rect 12624 12665 12633 12699
rect 12633 12665 12667 12699
rect 12667 12665 12676 12699
rect 12624 12656 12676 12665
rect 4068 12588 4120 12640
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 9496 12631 9548 12640
rect 9496 12597 9505 12631
rect 9505 12597 9539 12631
rect 9539 12597 9548 12631
rect 9496 12588 9548 12597
rect 10048 12588 10100 12640
rect 10968 12588 11020 12640
rect 11244 12588 11296 12640
rect 13820 12631 13872 12640
rect 13820 12597 13829 12631
rect 13829 12597 13863 12631
rect 13863 12597 13872 12631
rect 13820 12588 13872 12597
rect 14188 12631 14240 12640
rect 14188 12597 14197 12631
rect 14197 12597 14231 12631
rect 14231 12597 14240 12631
rect 15292 12733 15301 12767
rect 15301 12733 15335 12767
rect 15335 12733 15344 12767
rect 15292 12724 15344 12733
rect 15568 12767 15620 12776
rect 15568 12733 15577 12767
rect 15577 12733 15611 12767
rect 15611 12733 15620 12767
rect 15568 12724 15620 12733
rect 16948 12724 17000 12776
rect 19524 12792 19576 12844
rect 20628 12835 20680 12844
rect 20628 12801 20637 12835
rect 20637 12801 20671 12835
rect 20671 12801 20680 12835
rect 20628 12792 20680 12801
rect 21364 12724 21416 12776
rect 22468 12767 22520 12776
rect 22468 12733 22512 12767
rect 22512 12733 22520 12767
rect 22468 12724 22520 12733
rect 15844 12699 15896 12708
rect 15844 12665 15853 12699
rect 15853 12665 15887 12699
rect 15887 12665 15896 12699
rect 15844 12656 15896 12665
rect 14188 12588 14240 12597
rect 15568 12588 15620 12640
rect 16856 12656 16908 12708
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 20996 12656 21048 12708
rect 21180 12588 21232 12640
rect 22652 12588 22704 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 4160 12384 4212 12436
rect 12072 12427 12124 12436
rect 12072 12393 12081 12427
rect 12081 12393 12115 12427
rect 12115 12393 12124 12427
rect 12072 12384 12124 12393
rect 13820 12384 13872 12436
rect 15292 12384 15344 12436
rect 20904 12384 20956 12436
rect 24768 12427 24820 12436
rect 2688 12291 2740 12300
rect 2688 12257 2697 12291
rect 2697 12257 2731 12291
rect 2731 12257 2740 12291
rect 2688 12248 2740 12257
rect 4620 12248 4672 12300
rect 6184 12316 6236 12368
rect 7564 12359 7616 12368
rect 7564 12325 7573 12359
rect 7573 12325 7607 12359
rect 7607 12325 7616 12359
rect 7564 12316 7616 12325
rect 4896 12291 4948 12300
rect 4896 12257 4905 12291
rect 4905 12257 4939 12291
rect 4939 12257 4948 12291
rect 4896 12248 4948 12257
rect 2044 12180 2096 12232
rect 4160 12180 4212 12232
rect 5172 12248 5224 12300
rect 5540 12248 5592 12300
rect 6368 12291 6420 12300
rect 6368 12257 6377 12291
rect 6377 12257 6411 12291
rect 6411 12257 6420 12291
rect 6368 12248 6420 12257
rect 7196 12291 7248 12300
rect 7196 12257 7205 12291
rect 7205 12257 7239 12291
rect 7239 12257 7248 12291
rect 7196 12248 7248 12257
rect 8300 12248 8352 12300
rect 9036 12248 9088 12300
rect 9680 12248 9732 12300
rect 10048 12248 10100 12300
rect 10140 12248 10192 12300
rect 10416 12291 10468 12300
rect 10416 12257 10425 12291
rect 10425 12257 10459 12291
rect 10459 12257 10468 12291
rect 10416 12248 10468 12257
rect 11520 12291 11572 12300
rect 11520 12257 11564 12291
rect 11564 12257 11572 12291
rect 11520 12248 11572 12257
rect 12164 12248 12216 12300
rect 13360 12291 13412 12300
rect 13360 12257 13369 12291
rect 13369 12257 13403 12291
rect 13403 12257 13412 12291
rect 13360 12248 13412 12257
rect 10784 12180 10836 12232
rect 11704 12180 11756 12232
rect 14004 12248 14056 12300
rect 14464 12316 14516 12368
rect 18880 12316 18932 12368
rect 24768 12393 24777 12427
rect 24777 12393 24811 12427
rect 24811 12393 24820 12427
rect 24768 12384 24820 12393
rect 15292 12291 15344 12300
rect 15292 12257 15301 12291
rect 15301 12257 15335 12291
rect 15335 12257 15344 12291
rect 15292 12248 15344 12257
rect 16764 12291 16816 12300
rect 2504 12155 2556 12164
rect 2504 12121 2513 12155
rect 2513 12121 2547 12155
rect 2547 12121 2556 12155
rect 2504 12112 2556 12121
rect 8760 12155 8812 12164
rect 8760 12121 8769 12155
rect 8769 12121 8803 12155
rect 8803 12121 8812 12155
rect 8760 12112 8812 12121
rect 15476 12180 15528 12232
rect 16028 12180 16080 12232
rect 16764 12257 16773 12291
rect 16773 12257 16807 12291
rect 16807 12257 16816 12291
rect 16764 12248 16816 12257
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 17500 12291 17552 12300
rect 17500 12257 17509 12291
rect 17509 12257 17543 12291
rect 17543 12257 17552 12291
rect 17500 12248 17552 12257
rect 18788 12291 18840 12300
rect 18788 12257 18797 12291
rect 18797 12257 18831 12291
rect 18831 12257 18840 12291
rect 18788 12248 18840 12257
rect 22468 12291 22520 12300
rect 22468 12257 22512 12291
rect 22512 12257 22520 12291
rect 22468 12248 22520 12257
rect 20996 12223 21048 12232
rect 20996 12189 21005 12223
rect 21005 12189 21039 12223
rect 21039 12189 21048 12223
rect 20996 12180 21048 12189
rect 21088 12180 21140 12232
rect 14280 12155 14332 12164
rect 14280 12121 14289 12155
rect 14289 12121 14323 12155
rect 14323 12121 14332 12155
rect 14280 12112 14332 12121
rect 17684 12155 17736 12164
rect 17684 12121 17693 12155
rect 17693 12121 17727 12155
rect 17727 12121 17736 12155
rect 17684 12112 17736 12121
rect 6552 12087 6604 12096
rect 6552 12053 6561 12087
rect 6561 12053 6595 12087
rect 6595 12053 6604 12087
rect 6552 12044 6604 12053
rect 11428 12044 11480 12096
rect 12440 12087 12492 12096
rect 12440 12053 12449 12087
rect 12449 12053 12483 12087
rect 12483 12053 12492 12087
rect 12440 12044 12492 12053
rect 12624 12044 12676 12096
rect 14372 12044 14424 12096
rect 14648 12087 14700 12096
rect 14648 12053 14657 12087
rect 14657 12053 14691 12087
rect 14691 12053 14700 12087
rect 14648 12044 14700 12053
rect 16396 12044 16448 12096
rect 19524 12044 19576 12096
rect 22192 12044 22244 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2504 11840 2556 11892
rect 2688 11840 2740 11892
rect 4160 11883 4212 11892
rect 4160 11849 4169 11883
rect 4169 11849 4203 11883
rect 4203 11849 4212 11883
rect 4160 11840 4212 11849
rect 4436 11883 4488 11892
rect 4436 11849 4445 11883
rect 4445 11849 4479 11883
rect 4479 11849 4488 11883
rect 4436 11840 4488 11849
rect 4804 11772 4856 11824
rect 2044 11679 2096 11688
rect 2044 11645 2053 11679
rect 2053 11645 2087 11679
rect 2087 11645 2096 11679
rect 2044 11636 2096 11645
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 6184 11840 6236 11892
rect 6368 11883 6420 11892
rect 6368 11849 6377 11883
rect 6377 11849 6411 11883
rect 6411 11849 6420 11883
rect 6368 11840 6420 11849
rect 8300 11883 8352 11892
rect 8300 11849 8309 11883
rect 8309 11849 8343 11883
rect 8343 11849 8352 11883
rect 8300 11840 8352 11849
rect 8576 11883 8628 11892
rect 8576 11849 8585 11883
rect 8585 11849 8619 11883
rect 8619 11849 8628 11883
rect 8576 11840 8628 11849
rect 10416 11840 10468 11892
rect 11520 11840 11572 11892
rect 12900 11840 12952 11892
rect 13360 11840 13412 11892
rect 14188 11883 14240 11892
rect 14188 11849 14197 11883
rect 14197 11849 14231 11883
rect 14231 11849 14240 11883
rect 14188 11840 14240 11849
rect 18880 11840 18932 11892
rect 20996 11840 21048 11892
rect 7840 11772 7892 11824
rect 8760 11772 8812 11824
rect 5356 11747 5408 11756
rect 5356 11713 5365 11747
rect 5365 11713 5399 11747
rect 5399 11713 5408 11747
rect 5356 11704 5408 11713
rect 8208 11704 8260 11756
rect 17500 11815 17552 11824
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 7380 11636 7432 11688
rect 8576 11636 8628 11688
rect 9036 11679 9088 11688
rect 9036 11645 9045 11679
rect 9045 11645 9079 11679
rect 9079 11645 9088 11679
rect 9036 11636 9088 11645
rect 11704 11636 11756 11688
rect 12072 11636 12124 11688
rect 13636 11636 13688 11688
rect 14648 11679 14700 11688
rect 14648 11645 14657 11679
rect 14657 11645 14691 11679
rect 14691 11645 14700 11679
rect 14648 11636 14700 11645
rect 17500 11781 17509 11815
rect 17509 11781 17543 11815
rect 17543 11781 17552 11815
rect 17500 11772 17552 11781
rect 15384 11679 15436 11688
rect 4804 11568 4856 11620
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 2872 11543 2924 11552
rect 2872 11509 2881 11543
rect 2881 11509 2915 11543
rect 2915 11509 2924 11543
rect 2872 11500 2924 11509
rect 9496 11611 9548 11620
rect 9496 11577 9505 11611
rect 9505 11577 9539 11611
rect 9539 11577 9548 11611
rect 9496 11568 9548 11577
rect 13728 11568 13780 11620
rect 15384 11645 15393 11679
rect 15393 11645 15427 11679
rect 15427 11645 15436 11679
rect 15384 11636 15436 11645
rect 15752 11679 15804 11688
rect 15752 11645 15761 11679
rect 15761 11645 15795 11679
rect 15795 11645 15804 11679
rect 15752 11636 15804 11645
rect 16120 11568 16172 11620
rect 16764 11636 16816 11688
rect 18880 11568 18932 11620
rect 8392 11500 8444 11552
rect 9680 11500 9732 11552
rect 10968 11500 11020 11552
rect 12164 11543 12216 11552
rect 12164 11509 12173 11543
rect 12173 11509 12207 11543
rect 12207 11509 12216 11543
rect 12164 11500 12216 11509
rect 16580 11500 16632 11552
rect 20904 11543 20956 11552
rect 20904 11509 20913 11543
rect 20913 11509 20947 11543
rect 20947 11509 20956 11543
rect 20904 11500 20956 11509
rect 21088 11568 21140 11620
rect 22100 11611 22152 11620
rect 21364 11500 21416 11552
rect 22100 11577 22109 11611
rect 22109 11577 22143 11611
rect 22143 11577 22152 11611
rect 22100 11568 22152 11577
rect 22468 11543 22520 11552
rect 22468 11509 22477 11543
rect 22477 11509 22511 11543
rect 22511 11509 22520 11543
rect 22468 11500 22520 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 4804 11296 4856 11348
rect 6460 11296 6512 11348
rect 7932 11339 7984 11348
rect 7932 11305 7941 11339
rect 7941 11305 7975 11339
rect 7975 11305 7984 11339
rect 7932 11296 7984 11305
rect 9036 11339 9088 11348
rect 2228 11160 2280 11212
rect 2596 11160 2648 11212
rect 5448 11228 5500 11280
rect 7380 11271 7432 11280
rect 7380 11237 7389 11271
rect 7389 11237 7423 11271
rect 7423 11237 7432 11271
rect 9036 11305 9045 11339
rect 9045 11305 9079 11339
rect 9079 11305 9088 11339
rect 9036 11296 9088 11305
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 12072 11339 12124 11348
rect 12072 11305 12081 11339
rect 12081 11305 12115 11339
rect 12115 11305 12124 11339
rect 12072 11296 12124 11305
rect 12440 11339 12492 11348
rect 12440 11305 12449 11339
rect 12449 11305 12483 11339
rect 12483 11305 12492 11339
rect 12440 11296 12492 11305
rect 15384 11296 15436 11348
rect 15660 11296 15712 11348
rect 16672 11296 16724 11348
rect 18788 11339 18840 11348
rect 18788 11305 18797 11339
rect 18797 11305 18831 11339
rect 18831 11305 18840 11339
rect 18788 11296 18840 11305
rect 21364 11339 21416 11348
rect 21364 11305 21373 11339
rect 21373 11305 21407 11339
rect 21407 11305 21416 11339
rect 21364 11296 21416 11305
rect 7380 11228 7432 11237
rect 8760 11228 8812 11280
rect 9864 11228 9916 11280
rect 2044 11092 2096 11144
rect 4896 11160 4948 11212
rect 5264 11203 5316 11212
rect 5264 11169 5273 11203
rect 5273 11169 5307 11203
rect 5307 11169 5316 11203
rect 5264 11160 5316 11169
rect 6460 11160 6512 11212
rect 7840 11160 7892 11212
rect 10048 11203 10100 11212
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 6828 11092 6880 11144
rect 5080 11067 5132 11076
rect 5080 11033 5089 11067
rect 5089 11033 5123 11067
rect 5123 11033 5132 11067
rect 5080 11024 5132 11033
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 12256 11228 12308 11280
rect 9588 11092 9640 11144
rect 11060 11203 11112 11212
rect 11060 11169 11069 11203
rect 11069 11169 11103 11203
rect 11103 11169 11112 11203
rect 11060 11160 11112 11169
rect 12164 11203 12216 11212
rect 12164 11169 12173 11203
rect 12173 11169 12207 11203
rect 12207 11169 12216 11203
rect 12164 11160 12216 11169
rect 12900 11203 12952 11212
rect 12900 11169 12909 11203
rect 12909 11169 12943 11203
rect 12943 11169 12952 11203
rect 12900 11160 12952 11169
rect 15568 11228 15620 11280
rect 17132 11228 17184 11280
rect 13544 11203 13596 11212
rect 13544 11169 13553 11203
rect 13553 11169 13587 11203
rect 13587 11169 13596 11203
rect 13544 11160 13596 11169
rect 15292 11203 15344 11212
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 15292 11160 15344 11169
rect 16396 11160 16448 11212
rect 16580 11160 16632 11212
rect 20904 11228 20956 11280
rect 21916 11271 21968 11280
rect 21916 11237 21925 11271
rect 21925 11237 21959 11271
rect 21959 11237 21968 11271
rect 21916 11228 21968 11237
rect 22100 11228 22152 11280
rect 17500 11160 17552 11212
rect 19524 11203 19576 11212
rect 19524 11169 19533 11203
rect 19533 11169 19567 11203
rect 19567 11169 19576 11203
rect 19524 11160 19576 11169
rect 24124 11160 24176 11212
rect 21456 11092 21508 11144
rect 7932 10956 7984 11008
rect 9404 10956 9456 11008
rect 12256 11024 12308 11076
rect 14832 11024 14884 11076
rect 14004 10999 14056 11008
rect 14004 10965 14013 10999
rect 14013 10965 14047 10999
rect 14047 10965 14056 10999
rect 14004 10956 14056 10965
rect 18052 11024 18104 11076
rect 16948 10956 17000 11008
rect 24676 10956 24728 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2044 10795 2096 10804
rect 2044 10761 2053 10795
rect 2053 10761 2087 10795
rect 2087 10761 2096 10795
rect 2044 10752 2096 10761
rect 2228 10752 2280 10804
rect 2780 10752 2832 10804
rect 3148 10752 3200 10804
rect 7840 10752 7892 10804
rect 8392 10752 8444 10804
rect 9404 10752 9456 10804
rect 10048 10752 10100 10804
rect 12164 10752 12216 10804
rect 12256 10795 12308 10804
rect 12256 10761 12265 10795
rect 12265 10761 12299 10795
rect 12299 10761 12308 10795
rect 12256 10752 12308 10761
rect 12900 10752 12952 10804
rect 3700 10727 3752 10736
rect 3700 10693 3709 10727
rect 3709 10693 3743 10727
rect 3743 10693 3752 10727
rect 3700 10684 3752 10693
rect 8300 10684 8352 10736
rect 8484 10659 8536 10668
rect 3148 10548 3200 10600
rect 5540 10548 5592 10600
rect 5172 10480 5224 10532
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 8484 10625 8493 10659
rect 8493 10625 8527 10659
rect 8527 10625 8536 10659
rect 8484 10616 8536 10625
rect 10140 10616 10192 10668
rect 16580 10752 16632 10804
rect 19524 10752 19576 10804
rect 20536 10752 20588 10804
rect 21456 10795 21508 10804
rect 21456 10761 21465 10795
rect 21465 10761 21499 10795
rect 21499 10761 21508 10795
rect 21456 10752 21508 10761
rect 21916 10752 21968 10804
rect 24768 10795 24820 10804
rect 24768 10761 24777 10795
rect 24777 10761 24811 10795
rect 24811 10761 24820 10795
rect 24768 10752 24820 10761
rect 15292 10727 15344 10736
rect 15292 10693 15301 10727
rect 15301 10693 15335 10727
rect 15335 10693 15344 10727
rect 15292 10684 15344 10693
rect 6920 10548 6972 10557
rect 12164 10548 12216 10600
rect 13360 10591 13412 10600
rect 13360 10557 13369 10591
rect 13369 10557 13403 10591
rect 13403 10557 13412 10591
rect 13360 10548 13412 10557
rect 14004 10616 14056 10668
rect 17224 10616 17276 10668
rect 20444 10659 20496 10668
rect 20444 10625 20453 10659
rect 20453 10625 20487 10659
rect 20487 10625 20496 10659
rect 20444 10616 20496 10625
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 7564 10480 7616 10532
rect 8484 10480 8536 10532
rect 11244 10480 11296 10532
rect 2688 10455 2740 10464
rect 2688 10421 2697 10455
rect 2697 10421 2731 10455
rect 2731 10421 2740 10455
rect 2688 10412 2740 10421
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 4896 10412 4948 10464
rect 6644 10412 6696 10464
rect 7288 10455 7340 10464
rect 7288 10421 7297 10455
rect 7297 10421 7331 10455
rect 7331 10421 7340 10455
rect 7288 10412 7340 10421
rect 9680 10412 9732 10464
rect 11060 10412 11112 10464
rect 11704 10412 11756 10464
rect 12624 10480 12676 10532
rect 15476 10548 15528 10600
rect 16120 10591 16172 10600
rect 16120 10557 16129 10591
rect 16129 10557 16163 10591
rect 16163 10557 16172 10591
rect 16120 10548 16172 10557
rect 16672 10591 16724 10600
rect 16672 10557 16681 10591
rect 16681 10557 16715 10591
rect 16715 10557 16724 10591
rect 16672 10548 16724 10557
rect 16948 10591 17000 10600
rect 16948 10557 16957 10591
rect 16957 10557 16991 10591
rect 16991 10557 17000 10591
rect 16948 10548 17000 10557
rect 18972 10548 19024 10600
rect 21364 10548 21416 10600
rect 22008 10591 22060 10600
rect 22008 10557 22017 10591
rect 22017 10557 22051 10591
rect 22051 10557 22060 10591
rect 22008 10548 22060 10557
rect 24124 10548 24176 10600
rect 24308 10591 24360 10600
rect 24308 10557 24317 10591
rect 24317 10557 24351 10591
rect 24351 10557 24360 10591
rect 24308 10548 24360 10557
rect 24676 10548 24728 10600
rect 14832 10523 14884 10532
rect 14832 10489 14841 10523
rect 14841 10489 14875 10523
rect 14875 10489 14884 10523
rect 14832 10480 14884 10489
rect 16396 10480 16448 10532
rect 20536 10523 20588 10532
rect 20536 10489 20545 10523
rect 20545 10489 20579 10523
rect 20579 10489 20588 10523
rect 20536 10480 20588 10489
rect 13084 10412 13136 10464
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 19064 10455 19116 10464
rect 19064 10421 19073 10455
rect 19073 10421 19107 10455
rect 19107 10421 19116 10455
rect 19064 10412 19116 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 5080 10208 5132 10260
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 8392 10208 8444 10260
rect 10140 10208 10192 10260
rect 6460 10140 6512 10192
rect 6736 10140 6788 10192
rect 8116 10183 8168 10192
rect 8116 10149 8125 10183
rect 8125 10149 8159 10183
rect 8159 10149 8168 10183
rect 8116 10140 8168 10149
rect 8208 10183 8260 10192
rect 8208 10149 8217 10183
rect 8217 10149 8251 10183
rect 8251 10149 8260 10183
rect 8208 10140 8260 10149
rect 10048 10140 10100 10192
rect 12072 10208 12124 10260
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 13636 10251 13688 10260
rect 13636 10217 13645 10251
rect 13645 10217 13679 10251
rect 13679 10217 13688 10251
rect 13636 10208 13688 10217
rect 14924 10208 14976 10260
rect 16120 10208 16172 10260
rect 20444 10251 20496 10260
rect 20444 10217 20453 10251
rect 20453 10217 20487 10251
rect 20487 10217 20496 10251
rect 20444 10208 20496 10217
rect 22008 10251 22060 10260
rect 22008 10217 22017 10251
rect 22017 10217 22051 10251
rect 22051 10217 22060 10251
rect 22008 10208 22060 10217
rect 11888 10183 11940 10192
rect 11888 10149 11897 10183
rect 11897 10149 11931 10183
rect 11931 10149 11940 10183
rect 11888 10140 11940 10149
rect 13084 10183 13136 10192
rect 13084 10149 13087 10183
rect 13087 10149 13121 10183
rect 13121 10149 13136 10183
rect 13084 10140 13136 10149
rect 13360 10140 13412 10192
rect 2136 10072 2188 10124
rect 2596 10072 2648 10124
rect 3148 10115 3200 10124
rect 3148 10081 3157 10115
rect 3157 10081 3191 10115
rect 3191 10081 3200 10115
rect 3148 10072 3200 10081
rect 4896 10072 4948 10124
rect 5356 10072 5408 10124
rect 6644 10072 6696 10124
rect 7288 10072 7340 10124
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 9864 10072 9916 10124
rect 12440 10072 12492 10124
rect 13268 10072 13320 10124
rect 14004 10140 14056 10192
rect 15752 10140 15804 10192
rect 16948 10140 17000 10192
rect 17316 10140 17368 10192
rect 16396 10115 16448 10124
rect 16396 10081 16405 10115
rect 16405 10081 16439 10115
rect 16439 10081 16448 10115
rect 16396 10072 16448 10081
rect 16580 10072 16632 10124
rect 17224 10115 17276 10124
rect 17224 10081 17233 10115
rect 17233 10081 17267 10115
rect 17267 10081 17276 10115
rect 17224 10072 17276 10081
rect 18880 10140 18932 10192
rect 20812 10140 20864 10192
rect 18052 10072 18104 10124
rect 18604 10072 18656 10124
rect 22100 10072 22152 10124
rect 23112 10115 23164 10124
rect 23112 10081 23156 10115
rect 23156 10081 23164 10115
rect 23112 10072 23164 10081
rect 5172 10004 5224 10056
rect 8300 10004 8352 10056
rect 11520 10004 11572 10056
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 17960 10004 18012 10056
rect 20720 10004 20772 10056
rect 21732 10004 21784 10056
rect 2504 9979 2556 9988
rect 2504 9945 2513 9979
rect 2513 9945 2547 9979
rect 2547 9945 2556 9979
rect 2504 9936 2556 9945
rect 4988 9936 5040 9988
rect 6276 9936 6328 9988
rect 6920 9868 6972 9920
rect 7564 9868 7616 9920
rect 8484 9868 8536 9920
rect 9864 9911 9916 9920
rect 9864 9877 9873 9911
rect 9873 9877 9907 9911
rect 9907 9877 9916 9911
rect 9864 9868 9916 9877
rect 12164 9911 12216 9920
rect 12164 9877 12173 9911
rect 12173 9877 12207 9911
rect 12207 9877 12216 9911
rect 12164 9868 12216 9877
rect 13544 9868 13596 9920
rect 20812 9868 20864 9920
rect 23388 9868 23440 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2136 9707 2188 9716
rect 2136 9673 2145 9707
rect 2145 9673 2179 9707
rect 2179 9673 2188 9707
rect 2136 9664 2188 9673
rect 2504 9664 2556 9716
rect 5080 9664 5132 9716
rect 6644 9707 6696 9716
rect 6644 9673 6653 9707
rect 6653 9673 6687 9707
rect 6687 9673 6696 9707
rect 6644 9664 6696 9673
rect 6920 9664 6972 9716
rect 8116 9664 8168 9716
rect 9680 9664 9732 9716
rect 12072 9664 12124 9716
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 4988 9528 5040 9580
rect 9404 9596 9456 9648
rect 10968 9596 11020 9648
rect 13820 9639 13872 9648
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 14648 9639 14700 9648
rect 14648 9605 14657 9639
rect 14657 9605 14691 9639
rect 14691 9605 14700 9639
rect 14648 9596 14700 9605
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 14372 9528 14424 9580
rect 15292 9664 15344 9716
rect 15476 9707 15528 9716
rect 15476 9673 15485 9707
rect 15485 9673 15519 9707
rect 15519 9673 15528 9707
rect 15476 9664 15528 9673
rect 17316 9707 17368 9716
rect 17316 9673 17325 9707
rect 17325 9673 17359 9707
rect 17359 9673 17368 9707
rect 17316 9664 17368 9673
rect 18972 9707 19024 9716
rect 18972 9673 18981 9707
rect 18981 9673 19015 9707
rect 19015 9673 19024 9707
rect 18972 9664 19024 9673
rect 20720 9664 20772 9716
rect 23112 9707 23164 9716
rect 16488 9596 16540 9648
rect 17224 9596 17276 9648
rect 19984 9596 20036 9648
rect 20812 9639 20864 9648
rect 20812 9605 20821 9639
rect 20821 9605 20855 9639
rect 20855 9605 20864 9639
rect 20812 9596 20864 9605
rect 23112 9673 23121 9707
rect 23121 9673 23155 9707
rect 23155 9673 23164 9707
rect 23112 9664 23164 9673
rect 24768 9639 24820 9648
rect 24768 9605 24777 9639
rect 24777 9605 24811 9639
rect 24811 9605 24820 9639
rect 24768 9596 24820 9605
rect 17960 9528 18012 9580
rect 18880 9528 18932 9580
rect 20168 9571 20220 9580
rect 20168 9537 20177 9571
rect 20177 9537 20211 9571
rect 20211 9537 20220 9571
rect 20168 9528 20220 9537
rect 20720 9528 20772 9580
rect 21272 9528 21324 9580
rect 21732 9571 21784 9580
rect 21732 9537 21741 9571
rect 21741 9537 21775 9571
rect 21775 9537 21784 9571
rect 21732 9528 21784 9537
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 5356 9503 5408 9512
rect 5356 9469 5365 9503
rect 5365 9469 5399 9503
rect 5399 9469 5408 9503
rect 5356 9460 5408 9469
rect 9312 9503 9364 9512
rect 9312 9469 9321 9503
rect 9321 9469 9355 9503
rect 9355 9469 9364 9503
rect 9312 9460 9364 9469
rect 2596 9324 2648 9376
rect 4896 9367 4948 9376
rect 4896 9333 4905 9367
rect 4905 9333 4939 9367
rect 4939 9333 4948 9367
rect 4896 9324 4948 9333
rect 7012 9367 7064 9376
rect 7012 9333 7021 9367
rect 7021 9333 7055 9367
rect 7055 9333 7064 9367
rect 7012 9324 7064 9333
rect 10968 9435 11020 9444
rect 10968 9401 10977 9435
rect 10977 9401 11011 9435
rect 11011 9401 11020 9435
rect 11520 9435 11572 9444
rect 10968 9392 11020 9401
rect 11520 9401 11529 9435
rect 11529 9401 11563 9435
rect 11563 9401 11572 9435
rect 11520 9392 11572 9401
rect 8116 9324 8168 9376
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 8760 9324 8812 9333
rect 10784 9324 10836 9376
rect 11336 9324 11388 9376
rect 12256 9367 12308 9376
rect 12256 9333 12265 9367
rect 12265 9333 12299 9367
rect 12299 9333 12308 9367
rect 13820 9392 13872 9444
rect 16028 9435 16080 9444
rect 12256 9324 12308 9333
rect 13084 9324 13136 9376
rect 13728 9324 13780 9376
rect 16028 9401 16037 9435
rect 16037 9401 16071 9435
rect 16071 9401 16080 9435
rect 16028 9392 16080 9401
rect 16672 9435 16724 9444
rect 16672 9401 16681 9435
rect 16681 9401 16715 9435
rect 16715 9401 16724 9435
rect 16672 9392 16724 9401
rect 17868 9435 17920 9444
rect 17868 9401 17877 9435
rect 17877 9401 17911 9435
rect 17911 9401 17920 9435
rect 17868 9392 17920 9401
rect 24584 9503 24636 9512
rect 24584 9469 24593 9503
rect 24593 9469 24627 9503
rect 24627 9469 24636 9503
rect 24584 9460 24636 9469
rect 19524 9392 19576 9444
rect 19984 9435 20036 9444
rect 19984 9401 19993 9435
rect 19993 9401 20027 9435
rect 20027 9401 20036 9435
rect 19984 9392 20036 9401
rect 21548 9435 21600 9444
rect 21548 9401 21557 9435
rect 21557 9401 21591 9435
rect 21591 9401 21600 9435
rect 21548 9392 21600 9401
rect 16212 9324 16264 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 4988 9120 5040 9172
rect 7380 9120 7432 9172
rect 7748 9120 7800 9172
rect 8208 9120 8260 9172
rect 8576 9120 8628 9172
rect 8760 9120 8812 9172
rect 11336 9163 11388 9172
rect 11336 9129 11345 9163
rect 11345 9129 11379 9163
rect 11379 9129 11388 9163
rect 11336 9120 11388 9129
rect 13268 9163 13320 9172
rect 13268 9129 13277 9163
rect 13277 9129 13311 9163
rect 13311 9129 13320 9163
rect 13268 9120 13320 9129
rect 14004 9163 14056 9172
rect 14004 9129 14013 9163
rect 14013 9129 14047 9163
rect 14047 9129 14056 9163
rect 14004 9120 14056 9129
rect 14372 9163 14424 9172
rect 14372 9129 14381 9163
rect 14381 9129 14415 9163
rect 14415 9129 14424 9163
rect 14372 9120 14424 9129
rect 16028 9120 16080 9172
rect 16212 9163 16264 9172
rect 16212 9129 16221 9163
rect 16221 9129 16255 9163
rect 16255 9129 16264 9163
rect 16212 9120 16264 9129
rect 16580 9163 16632 9172
rect 16580 9129 16589 9163
rect 16589 9129 16623 9163
rect 16623 9129 16632 9163
rect 16580 9120 16632 9129
rect 17960 9120 18012 9172
rect 18604 9163 18656 9172
rect 18604 9129 18613 9163
rect 18613 9129 18647 9163
rect 18647 9129 18656 9163
rect 18604 9120 18656 9129
rect 24584 9120 24636 9172
rect 5356 9052 5408 9104
rect 8116 9052 8168 9104
rect 8392 9052 8444 9104
rect 9312 9052 9364 9104
rect 10140 9052 10192 9104
rect 12164 9052 12216 9104
rect 12992 9095 13044 9104
rect 12992 9061 13001 9095
rect 13001 9061 13035 9095
rect 13035 9061 13044 9095
rect 12992 9052 13044 9061
rect 15384 9052 15436 9104
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 5172 8984 5224 9036
rect 6092 9027 6144 9036
rect 6092 8993 6101 9027
rect 6101 8993 6135 9027
rect 6135 8993 6144 9027
rect 6092 8984 6144 8993
rect 11520 8984 11572 9036
rect 13544 8984 13596 9036
rect 14832 8984 14884 9036
rect 7840 8916 7892 8968
rect 10048 8916 10100 8968
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 10784 8848 10836 8900
rect 12532 8848 12584 8900
rect 18512 9052 18564 9104
rect 19064 9052 19116 9104
rect 20168 9052 20220 9104
rect 21088 9095 21140 9104
rect 21088 9061 21097 9095
rect 21097 9061 21131 9095
rect 21131 9061 21140 9095
rect 21088 9052 21140 9061
rect 17132 9027 17184 9036
rect 17132 8993 17141 9027
rect 17141 8993 17175 9027
rect 17175 8993 17184 9027
rect 17132 8984 17184 8993
rect 23572 9027 23624 9036
rect 23572 8993 23616 9027
rect 23616 8993 23624 9027
rect 23572 8984 23624 8993
rect 16212 8916 16264 8968
rect 20996 8959 21048 8968
rect 20996 8925 21005 8959
rect 21005 8925 21039 8959
rect 21039 8925 21048 8959
rect 20996 8916 21048 8925
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 17868 8848 17920 8900
rect 19524 8780 19576 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2596 8576 2648 8628
rect 4620 8576 4672 8628
rect 8668 8619 8720 8628
rect 8668 8585 8677 8619
rect 8677 8585 8711 8619
rect 8711 8585 8720 8619
rect 8668 8576 8720 8585
rect 13544 8576 13596 8628
rect 13728 8619 13780 8628
rect 13728 8585 13737 8619
rect 13737 8585 13771 8619
rect 13771 8585 13780 8619
rect 15384 8619 15436 8628
rect 13728 8576 13780 8585
rect 4988 8508 5040 8560
rect 4160 8372 4212 8424
rect 4896 8372 4948 8424
rect 6092 8440 6144 8492
rect 8116 8440 8168 8492
rect 10140 8508 10192 8560
rect 10048 8440 10100 8492
rect 14280 8440 14332 8492
rect 7380 8415 7432 8424
rect 7380 8381 7389 8415
rect 7389 8381 7423 8415
rect 7423 8381 7432 8415
rect 7380 8372 7432 8381
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 8668 8372 8720 8424
rect 9312 8415 9364 8424
rect 9312 8381 9321 8415
rect 9321 8381 9355 8415
rect 9355 8381 9364 8415
rect 9312 8372 9364 8381
rect 9680 8372 9732 8424
rect 10876 8372 10928 8424
rect 11336 8415 11388 8424
rect 11336 8381 11345 8415
rect 11345 8381 11379 8415
rect 11379 8381 11388 8415
rect 12164 8415 12216 8424
rect 11336 8372 11388 8381
rect 12164 8381 12173 8415
rect 12173 8381 12207 8415
rect 12207 8381 12216 8415
rect 12164 8372 12216 8381
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 12440 8372 12492 8381
rect 7840 8347 7892 8356
rect 7840 8313 7849 8347
rect 7849 8313 7883 8347
rect 7883 8313 7892 8347
rect 7840 8304 7892 8313
rect 8116 8279 8168 8288
rect 8116 8245 8125 8279
rect 8125 8245 8159 8279
rect 8159 8245 8168 8279
rect 8116 8236 8168 8245
rect 8208 8236 8260 8288
rect 9404 8304 9456 8356
rect 9588 8347 9640 8356
rect 9588 8313 9597 8347
rect 9597 8313 9631 8347
rect 9631 8313 9640 8347
rect 9588 8304 9640 8313
rect 10140 8304 10192 8356
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 17132 8619 17184 8628
rect 17132 8585 17141 8619
rect 17141 8585 17175 8619
rect 17175 8585 17184 8619
rect 17132 8576 17184 8585
rect 18512 8576 18564 8628
rect 19064 8576 19116 8628
rect 16672 8551 16724 8560
rect 16672 8517 16681 8551
rect 16681 8517 16715 8551
rect 16715 8517 16724 8551
rect 16672 8508 16724 8517
rect 19984 8576 20036 8628
rect 21548 8576 21600 8628
rect 23572 8576 23624 8628
rect 21088 8508 21140 8560
rect 16212 8440 16264 8492
rect 18788 8483 18840 8492
rect 18788 8449 18797 8483
rect 18797 8449 18831 8483
rect 18831 8449 18840 8483
rect 18788 8440 18840 8449
rect 19984 8440 20036 8492
rect 21272 8440 21324 8492
rect 15200 8372 15252 8424
rect 20812 8372 20864 8424
rect 21640 8372 21692 8424
rect 23480 8372 23532 8424
rect 16120 8347 16172 8356
rect 16120 8313 16129 8347
rect 16129 8313 16163 8347
rect 16163 8313 16172 8347
rect 16120 8304 16172 8313
rect 16212 8347 16264 8356
rect 16212 8313 16221 8347
rect 16221 8313 16255 8347
rect 16255 8313 16264 8347
rect 16212 8304 16264 8313
rect 20076 8304 20128 8356
rect 10968 8236 11020 8288
rect 24676 8236 24728 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 7564 8075 7616 8084
rect 5172 7939 5224 7948
rect 5172 7905 5181 7939
rect 5181 7905 5215 7939
rect 5215 7905 5224 7939
rect 5172 7896 5224 7905
rect 5540 7896 5592 7948
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 7840 8075 7892 8084
rect 7840 8041 7849 8075
rect 7849 8041 7883 8075
rect 7883 8041 7892 8075
rect 7840 8032 7892 8041
rect 10048 8075 10100 8084
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 10876 8075 10928 8084
rect 10876 8041 10885 8075
rect 10885 8041 10919 8075
rect 10919 8041 10928 8075
rect 10876 8032 10928 8041
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 14280 8032 14332 8084
rect 14832 8032 14884 8084
rect 19524 8032 19576 8084
rect 20996 8032 21048 8084
rect 21640 8032 21692 8084
rect 24768 8075 24820 8084
rect 24768 8041 24777 8075
rect 24777 8041 24811 8075
rect 24811 8041 24820 8075
rect 24768 8032 24820 8041
rect 6460 7939 6512 7948
rect 6460 7905 6469 7939
rect 6469 7905 6503 7939
rect 6503 7905 6512 7939
rect 6460 7896 6512 7905
rect 6552 7896 6604 7948
rect 7932 7896 7984 7948
rect 8208 7939 8260 7948
rect 8208 7905 8217 7939
rect 8217 7905 8251 7939
rect 8251 7905 8260 7939
rect 8208 7896 8260 7905
rect 8668 7896 8720 7948
rect 9312 7896 9364 7948
rect 9772 7939 9824 7948
rect 9772 7905 9781 7939
rect 9781 7905 9815 7939
rect 9815 7905 9824 7939
rect 9772 7896 9824 7905
rect 11428 8007 11480 8016
rect 11428 7973 11437 8007
rect 11437 7973 11471 8007
rect 11471 7973 11480 8007
rect 11428 7964 11480 7973
rect 11704 7964 11756 8016
rect 13820 8007 13872 8016
rect 13820 7973 13829 8007
rect 13829 7973 13863 8007
rect 13863 7973 13872 8007
rect 13820 7964 13872 7973
rect 15200 7964 15252 8016
rect 15476 8007 15528 8016
rect 15476 7973 15485 8007
rect 15485 7973 15519 8007
rect 15519 7973 15528 8007
rect 15476 7964 15528 7973
rect 16028 8007 16080 8016
rect 16028 7973 16037 8007
rect 16037 7973 16071 8007
rect 16071 7973 16080 8007
rect 16028 7964 16080 7973
rect 17868 7964 17920 8016
rect 10876 7896 10928 7948
rect 17684 7896 17736 7948
rect 21180 7896 21232 7948
rect 21732 7896 21784 7948
rect 24584 7939 24636 7948
rect 24584 7905 24593 7939
rect 24593 7905 24627 7939
rect 24627 7905 24636 7939
rect 24584 7896 24636 7905
rect 25412 7896 25464 7948
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 8760 7871 8812 7880
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 11520 7828 11572 7880
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 15384 7871 15436 7880
rect 15384 7837 15393 7871
rect 15393 7837 15427 7871
rect 15427 7837 15436 7871
rect 15384 7828 15436 7837
rect 19984 7828 20036 7880
rect 12440 7803 12492 7812
rect 12440 7769 12449 7803
rect 12449 7769 12483 7803
rect 12483 7769 12492 7803
rect 12440 7760 12492 7769
rect 16120 7760 16172 7812
rect 18972 7760 19024 7812
rect 9220 7735 9272 7744
rect 9220 7701 9229 7735
rect 9229 7701 9263 7735
rect 9263 7701 9272 7735
rect 9220 7692 9272 7701
rect 18880 7735 18932 7744
rect 18880 7701 18889 7735
rect 18889 7701 18923 7735
rect 18923 7701 18932 7735
rect 18880 7692 18932 7701
rect 19892 7735 19944 7744
rect 19892 7701 19901 7735
rect 19901 7701 19935 7735
rect 19935 7701 19944 7735
rect 19892 7692 19944 7701
rect 21272 7692 21324 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 5172 7488 5224 7540
rect 6552 7531 6604 7540
rect 6552 7497 6561 7531
rect 6561 7497 6595 7531
rect 6595 7497 6604 7531
rect 6552 7488 6604 7497
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 9772 7488 9824 7540
rect 11704 7531 11756 7540
rect 11704 7497 11713 7531
rect 11713 7497 11747 7531
rect 11747 7497 11756 7531
rect 11704 7488 11756 7497
rect 10508 7463 10560 7472
rect 10508 7429 10517 7463
rect 10517 7429 10551 7463
rect 10551 7429 10560 7463
rect 10508 7420 10560 7429
rect 8300 7352 8352 7404
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 9680 7395 9732 7404
rect 9680 7361 9689 7395
rect 9689 7361 9723 7395
rect 9723 7361 9732 7395
rect 9680 7352 9732 7361
rect 3700 7327 3752 7336
rect 3700 7293 3709 7327
rect 3709 7293 3743 7327
rect 3743 7293 3752 7327
rect 3700 7284 3752 7293
rect 2780 7216 2832 7268
rect 5080 7284 5132 7336
rect 5448 7327 5500 7336
rect 5448 7293 5457 7327
rect 5457 7293 5491 7327
rect 5491 7293 5500 7327
rect 5448 7284 5500 7293
rect 5540 7284 5592 7336
rect 7012 7284 7064 7336
rect 11244 7395 11296 7404
rect 11244 7361 11253 7395
rect 11253 7361 11287 7395
rect 11287 7361 11296 7395
rect 11244 7352 11296 7361
rect 10876 7284 10928 7336
rect 6184 7216 6236 7268
rect 3884 7191 3936 7200
rect 3884 7157 3893 7191
rect 3893 7157 3927 7191
rect 3927 7157 3936 7191
rect 3884 7148 3936 7157
rect 7104 7148 7156 7200
rect 8116 7216 8168 7268
rect 9128 7148 9180 7200
rect 11612 7148 11664 7200
rect 13084 7488 13136 7540
rect 15384 7488 15436 7540
rect 17684 7488 17736 7540
rect 20536 7488 20588 7540
rect 21180 7531 21232 7540
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 23480 7488 23532 7540
rect 25412 7531 25464 7540
rect 25412 7497 25421 7531
rect 25421 7497 25455 7531
rect 25455 7497 25464 7531
rect 25412 7488 25464 7497
rect 13728 7420 13780 7472
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 14924 7395 14976 7404
rect 12440 7352 12492 7361
rect 14924 7361 14933 7395
rect 14933 7361 14967 7395
rect 14967 7361 14976 7395
rect 14924 7352 14976 7361
rect 15200 7352 15252 7404
rect 15936 7395 15988 7404
rect 15936 7361 15945 7395
rect 15945 7361 15979 7395
rect 15979 7361 15988 7395
rect 15936 7352 15988 7361
rect 17868 7352 17920 7404
rect 18880 7395 18932 7404
rect 18880 7361 18889 7395
rect 18889 7361 18923 7395
rect 18923 7361 18932 7395
rect 18880 7352 18932 7361
rect 13728 7284 13780 7336
rect 13912 7284 13964 7336
rect 24676 7327 24728 7336
rect 24676 7293 24694 7327
rect 24694 7293 24728 7327
rect 24676 7284 24728 7293
rect 13084 7216 13136 7268
rect 13820 7216 13872 7268
rect 18972 7259 19024 7268
rect 18972 7225 18981 7259
rect 18981 7225 19015 7259
rect 19015 7225 19024 7259
rect 18972 7216 19024 7225
rect 19524 7259 19576 7268
rect 19524 7225 19533 7259
rect 19533 7225 19567 7259
rect 19567 7225 19576 7259
rect 19524 7216 19576 7225
rect 15292 7191 15344 7200
rect 15292 7157 15301 7191
rect 15301 7157 15335 7191
rect 15335 7157 15344 7191
rect 15292 7148 15344 7157
rect 15476 7148 15528 7200
rect 19984 7148 20036 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 3700 6987 3752 6996
rect 3700 6953 3709 6987
rect 3709 6953 3743 6987
rect 3743 6953 3752 6987
rect 6460 6987 6512 6996
rect 3700 6944 3752 6953
rect 6460 6953 6469 6987
rect 6469 6953 6503 6987
rect 6503 6953 6512 6987
rect 6460 6944 6512 6953
rect 7012 6944 7064 6996
rect 5080 6876 5132 6928
rect 7104 6876 7156 6928
rect 7932 6944 7984 6996
rect 9128 6987 9180 6996
rect 9128 6953 9137 6987
rect 9137 6953 9171 6987
rect 9171 6953 9180 6987
rect 9128 6944 9180 6953
rect 10876 6944 10928 6996
rect 11244 6944 11296 6996
rect 9864 6919 9916 6928
rect 5540 6808 5592 6860
rect 6000 6808 6052 6860
rect 6920 6851 6972 6860
rect 6920 6817 6929 6851
rect 6929 6817 6963 6851
rect 6963 6817 6972 6851
rect 6920 6808 6972 6817
rect 9864 6885 9873 6919
rect 9873 6885 9907 6919
rect 9907 6885 9916 6919
rect 9864 6876 9916 6885
rect 11612 6919 11664 6928
rect 11612 6885 11615 6919
rect 11615 6885 11649 6919
rect 11649 6885 11664 6919
rect 11612 6876 11664 6885
rect 13176 6919 13228 6928
rect 13176 6885 13185 6919
rect 13185 6885 13219 6919
rect 13219 6885 13228 6919
rect 13176 6876 13228 6885
rect 15476 6919 15528 6928
rect 15476 6885 15485 6919
rect 15485 6885 15519 6919
rect 15519 6885 15528 6919
rect 15476 6876 15528 6885
rect 16120 6876 16172 6928
rect 17408 6876 17460 6928
rect 17868 6876 17920 6928
rect 18788 6919 18840 6928
rect 18788 6885 18797 6919
rect 18797 6885 18831 6919
rect 18831 6885 18840 6919
rect 18788 6876 18840 6885
rect 11152 6808 11204 6860
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 16856 6851 16908 6860
rect 16856 6817 16865 6851
rect 16865 6817 16899 6851
rect 16899 6817 16908 6851
rect 16856 6808 16908 6817
rect 20996 6851 21048 6860
rect 20996 6817 21005 6851
rect 21005 6817 21039 6851
rect 21039 6817 21048 6851
rect 20996 6808 21048 6817
rect 6092 6783 6144 6792
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 9036 6740 9088 6792
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 13268 6740 13320 6792
rect 15384 6783 15436 6792
rect 12992 6672 13044 6724
rect 15384 6749 15393 6783
rect 15393 6749 15427 6783
rect 15427 6749 15436 6783
rect 15384 6740 15436 6749
rect 18696 6783 18748 6792
rect 18696 6749 18705 6783
rect 18705 6749 18739 6783
rect 18739 6749 18748 6783
rect 18696 6740 18748 6749
rect 18880 6740 18932 6792
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 14004 6672 14056 6724
rect 15108 6672 15160 6724
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 12164 6647 12216 6656
rect 12164 6613 12173 6647
rect 12173 6613 12207 6647
rect 12207 6613 12216 6647
rect 12164 6604 12216 6613
rect 14280 6647 14332 6656
rect 14280 6613 14289 6647
rect 14289 6613 14323 6647
rect 14323 6613 14332 6647
rect 14280 6604 14332 6613
rect 14832 6604 14884 6656
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 17960 6604 18012 6656
rect 19432 6604 19484 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 5080 6443 5132 6452
rect 5080 6409 5089 6443
rect 5089 6409 5123 6443
rect 5123 6409 5132 6443
rect 5080 6400 5132 6409
rect 6000 6400 6052 6452
rect 6920 6400 6972 6452
rect 9036 6443 9088 6452
rect 9036 6409 9045 6443
rect 9045 6409 9079 6443
rect 9079 6409 9088 6443
rect 9036 6400 9088 6409
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 9864 6400 9916 6452
rect 10232 6400 10284 6452
rect 6092 6264 6144 6316
rect 8300 6264 8352 6316
rect 5448 6239 5500 6248
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 5448 6196 5500 6205
rect 5540 6196 5592 6248
rect 7012 6196 7064 6248
rect 9128 6196 9180 6248
rect 7104 6103 7156 6112
rect 7104 6069 7113 6103
rect 7113 6069 7147 6103
rect 7147 6069 7156 6103
rect 11796 6400 11848 6452
rect 13176 6400 13228 6452
rect 15476 6400 15528 6452
rect 17408 6443 17460 6452
rect 17408 6409 17417 6443
rect 17417 6409 17451 6443
rect 17451 6409 17460 6443
rect 17408 6400 17460 6409
rect 18788 6400 18840 6452
rect 20996 6443 21048 6452
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 11244 6264 11296 6316
rect 12532 6264 12584 6316
rect 14280 6307 14332 6316
rect 14280 6273 14289 6307
rect 14289 6273 14323 6307
rect 14323 6273 14332 6307
rect 14280 6264 14332 6273
rect 14372 6264 14424 6316
rect 14740 6264 14792 6316
rect 15384 6264 15436 6316
rect 19800 6332 19852 6384
rect 24768 6375 24820 6384
rect 24768 6341 24777 6375
rect 24777 6341 24811 6375
rect 24811 6341 24820 6375
rect 24768 6332 24820 6341
rect 18880 6264 18932 6316
rect 19340 6264 19392 6316
rect 17776 6239 17828 6248
rect 11612 6128 11664 6180
rect 7104 6060 7156 6069
rect 9496 6060 9548 6112
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 17776 6205 17785 6239
rect 17785 6205 17819 6239
rect 17819 6205 17828 6239
rect 17776 6196 17828 6205
rect 19432 6196 19484 6248
rect 24584 6239 24636 6248
rect 24584 6205 24593 6239
rect 24593 6205 24627 6239
rect 24627 6205 24636 6239
rect 24584 6196 24636 6205
rect 17960 6128 18012 6180
rect 17776 6060 17828 6112
rect 19800 6171 19852 6180
rect 19800 6137 19809 6171
rect 19809 6137 19843 6171
rect 19843 6137 19852 6171
rect 19800 6128 19852 6137
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 5540 5856 5592 5908
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 9036 5856 9088 5908
rect 9220 5856 9272 5908
rect 10140 5856 10192 5908
rect 11152 5856 11204 5908
rect 12900 5856 12952 5908
rect 13176 5856 13228 5908
rect 14004 5899 14056 5908
rect 14004 5865 14013 5899
rect 14013 5865 14047 5899
rect 14047 5865 14056 5899
rect 14004 5856 14056 5865
rect 14832 5856 14884 5908
rect 16856 5899 16908 5908
rect 16856 5865 16865 5899
rect 16865 5865 16899 5899
rect 16899 5865 16908 5899
rect 16856 5856 16908 5865
rect 7104 5831 7156 5840
rect 7104 5797 7107 5831
rect 7107 5797 7141 5831
rect 7141 5797 7156 5831
rect 7104 5788 7156 5797
rect 6184 5720 6236 5772
rect 7564 5720 7616 5772
rect 9404 5788 9456 5840
rect 9864 5831 9916 5840
rect 9864 5797 9873 5831
rect 9873 5797 9907 5831
rect 9907 5797 9916 5831
rect 9864 5788 9916 5797
rect 12624 5831 12676 5840
rect 12624 5797 12633 5831
rect 12633 5797 12667 5831
rect 12667 5797 12676 5831
rect 12624 5788 12676 5797
rect 15292 5831 15344 5840
rect 15292 5797 15301 5831
rect 15301 5797 15335 5831
rect 15335 5797 15344 5831
rect 15292 5788 15344 5797
rect 17776 5831 17828 5840
rect 17776 5797 17785 5831
rect 17785 5797 17819 5831
rect 17819 5797 17828 5831
rect 17776 5788 17828 5797
rect 19248 5788 19300 5840
rect 20904 5788 20956 5840
rect 8668 5763 8720 5772
rect 8668 5729 8686 5763
rect 8686 5729 8720 5763
rect 8668 5720 8720 5729
rect 14556 5720 14608 5772
rect 15476 5763 15528 5772
rect 15476 5729 15485 5763
rect 15485 5729 15519 5763
rect 15519 5729 15528 5763
rect 15476 5720 15528 5729
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 9680 5584 9732 5636
rect 10968 5652 11020 5704
rect 13268 5652 13320 5704
rect 13636 5695 13688 5704
rect 13636 5661 13645 5695
rect 13645 5661 13679 5695
rect 13679 5661 13688 5695
rect 13636 5652 13688 5661
rect 16764 5652 16816 5704
rect 19340 5652 19392 5704
rect 19524 5695 19576 5704
rect 19524 5661 19533 5695
rect 19533 5661 19567 5695
rect 19567 5661 19576 5695
rect 19524 5652 19576 5661
rect 11060 5584 11112 5636
rect 11796 5584 11848 5636
rect 13084 5584 13136 5636
rect 14280 5584 14332 5636
rect 17776 5516 17828 5568
rect 18696 5516 18748 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 6184 5355 6236 5364
rect 6184 5321 6193 5355
rect 6193 5321 6227 5355
rect 6227 5321 6236 5355
rect 6184 5312 6236 5321
rect 7104 5355 7156 5364
rect 7104 5321 7113 5355
rect 7113 5321 7147 5355
rect 7147 5321 7156 5355
rect 7104 5312 7156 5321
rect 8668 5355 8720 5364
rect 8668 5321 8677 5355
rect 8677 5321 8711 5355
rect 8711 5321 8720 5355
rect 8668 5312 8720 5321
rect 9864 5312 9916 5364
rect 11796 5355 11848 5364
rect 11796 5321 11805 5355
rect 11805 5321 11839 5355
rect 11839 5321 11848 5355
rect 11796 5312 11848 5321
rect 13820 5355 13872 5364
rect 13820 5321 13829 5355
rect 13829 5321 13863 5355
rect 13863 5321 13872 5355
rect 13820 5312 13872 5321
rect 14556 5312 14608 5364
rect 15476 5355 15528 5364
rect 15476 5321 15485 5355
rect 15485 5321 15519 5355
rect 15519 5321 15528 5355
rect 15476 5312 15528 5321
rect 17776 5312 17828 5364
rect 19248 5355 19300 5364
rect 19248 5321 19257 5355
rect 19257 5321 19291 5355
rect 19291 5321 19300 5355
rect 19248 5312 19300 5321
rect 19340 5312 19392 5364
rect 23480 5312 23532 5364
rect 9404 5244 9456 5296
rect 9588 5287 9640 5296
rect 9588 5253 9597 5287
rect 9597 5253 9631 5287
rect 9631 5253 9640 5287
rect 9588 5244 9640 5253
rect 12624 5244 12676 5296
rect 13084 5287 13136 5296
rect 13084 5253 13093 5287
rect 13093 5253 13127 5287
rect 13127 5253 13136 5287
rect 13084 5244 13136 5253
rect 14004 5244 14056 5296
rect 9220 5176 9272 5228
rect 10968 5176 11020 5228
rect 12532 5219 12584 5228
rect 12532 5185 12541 5219
rect 12541 5185 12575 5219
rect 12575 5185 12584 5219
rect 12532 5176 12584 5185
rect 14372 5219 14424 5228
rect 14372 5185 14381 5219
rect 14381 5185 14415 5219
rect 14415 5185 14424 5219
rect 14372 5176 14424 5185
rect 17132 5176 17184 5228
rect 17684 5176 17736 5228
rect 19432 5176 19484 5228
rect 6368 5040 6420 5092
rect 7564 5083 7616 5092
rect 7564 5049 7573 5083
rect 7573 5049 7607 5083
rect 7607 5049 7616 5083
rect 8116 5083 8168 5092
rect 7564 5040 7616 5049
rect 8116 5049 8125 5083
rect 8125 5049 8159 5083
rect 8159 5049 8168 5083
rect 8116 5040 8168 5049
rect 9128 5083 9180 5092
rect 9128 5049 9137 5083
rect 9137 5049 9171 5083
rect 9171 5049 9180 5083
rect 9128 5040 9180 5049
rect 11060 5040 11112 5092
rect 11520 5083 11572 5092
rect 11520 5049 11529 5083
rect 11529 5049 11563 5083
rect 11563 5049 11572 5083
rect 11520 5040 11572 5049
rect 11980 5040 12032 5092
rect 12532 5040 12584 5092
rect 12624 5083 12676 5092
rect 12624 5049 12633 5083
rect 12633 5049 12667 5083
rect 12667 5049 12676 5083
rect 12624 5040 12676 5049
rect 10876 4972 10928 5024
rect 11336 4972 11388 5024
rect 13820 4972 13872 5024
rect 15752 4972 15804 5024
rect 16764 5015 16816 5024
rect 16764 4981 16773 5015
rect 16773 4981 16807 5015
rect 16807 4981 16816 5015
rect 16764 4972 16816 4981
rect 25136 5015 25188 5024
rect 25136 4981 25145 5015
rect 25145 4981 25179 5015
rect 25179 4981 25188 5015
rect 25136 4972 25188 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 9128 4768 9180 4820
rect 9772 4768 9824 4820
rect 12900 4768 12952 4820
rect 17868 4768 17920 4820
rect 24768 4811 24820 4820
rect 24768 4777 24777 4811
rect 24777 4777 24811 4811
rect 24811 4777 24820 4811
rect 24768 4768 24820 4777
rect 7564 4743 7616 4752
rect 7564 4709 7573 4743
rect 7573 4709 7607 4743
rect 7607 4709 7616 4743
rect 7564 4700 7616 4709
rect 8208 4700 8260 4752
rect 10876 4743 10928 4752
rect 10876 4709 10885 4743
rect 10885 4709 10919 4743
rect 10919 4709 10928 4743
rect 10876 4700 10928 4709
rect 11520 4700 11572 4752
rect 12072 4700 12124 4752
rect 12348 4700 12400 4752
rect 13084 4700 13136 4752
rect 9864 4632 9916 4684
rect 10600 4632 10652 4684
rect 14188 4632 14240 4684
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 17592 4632 17644 4684
rect 24216 4632 24268 4684
rect 7196 4564 7248 4616
rect 10140 4564 10192 4616
rect 12348 4607 12400 4616
rect 12348 4573 12357 4607
rect 12357 4573 12391 4607
rect 12391 4573 12400 4607
rect 12348 4564 12400 4573
rect 9680 4428 9732 4480
rect 15936 4471 15988 4480
rect 15936 4437 15945 4471
rect 15945 4437 15979 4471
rect 15979 4437 15988 4471
rect 15936 4428 15988 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 7564 4224 7616 4276
rect 9864 4267 9916 4276
rect 9864 4233 9873 4267
rect 9873 4233 9907 4267
rect 9907 4233 9916 4267
rect 9864 4224 9916 4233
rect 10876 4224 10928 4276
rect 12348 4224 12400 4276
rect 14188 4224 14240 4276
rect 15752 4267 15804 4276
rect 7196 4156 7248 4208
rect 8116 4088 8168 4140
rect 9220 4156 9272 4208
rect 8576 4088 8628 4140
rect 8944 4131 8996 4140
rect 7380 3995 7432 4004
rect 7380 3961 7389 3995
rect 7389 3961 7423 3995
rect 7423 3961 7432 3995
rect 7380 3952 7432 3961
rect 8944 4097 8953 4131
rect 8953 4097 8987 4131
rect 8987 4097 8996 4131
rect 8944 4088 8996 4097
rect 9588 4088 9640 4140
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 12532 4088 12584 4140
rect 14372 4156 14424 4208
rect 15752 4233 15761 4267
rect 15761 4233 15795 4267
rect 15795 4233 15804 4267
rect 15752 4224 15804 4233
rect 17592 4224 17644 4276
rect 24216 4224 24268 4276
rect 16120 4156 16172 4208
rect 12072 4020 12124 4072
rect 10048 3952 10100 4004
rect 10876 3995 10928 4004
rect 10876 3961 10885 3995
rect 10885 3961 10919 3995
rect 10919 3961 10928 3995
rect 10876 3952 10928 3961
rect 10968 3995 11020 4004
rect 10968 3961 10977 3995
rect 10977 3961 11011 3995
rect 11011 3961 11020 3995
rect 12532 3995 12584 4004
rect 10968 3952 11020 3961
rect 12532 3961 12541 3995
rect 12541 3961 12575 3995
rect 12575 3961 12584 3995
rect 12532 3952 12584 3961
rect 10140 3884 10192 3936
rect 12440 3884 12492 3936
rect 19432 4020 19484 4072
rect 14740 3884 14792 3936
rect 14924 3927 14976 3936
rect 14924 3893 14933 3927
rect 14933 3893 14967 3927
rect 14967 3893 14976 3927
rect 14924 3884 14976 3893
rect 20444 3927 20496 3936
rect 20444 3893 20453 3927
rect 20453 3893 20487 3927
rect 20487 3893 20496 3927
rect 20444 3884 20496 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2688 3680 2740 3732
rect 5448 3680 5500 3732
rect 7380 3680 7432 3732
rect 8944 3723 8996 3732
rect 8944 3689 8953 3723
rect 8953 3689 8987 3723
rect 8987 3689 8996 3723
rect 8944 3680 8996 3689
rect 10876 3680 10928 3732
rect 11980 3680 12032 3732
rect 12440 3723 12492 3732
rect 12440 3689 12449 3723
rect 12449 3689 12483 3723
rect 12483 3689 12492 3723
rect 12440 3680 12492 3689
rect 7748 3612 7800 3664
rect 8116 3655 8168 3664
rect 8116 3621 8125 3655
rect 8125 3621 8159 3655
rect 8159 3621 8168 3655
rect 8116 3612 8168 3621
rect 9496 3612 9548 3664
rect 9772 3655 9824 3664
rect 9772 3621 9781 3655
rect 9781 3621 9815 3655
rect 9815 3621 9824 3655
rect 9772 3612 9824 3621
rect 9864 3655 9916 3664
rect 9864 3621 9873 3655
rect 9873 3621 9907 3655
rect 9907 3621 9916 3655
rect 9864 3612 9916 3621
rect 12532 3612 12584 3664
rect 2504 3544 2556 3596
rect 5448 3587 5500 3596
rect 5448 3553 5466 3587
rect 5466 3553 5500 3587
rect 5448 3544 5500 3553
rect 6368 3587 6420 3596
rect 6368 3553 6412 3587
rect 6412 3553 6420 3587
rect 6368 3544 6420 3553
rect 10968 3544 11020 3596
rect 11796 3587 11848 3596
rect 11796 3553 11814 3587
rect 11814 3553 11848 3587
rect 11796 3544 11848 3553
rect 21272 3544 21324 3596
rect 22100 3544 22152 3596
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 9220 3476 9272 3528
rect 21824 3451 21876 3460
rect 21824 3417 21833 3451
rect 21833 3417 21867 3451
rect 21867 3417 21876 3451
rect 21824 3408 21876 3417
rect 12900 3340 12952 3392
rect 15384 3340 15436 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 7472 3136 7524 3188
rect 9404 3136 9456 3188
rect 7748 3111 7800 3120
rect 7748 3077 7757 3111
rect 7757 3077 7791 3111
rect 7791 3077 7800 3111
rect 7748 3068 7800 3077
rect 6644 2932 6696 2984
rect 9772 3136 9824 3188
rect 11796 3179 11848 3188
rect 11796 3145 11805 3179
rect 11805 3145 11839 3179
rect 11839 3145 11848 3179
rect 11796 3136 11848 3145
rect 21732 3179 21784 3188
rect 21732 3145 21741 3179
rect 21741 3145 21775 3179
rect 21775 3145 21784 3179
rect 21732 3136 21784 3145
rect 22100 3179 22152 3188
rect 22100 3145 22109 3179
rect 22109 3145 22143 3179
rect 22143 3145 22152 3179
rect 22100 3136 22152 3145
rect 9864 3068 9916 3120
rect 20076 3068 20128 3120
rect 12716 2932 12768 2984
rect 17960 2932 18012 2984
rect 21732 2932 21784 2984
rect 24308 2975 24360 2984
rect 24308 2941 24317 2975
rect 24317 2941 24351 2975
rect 24351 2941 24360 2975
rect 24308 2932 24360 2941
rect 10968 2864 11020 2916
rect 13728 2864 13780 2916
rect 2504 2796 2556 2848
rect 5448 2839 5500 2848
rect 5448 2805 5457 2839
rect 5457 2805 5491 2839
rect 5491 2805 5500 2839
rect 5448 2796 5500 2805
rect 6368 2839 6420 2848
rect 6368 2805 6377 2839
rect 6377 2805 6411 2839
rect 6411 2805 6420 2839
rect 6368 2796 6420 2805
rect 23204 2796 23256 2848
rect 24492 2839 24544 2848
rect 24492 2805 24501 2839
rect 24501 2805 24535 2839
rect 24535 2805 24544 2839
rect 24492 2796 24544 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1584 2592 1636 2644
rect 4620 2592 4672 2644
rect 7380 2592 7432 2644
rect 9956 2592 10008 2644
rect 10784 2592 10836 2644
rect 16764 2592 16816 2644
rect 18972 2635 19024 2644
rect 18972 2601 18981 2635
rect 18981 2601 19015 2635
rect 19015 2601 19024 2635
rect 18972 2592 19024 2601
rect 1400 2499 1452 2508
rect 1400 2465 1444 2499
rect 1444 2465 1452 2499
rect 1400 2456 1452 2465
rect 4620 2388 4672 2440
rect 9864 2499 9916 2508
rect 9864 2465 9908 2499
rect 9908 2465 9916 2499
rect 9864 2456 9916 2465
rect 7656 2252 7708 2304
rect 17040 2456 17092 2508
rect 20260 2592 20312 2644
rect 21916 2635 21968 2644
rect 21916 2601 21925 2635
rect 21925 2601 21959 2635
rect 21959 2601 21968 2635
rect 21916 2592 21968 2601
rect 21732 2499 21784 2508
rect 21732 2465 21741 2499
rect 21741 2465 21775 2499
rect 21775 2465 21784 2499
rect 21732 2456 21784 2465
rect 22836 2499 22888 2508
rect 22836 2465 22845 2499
rect 22845 2465 22879 2499
rect 22879 2465 22888 2499
rect 22836 2456 22888 2465
rect 23664 2456 23716 2508
rect 19064 2320 19116 2372
rect 21180 2320 21232 2372
rect 25320 2320 25372 2372
rect 11796 2252 11848 2304
rect 17040 2295 17092 2304
rect 17040 2261 17049 2295
rect 17049 2261 17083 2295
rect 17083 2261 17092 2295
rect 17040 2252 17092 2261
rect 24768 2295 24820 2304
rect 24768 2261 24777 2295
rect 24777 2261 24811 2295
rect 24811 2261 24820 2295
rect 24768 2252 24820 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 478 27520 534 28000
rect 1490 27520 1546 28000
rect 2502 27520 2558 28000
rect 3514 27520 3570 28000
rect 4618 27520 4674 28000
rect 5630 27520 5686 28000
rect 6642 27520 6698 28000
rect 7654 27520 7710 28000
rect 8758 27520 8814 28000
rect 9770 27520 9826 28000
rect 10782 27520 10838 28000
rect 11794 27520 11850 28000
rect 12898 27520 12954 28000
rect 13910 27520 13966 28000
rect 14922 27520 14978 28000
rect 15934 27520 15990 28000
rect 17038 27520 17094 28000
rect 18050 27520 18106 28000
rect 19062 27520 19118 28000
rect 20074 27520 20130 28000
rect 21178 27520 21234 28000
rect 22190 27520 22246 28000
rect 23202 27520 23258 28000
rect 24214 27520 24270 28000
rect 25318 27520 25374 28000
rect 26330 27520 26386 28000
rect 27342 27520 27398 28000
rect 492 23662 520 27520
rect 1504 24274 1532 27520
rect 1492 24268 1544 24274
rect 1492 24210 1544 24216
rect 1504 23866 1532 24210
rect 1492 23860 1544 23866
rect 1492 23802 1544 23808
rect 2516 23662 2544 27520
rect 2686 24168 2742 24177
rect 2686 24103 2688 24112
rect 2740 24103 2742 24112
rect 2688 24074 2740 24080
rect 3528 23662 3556 27520
rect 4066 26480 4122 26489
rect 4066 26415 4122 26424
rect 4080 26314 4108 26415
rect 4068 26308 4120 26314
rect 4068 26250 4120 26256
rect 4632 24274 4660 27520
rect 5644 25140 5672 27520
rect 6184 26308 6236 26314
rect 6184 26250 6236 26256
rect 5552 25112 5672 25140
rect 5552 24818 5580 25112
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 5448 24608 5500 24614
rect 5448 24550 5500 24556
rect 5460 24313 5488 24550
rect 5446 24304 5502 24313
rect 4620 24268 4672 24274
rect 5446 24239 5502 24248
rect 4620 24210 4672 24216
rect 4632 23866 4660 24210
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 5540 24064 5592 24070
rect 5540 24006 5592 24012
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 5276 23730 5304 24006
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 480 23656 532 23662
rect 480 23598 532 23604
rect 2504 23656 2556 23662
rect 3516 23656 3568 23662
rect 2504 23598 2556 23604
rect 2686 23624 2742 23633
rect 3516 23598 3568 23604
rect 2686 23559 2742 23568
rect 5356 23588 5408 23594
rect 2700 23526 2728 23559
rect 5356 23530 5408 23536
rect 2688 23520 2740 23526
rect 5368 23497 5396 23530
rect 2688 23462 2740 23468
rect 5354 23488 5410 23497
rect 5354 23423 5410 23432
rect 3422 23352 3478 23361
rect 5368 23322 5396 23423
rect 5552 23322 5580 24006
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5908 23588 5960 23594
rect 5908 23530 5960 23536
rect 3422 23287 3478 23296
rect 5356 23316 5408 23322
rect 3436 14929 3464 23287
rect 5356 23258 5408 23264
rect 5540 23316 5592 23322
rect 5540 23258 5592 23264
rect 5552 22778 5580 23258
rect 5920 23118 5948 23530
rect 6000 23248 6052 23254
rect 6000 23190 6052 23196
rect 5908 23112 5960 23118
rect 5908 23054 5960 23060
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 6012 22438 6040 23190
rect 6000 22432 6052 22438
rect 5078 22400 5134 22409
rect 6000 22374 6052 22380
rect 5078 22335 5134 22344
rect 5092 22234 5120 22335
rect 5080 22228 5132 22234
rect 5080 22170 5132 22176
rect 6196 22166 6224 26250
rect 6552 24336 6604 24342
rect 6552 24278 6604 24284
rect 6460 24200 6512 24206
rect 6460 24142 6512 24148
rect 6472 23526 6500 24142
rect 6564 23798 6592 24278
rect 6656 24138 6684 27520
rect 7668 24698 7696 27520
rect 8772 27418 8800 27520
rect 8772 27390 8892 27418
rect 8574 24848 8630 24857
rect 8574 24783 8576 24792
rect 8628 24783 8630 24792
rect 8576 24754 8628 24760
rect 7668 24670 7788 24698
rect 6828 24608 6880 24614
rect 6828 24550 6880 24556
rect 7656 24608 7708 24614
rect 7656 24550 7708 24556
rect 6736 24200 6788 24206
rect 6736 24142 6788 24148
rect 6644 24132 6696 24138
rect 6644 24074 6696 24080
rect 6656 23866 6684 24074
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 6552 23792 6604 23798
rect 6552 23734 6604 23740
rect 6460 23520 6512 23526
rect 6460 23462 6512 23468
rect 6472 23322 6500 23462
rect 6460 23316 6512 23322
rect 6460 23258 6512 23264
rect 6564 22506 6592 23734
rect 6748 23100 6776 24142
rect 6840 23202 6868 24550
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7576 23594 7604 24006
rect 7564 23588 7616 23594
rect 7564 23530 7616 23536
rect 7104 23520 7156 23526
rect 7102 23488 7104 23497
rect 7156 23488 7158 23497
rect 7102 23423 7158 23432
rect 6840 23174 6960 23202
rect 6932 23118 6960 23174
rect 6828 23112 6880 23118
rect 6748 23072 6828 23100
rect 6828 23054 6880 23060
rect 6920 23112 6972 23118
rect 6920 23054 6972 23060
rect 6552 22500 6604 22506
rect 6552 22442 6604 22448
rect 6184 22160 6236 22166
rect 6184 22102 6236 22108
rect 5080 22092 5132 22098
rect 5080 22034 5132 22040
rect 5448 22092 5500 22098
rect 5448 22034 5500 22040
rect 5092 21350 5120 22034
rect 4528 21344 4580 21350
rect 4528 21286 4580 21292
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 4540 20806 4568 21286
rect 5460 20806 5488 22034
rect 6000 21888 6052 21894
rect 5998 21856 6000 21865
rect 6052 21856 6054 21865
rect 5622 21788 5918 21808
rect 5998 21791 6054 21800
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6012 21554 6040 21791
rect 6196 21690 6224 22102
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6000 21548 6052 21554
rect 6000 21490 6052 21496
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5644 21010 5672 21422
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6196 21049 6224 21286
rect 6380 21078 6408 21966
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6368 21072 6420 21078
rect 6182 21040 6238 21049
rect 5632 21004 5684 21010
rect 6368 21014 6420 21020
rect 6182 20975 6184 20984
rect 5632 20946 5684 20952
rect 6236 20975 6238 20984
rect 6184 20946 6236 20952
rect 5644 20890 5672 20946
rect 5552 20862 5672 20890
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5460 20398 5488 20742
rect 5356 20392 5408 20398
rect 5356 20334 5408 20340
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 5092 19174 5120 19858
rect 5368 19242 5396 20334
rect 5552 20058 5580 20862
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6196 20602 6224 20946
rect 6184 20596 6236 20602
rect 6184 20538 6236 20544
rect 5724 20392 5776 20398
rect 5722 20360 5724 20369
rect 5776 20360 5778 20369
rect 5722 20295 5778 20304
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 5552 19310 5580 19994
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6012 19378 6040 19654
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 5540 19304 5592 19310
rect 5724 19304 5776 19310
rect 5540 19246 5592 19252
rect 5722 19272 5724 19281
rect 5776 19272 5778 19281
rect 5356 19236 5408 19242
rect 5356 19178 5408 19184
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 5092 18873 5120 19110
rect 5078 18864 5134 18873
rect 5552 18834 5580 19246
rect 5722 19207 5778 19216
rect 5078 18799 5134 18808
rect 5540 18828 5592 18834
rect 5540 18770 5592 18776
rect 5552 18426 5580 18770
rect 5736 18698 5764 19207
rect 5724 18692 5776 18698
rect 5724 18634 5776 18640
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5184 17746 5212 18362
rect 5540 18216 5592 18222
rect 5460 18164 5540 18170
rect 5460 18158 5592 18164
rect 5460 18142 5580 18158
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5184 17338 5212 17682
rect 5368 17649 5396 17682
rect 5460 17678 5488 18142
rect 5448 17672 5500 17678
rect 5354 17640 5410 17649
rect 5448 17614 5500 17620
rect 5354 17575 5410 17584
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 4066 17096 4122 17105
rect 4066 17031 4122 17040
rect 3422 14920 3478 14929
rect 3422 14855 3478 14864
rect 4080 14226 4108 17031
rect 5184 16794 5212 17274
rect 5368 17270 5396 17575
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5356 17264 5408 17270
rect 5356 17206 5408 17212
rect 6196 16946 6224 20538
rect 6564 19990 6592 21490
rect 6840 21026 6868 23054
rect 6932 22778 6960 23054
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 7024 21146 7052 21422
rect 7012 21140 7064 21146
rect 7012 21082 7064 21088
rect 6840 20998 6960 21026
rect 6840 20602 6868 20998
rect 6932 20942 6960 20998
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6552 19984 6604 19990
rect 6552 19926 6604 19932
rect 6564 19514 6592 19926
rect 6552 19508 6604 19514
rect 6552 19450 6604 19456
rect 6564 19242 6592 19450
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6552 19236 6604 19242
rect 6552 19178 6604 19184
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 6368 18624 6420 18630
rect 6368 18566 6420 18572
rect 6274 17776 6330 17785
rect 6274 17711 6330 17720
rect 6288 17338 6316 17711
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6196 16918 6316 16946
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 4356 16697 4384 16730
rect 4342 16688 4398 16697
rect 4252 16652 4304 16658
rect 6196 16658 6224 16730
rect 4342 16623 4398 16632
rect 5172 16652 5224 16658
rect 4252 16594 4304 16600
rect 6184 16652 6236 16658
rect 5224 16612 5304 16640
rect 5172 16594 5224 16600
rect 4264 15910 4292 16594
rect 5276 16046 5304 16612
rect 6184 16594 6236 16600
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6196 16250 6224 16594
rect 6288 16289 6316 16918
rect 6274 16280 6330 16289
rect 6184 16244 6236 16250
rect 6274 16215 6330 16224
rect 6184 16186 6236 16192
rect 5264 16040 5316 16046
rect 5262 16008 5264 16017
rect 5316 16008 5318 16017
rect 5262 15943 5318 15952
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 4264 15065 4292 15846
rect 5644 15706 5672 15846
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 4250 15056 4306 15065
rect 4250 14991 4306 15000
rect 5460 14822 5488 15438
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5552 15026 5580 15370
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5552 14929 5580 14962
rect 5538 14920 5594 14929
rect 5538 14855 5594 14864
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 4080 14198 4200 14226
rect 4172 14074 4200 14198
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4066 13968 4122 13977
rect 4066 13903 4122 13912
rect 2502 13696 2558 13705
rect 2502 13631 2558 13640
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2056 11694 2084 12174
rect 2516 12170 2544 13631
rect 4080 13410 4108 13903
rect 4172 13870 4200 14010
rect 5368 13870 5396 14418
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4356 13705 4384 13738
rect 4342 13696 4398 13705
rect 4342 13631 4398 13640
rect 4160 13456 4212 13462
rect 4080 13404 4160 13410
rect 4080 13398 4212 13404
rect 4080 13382 4200 13398
rect 4080 12968 4108 13382
rect 4356 13326 4384 13631
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4160 12980 4212 12986
rect 4080 12940 4160 12968
rect 4160 12922 4212 12928
rect 4436 12776 4488 12782
rect 2870 12744 2926 12753
rect 4436 12718 4488 12724
rect 2870 12679 2872 12688
rect 2924 12679 2926 12688
rect 2872 12650 2924 12656
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 4068 12640 4120 12646
rect 4120 12600 4200 12628
rect 4068 12582 4120 12588
rect 2608 12209 2636 12582
rect 3620 12345 3648 12582
rect 4172 12442 4200 12600
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 3606 12336 3662 12345
rect 2688 12300 2740 12306
rect 3606 12271 3662 12280
rect 2688 12242 2740 12248
rect 2594 12200 2650 12209
rect 2504 12164 2556 12170
rect 2594 12135 2650 12144
rect 2504 12106 2556 12112
rect 2516 11898 2544 12106
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 2226 11656 2282 11665
rect 2056 11354 2084 11630
rect 2226 11591 2282 11600
rect 2240 11558 2268 11591
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2240 11218 2268 11494
rect 2608 11218 2636 12135
rect 2700 11898 2728 12242
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4172 11898 4200 12174
rect 4448 11898 4476 12718
rect 4632 12306 4660 13330
rect 4908 12306 4936 13806
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5276 12986 5304 13262
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 5184 12306 5212 12650
rect 4620 12300 4672 12306
rect 4896 12300 4948 12306
rect 4620 12242 4672 12248
rect 4816 12260 4896 12288
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4632 11694 4660 12242
rect 4816 11830 4844 12260
rect 4896 12242 4948 12248
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4816 11626 4844 11766
rect 5368 11762 5396 13806
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 2056 10810 2084 11086
rect 2240 10810 2268 11154
rect 2608 11098 2636 11154
rect 2608 11070 2820 11098
rect 2792 10810 2820 11070
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2148 9722 2176 10066
rect 2504 9988 2556 9994
rect 2504 9930 2556 9936
rect 2516 9722 2544 9930
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2608 9382 2636 10066
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 8634 2636 9318
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2608 7721 2636 8570
rect 2594 7712 2650 7721
rect 2594 7647 2650 7656
rect 2700 7528 2728 10406
rect 2700 7500 2820 7528
rect 2792 7274 2820 7500
rect 2780 7268 2832 7274
rect 2780 7210 2832 7216
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2700 3641 2728 3674
rect 2686 3632 2742 3641
rect 2504 3596 2556 3602
rect 2686 3567 2742 3576
rect 2504 3538 2556 3544
rect 2516 2854 2544 3538
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 1582 2680 1638 2689
rect 1582 2615 1584 2624
rect 1636 2615 1638 2624
rect 1584 2586 1636 2592
rect 1490 2544 1546 2553
rect 1400 2508 1452 2514
rect 1490 2479 1546 2488
rect 1400 2450 1452 2456
rect 1412 1873 1440 2450
rect 478 1864 534 1873
rect 478 1799 534 1808
rect 1398 1864 1454 1873
rect 1398 1799 1454 1808
rect 492 480 520 1799
rect 1504 480 1532 2479
rect 2516 480 2544 2790
rect 2884 1601 2912 11494
rect 4816 11354 4844 11562
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 5460 11286 5488 14758
rect 6012 14278 6040 15506
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 6288 14226 6316 16215
rect 6380 15858 6408 18566
rect 6472 18290 6500 18770
rect 6564 18426 6592 19178
rect 6840 18902 6868 19246
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6472 18193 6500 18226
rect 6458 18184 6514 18193
rect 6564 18154 6592 18362
rect 6932 18222 6960 18566
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6458 18119 6514 18128
rect 6552 18148 6604 18154
rect 6552 18090 6604 18096
rect 6564 17814 6592 18090
rect 7116 17882 7144 23423
rect 7288 23248 7340 23254
rect 7288 23190 7340 23196
rect 7300 22438 7328 23190
rect 7472 22500 7524 22506
rect 7472 22442 7524 22448
rect 7288 22432 7340 22438
rect 7288 22374 7340 22380
rect 7300 21978 7328 22374
rect 7484 22234 7512 22442
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7208 21950 7328 21978
rect 7208 20058 7236 21950
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 7300 21078 7328 21830
rect 7288 21072 7340 21078
rect 7288 21014 7340 21020
rect 7300 20602 7328 21014
rect 7288 20596 7340 20602
rect 7288 20538 7340 20544
rect 7286 20224 7342 20233
rect 7286 20159 7342 20168
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 6552 17808 6604 17814
rect 6604 17756 6684 17762
rect 6552 17750 6684 17756
rect 6564 17734 6684 17750
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6550 17640 6606 17649
rect 6472 17066 6500 17614
rect 6550 17575 6606 17584
rect 6460 17060 6512 17066
rect 6460 17002 6512 17008
rect 6472 16794 6500 17002
rect 6460 16788 6512 16794
rect 6460 16730 6512 16736
rect 6458 15872 6514 15881
rect 6380 15830 6458 15858
rect 6458 15807 6514 15816
rect 6288 14198 6408 14226
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5552 12306 5580 13262
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6196 12374 6224 12582
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6196 11898 6224 12310
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10810 3188 11086
rect 3330 10840 3386 10849
rect 3148 10804 3200 10810
rect 3330 10775 3386 10784
rect 3148 10746 3200 10752
rect 3160 10606 3188 10746
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3146 10160 3202 10169
rect 3146 10095 3148 10104
rect 3200 10095 3202 10104
rect 3148 10066 3200 10072
rect 3344 9586 3372 10775
rect 3700 10736 3752 10742
rect 3698 10704 3700 10713
rect 3752 10704 3754 10713
rect 3698 10639 3754 10648
rect 4908 10470 4936 11154
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 4068 10464 4120 10470
rect 4066 10432 4068 10441
rect 4896 10464 4948 10470
rect 4120 10432 4122 10441
rect 4896 10406 4948 10412
rect 4066 10367 4122 10376
rect 4908 10130 4936 10406
rect 5092 10266 5120 11018
rect 5276 10554 5304 11154
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5998 10704 6054 10713
rect 5998 10639 6054 10648
rect 5540 10600 5592 10606
rect 5276 10548 5540 10554
rect 5276 10542 5592 10548
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5276 10526 5580 10542
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 4908 9382 4936 10066
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 5000 9586 5028 9930
rect 5092 9722 5120 10202
rect 5184 10062 5212 10474
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 5184 9602 5212 9998
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5092 9574 5212 9602
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4632 8634 4660 8978
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4908 8430 4936 9318
rect 5000 9178 5028 9522
rect 5092 9518 5120 9574
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5000 8566 5028 9114
rect 5172 9036 5224 9042
rect 5276 9024 5304 10526
rect 5538 10432 5594 10441
rect 5538 10367 5594 10376
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5368 9518 5396 10066
rect 5552 9586 5580 10367
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5368 9110 5396 9454
rect 5446 9344 5502 9353
rect 5446 9279 5502 9288
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5224 8996 5304 9024
rect 5172 8978 5224 8984
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 4160 8424 4212 8430
rect 4080 8384 4160 8412
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3712 7002 3740 7278
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3896 6905 3924 7142
rect 3882 6896 3938 6905
rect 3882 6831 3938 6840
rect 4080 4593 4108 8384
rect 4160 8366 4212 8372
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 5170 7984 5226 7993
rect 5170 7919 5172 7928
rect 5224 7919 5226 7928
rect 5172 7890 5224 7896
rect 5184 7546 5212 7890
rect 5460 7886 5488 9279
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6012 8673 6040 10639
rect 6288 9994 6316 14010
rect 6380 13938 6408 14198
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6380 11898 6408 12242
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6472 11354 6500 15807
rect 6564 14482 6592 17575
rect 6656 17338 6684 17734
rect 7116 17338 7144 17818
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6564 14074 6592 14418
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6564 12186 6592 13874
rect 6656 13705 6684 14758
rect 6642 13696 6698 13705
rect 6642 13631 6698 13640
rect 6564 12158 6684 12186
rect 6552 12096 6604 12102
rect 6550 12064 6552 12073
rect 6604 12064 6606 12073
rect 6550 11999 6606 12008
rect 6460 11348 6512 11354
rect 6380 11308 6460 11336
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 5998 8664 6054 8673
rect 5998 8599 6054 8608
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5446 7440 5502 7449
rect 5446 7375 5502 7384
rect 5460 7342 5488 7375
rect 5552 7342 5580 7890
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5092 6934 5120 7278
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 5092 6458 5120 6870
rect 5552 6866 5580 7278
rect 6012 6866 6040 8599
rect 6104 8498 6132 8978
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6288 7993 6316 9930
rect 6274 7984 6330 7993
rect 6274 7919 6330 7928
rect 6380 7449 6408 11308
rect 6460 11290 6512 11296
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6472 10198 6500 11154
rect 6656 10713 6684 12158
rect 6642 10704 6698 10713
rect 6642 10639 6698 10648
rect 6644 10464 6696 10470
rect 6642 10432 6644 10441
rect 6696 10432 6698 10441
rect 6642 10367 6698 10376
rect 6748 10198 6776 17070
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 7024 14550 7052 15438
rect 7116 15094 7144 15642
rect 7104 15088 7156 15094
rect 7104 15030 7156 15036
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 7116 14482 7144 15030
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 6828 14272 6880 14278
rect 6880 14220 6960 14226
rect 6828 14214 6960 14220
rect 6840 14198 6960 14214
rect 6932 12918 6960 14198
rect 7116 14074 7144 14418
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7300 13394 7328 20159
rect 7484 18970 7512 22170
rect 7576 22030 7604 23530
rect 7668 22642 7696 24550
rect 7760 23594 7788 24670
rect 8116 24336 8168 24342
rect 8116 24278 8168 24284
rect 8484 24336 8536 24342
rect 8484 24278 8536 24284
rect 8128 23866 8156 24278
rect 8496 23905 8524 24278
rect 8482 23896 8538 23905
rect 8116 23860 8168 23866
rect 8482 23831 8538 23840
rect 8116 23802 8168 23808
rect 8496 23798 8524 23831
rect 8484 23792 8536 23798
rect 8484 23734 8536 23740
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7748 23588 7800 23594
rect 7748 23530 7800 23536
rect 7852 23254 7880 23666
rect 7840 23248 7892 23254
rect 7840 23190 7892 23196
rect 7852 22642 7880 23190
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7668 22166 7696 22578
rect 7852 22234 7880 22578
rect 7840 22228 7892 22234
rect 7840 22170 7892 22176
rect 7656 22160 7708 22166
rect 7656 22102 7708 22108
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 8668 22092 8720 22098
rect 8668 22034 8720 22040
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 8128 21978 8156 22034
rect 8128 21950 8248 21978
rect 8220 21350 8248 21950
rect 8680 21554 8708 22034
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8668 21412 8720 21418
rect 8668 21354 8720 21360
rect 8208 21344 8260 21350
rect 8206 21312 8208 21321
rect 8260 21312 8262 21321
rect 8206 21247 8262 21256
rect 8680 21146 8708 21354
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8208 21072 8260 21078
rect 8208 21014 8260 21020
rect 8220 20534 8248 21014
rect 8208 20528 8260 20534
rect 8208 20470 8260 20476
rect 8864 20482 8892 27390
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9128 24676 9180 24682
rect 9128 24618 9180 24624
rect 9220 24676 9272 24682
rect 9220 24618 9272 24624
rect 9140 24410 9168 24618
rect 9128 24404 9180 24410
rect 9128 24346 9180 24352
rect 9140 23866 9168 24346
rect 9232 24342 9260 24618
rect 9220 24336 9272 24342
rect 9220 24278 9272 24284
rect 9692 24177 9720 25230
rect 9784 24834 9812 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10140 25288 10192 25294
rect 10140 25230 10192 25236
rect 9784 24806 10088 24834
rect 10152 24818 10180 25230
rect 10692 25152 10744 25158
rect 10692 25094 10744 25100
rect 9956 24744 10008 24750
rect 9956 24686 10008 24692
rect 9968 24274 9996 24686
rect 9956 24268 10008 24274
rect 9956 24210 10008 24216
rect 9678 24168 9734 24177
rect 9678 24103 9734 24112
rect 9862 24168 9918 24177
rect 9862 24103 9864 24112
rect 9916 24103 9918 24112
rect 9864 24074 9916 24080
rect 9968 23866 9996 24210
rect 9128 23860 9180 23866
rect 9128 23802 9180 23808
rect 9956 23860 10008 23866
rect 9956 23802 10008 23808
rect 9956 22500 10008 22506
rect 9956 22442 10008 22448
rect 9128 22432 9180 22438
rect 9126 22400 9128 22409
rect 9180 22400 9182 22409
rect 9126 22335 9182 22344
rect 9968 22166 9996 22442
rect 9956 22160 10008 22166
rect 9956 22102 10008 22108
rect 9310 21992 9366 22001
rect 9310 21927 9366 21936
rect 9034 21856 9090 21865
rect 9034 21791 9090 21800
rect 8864 20454 8984 20482
rect 8850 20360 8906 20369
rect 7748 20324 7800 20330
rect 8850 20295 8906 20304
rect 7748 20266 7800 20272
rect 7760 20058 7788 20266
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7760 19514 7788 19994
rect 8024 19984 8076 19990
rect 8024 19926 8076 19932
rect 8036 19514 8064 19926
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8208 19780 8260 19786
rect 8208 19722 8260 19728
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 8024 19508 8076 19514
rect 8024 19450 8076 19456
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7484 18426 7512 18906
rect 8220 18766 8248 19722
rect 8312 19310 8340 19790
rect 8588 19786 8616 20198
rect 8576 19780 8628 19786
rect 8576 19722 8628 19728
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7576 17882 7604 18702
rect 7840 18148 7892 18154
rect 7840 18090 7892 18096
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7760 17066 7788 17274
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7748 17060 7800 17066
rect 7748 17002 7800 17008
rect 7668 16726 7696 17002
rect 7656 16720 7708 16726
rect 7656 16662 7708 16668
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7576 15706 7604 15982
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7760 15026 7788 15914
rect 7852 15638 7880 18090
rect 8220 17270 8248 18702
rect 8772 18154 8800 20198
rect 8864 19174 8892 20295
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8760 18148 8812 18154
rect 8760 18090 8812 18096
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8680 17270 8708 17682
rect 8208 17264 8260 17270
rect 8668 17264 8720 17270
rect 8208 17206 8260 17212
rect 8666 17232 8668 17241
rect 8720 17232 8722 17241
rect 8666 17167 8722 17176
rect 8864 16794 8892 19110
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 7932 16652 7984 16658
rect 7932 16594 7984 16600
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 7944 16182 7972 16594
rect 8496 16250 8524 16594
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 7932 16176 7984 16182
rect 7932 16118 7984 16124
rect 7944 15910 7972 16118
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8772 15910 8800 15982
rect 7932 15904 7984 15910
rect 8760 15904 8812 15910
rect 7932 15846 7984 15852
rect 8758 15872 8760 15881
rect 8812 15872 8814 15881
rect 7840 15632 7892 15638
rect 7840 15574 7892 15580
rect 7852 15162 7880 15574
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7852 14890 7880 15098
rect 7840 14884 7892 14890
rect 7840 14826 7892 14832
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7300 12986 7328 13330
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 7194 12336 7250 12345
rect 7194 12271 7196 12280
rect 7248 12271 7250 12280
rect 7196 12242 7248 12248
rect 7208 11694 7236 12242
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7392 11286 7420 11630
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6656 9722 6684 10066
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6840 9625 6868 11086
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6932 9926 6960 10542
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7300 10130 7328 10406
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9722 6960 9862
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6826 9616 6882 9625
rect 6826 9551 6882 9560
rect 7012 9376 7064 9382
rect 7010 9344 7012 9353
rect 7064 9344 7066 9353
rect 7010 9279 7066 9288
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7392 8430 7420 9114
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 6458 8256 6514 8265
rect 6458 8191 6514 8200
rect 6472 7954 6500 8191
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6366 7440 6422 7449
rect 6366 7375 6422 7384
rect 6184 7268 6236 7274
rect 6184 7210 6236 7216
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5446 6352 5502 6361
rect 5446 6287 5502 6296
rect 5460 6254 5488 6287
rect 5552 6254 5580 6802
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6012 6458 6040 6802
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6104 6322 6132 6734
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5552 5914 5580 6190
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 6196 5778 6224 7210
rect 6472 7002 6500 7890
rect 6564 7546 6592 7890
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7024 7002 7052 7278
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6918 6896 6974 6905
rect 6918 6831 6920 6840
rect 6972 6831 6974 6840
rect 6920 6802 6972 6808
rect 6932 6458 6960 6802
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 7024 6254 7052 6938
rect 7116 6934 7144 7142
rect 7104 6928 7156 6934
rect 7208 6905 7236 7822
rect 7104 6870 7156 6876
rect 7194 6896 7250 6905
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 7116 6118 7144 6870
rect 7194 6831 7250 6840
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7116 5846 7144 6054
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6196 5370 6224 5714
rect 7116 5370 7144 5782
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 6368 5092 6420 5098
rect 6368 5034 6420 5040
rect 6380 4826 6408 5034
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 7196 4616 7248 4622
rect 4066 4584 4122 4593
rect 7196 4558 7248 4564
rect 4066 4519 4122 4528
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 7208 4214 7236 4558
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 5446 3904 5502 3913
rect 5446 3839 5502 3848
rect 5460 3738 5488 3839
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 5460 2854 5488 3538
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6380 2854 6408 3538
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 5448 2848 5500 2854
rect 3514 2816 3570 2825
rect 6368 2848 6420 2854
rect 5500 2808 5580 2836
rect 5448 2790 5500 2796
rect 3514 2751 3570 2760
rect 2870 1592 2926 1601
rect 2870 1527 2926 1536
rect 3528 480 3556 2751
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4632 2553 4660 2586
rect 4618 2544 4674 2553
rect 4618 2479 4674 2488
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4632 480 4660 2382
rect 5552 1442 5580 2808
rect 6366 2816 6368 2825
rect 6420 2816 6422 2825
rect 6366 2751 6422 2760
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5552 1414 5672 1442
rect 5644 480 5672 1414
rect 6656 480 6684 2926
rect 7208 2689 7236 4150
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7392 3738 7420 3946
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7484 3618 7512 14350
rect 7576 13870 7604 14758
rect 7852 14618 7880 14826
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7562 12744 7618 12753
rect 7562 12679 7564 12688
rect 7616 12679 7618 12688
rect 7838 12744 7894 12753
rect 7838 12679 7894 12688
rect 7564 12650 7616 12656
rect 7576 12374 7604 12650
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7852 11830 7880 12679
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7944 11506 7972 15846
rect 8758 15807 8814 15816
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8220 15178 8248 15438
rect 8220 15162 8340 15178
rect 8220 15156 8352 15162
rect 8220 15150 8300 15156
rect 8300 15098 8352 15104
rect 8206 14920 8262 14929
rect 8206 14855 8262 14864
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 8036 13258 8064 13874
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 7852 11478 7972 11506
rect 7852 11218 7880 11478
rect 7930 11384 7986 11393
rect 7930 11319 7932 11328
rect 7984 11319 7986 11328
rect 7932 11290 7984 11296
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7852 10810 7880 11154
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7576 9926 7604 10474
rect 7564 9920 7616 9926
rect 7562 9888 7564 9897
rect 7616 9888 7618 9897
rect 7562 9823 7618 9832
rect 7852 9194 7880 10746
rect 7944 10266 7972 10950
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7760 9178 7880 9194
rect 7748 9172 7880 9178
rect 7800 9166 7880 9172
rect 7748 9114 7800 9120
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7576 8090 7604 8366
rect 7852 8362 7880 8910
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7852 8090 7880 8298
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7944 7002 7972 7890
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7852 5953 7880 6598
rect 7944 6361 7972 6938
rect 7930 6352 7986 6361
rect 7930 6287 7986 6296
rect 7838 5944 7894 5953
rect 7838 5879 7894 5888
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7576 5098 7604 5714
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7576 4758 7604 5034
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7576 4282 7604 4694
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7392 3590 7512 3618
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 7194 2680 7250 2689
rect 7392 2650 7420 3590
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7484 3194 7512 3470
rect 7760 3233 7788 3606
rect 7746 3224 7802 3233
rect 7472 3188 7524 3194
rect 7746 3159 7802 3168
rect 7472 3130 7524 3136
rect 7760 3126 7788 3159
rect 7748 3120 7800 3126
rect 7748 3062 7800 3068
rect 7194 2615 7250 2624
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 8036 2553 8064 13194
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12889 8156 13126
rect 8114 12880 8170 12889
rect 8114 12815 8170 12824
rect 8128 12782 8156 12815
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8220 11762 8248 14855
rect 8404 14550 8432 15506
rect 8392 14544 8444 14550
rect 8444 14492 8524 14498
rect 8392 14486 8524 14492
rect 8404 14470 8524 14486
rect 8392 14340 8444 14346
rect 8392 14282 8444 14288
rect 8404 13938 8432 14282
rect 8496 14074 8524 14470
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8298 13696 8354 13705
rect 8298 13631 8354 13640
rect 8312 12850 8340 13631
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8496 13025 8524 13126
rect 8482 13016 8538 13025
rect 8482 12951 8538 12960
rect 8496 12918 8524 12951
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8312 11898 8340 12242
rect 8588 12073 8616 13194
rect 8772 12986 8800 13330
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8758 12200 8814 12209
rect 8758 12135 8760 12144
rect 8812 12135 8814 12144
rect 8760 12106 8812 12112
rect 8574 12064 8630 12073
rect 8574 11999 8630 12008
rect 8588 11898 8616 11999
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8588 11694 8616 11834
rect 8772 11830 8800 12106
rect 8760 11824 8812 11830
rect 8760 11766 8812 11772
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 10810 8432 11494
rect 8482 11384 8538 11393
rect 8482 11319 8538 11328
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8128 9722 8156 10134
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8128 9110 8156 9318
rect 8220 9178 8248 10134
rect 8312 10062 8340 10678
rect 8496 10674 8524 11319
rect 8772 11286 8800 11766
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8850 11248 8906 11257
rect 8850 11183 8906 11192
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 8128 8498 8156 9046
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8128 8294 8156 8434
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8128 7274 8156 8230
rect 8220 7954 8248 8230
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8312 7410 8340 9998
rect 8404 9110 8432 10202
rect 8496 9926 8524 10474
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8496 9382 8524 9862
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 8300 7404 8352 7410
rect 8220 7364 8300 7392
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8114 5128 8170 5137
rect 8114 5063 8116 5072
rect 8168 5063 8170 5072
rect 8116 5034 8168 5040
rect 8128 4146 8156 5034
rect 8220 4758 8248 7364
rect 8300 7346 8352 7352
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8312 5914 8340 6258
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8128 3670 8156 4082
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8496 3233 8524 9318
rect 8772 9178 8800 9318
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8588 4146 8616 9114
rect 8666 8664 8722 8673
rect 8666 8599 8668 8608
rect 8720 8599 8722 8608
rect 8668 8570 8720 8576
rect 8680 8430 8708 8570
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8680 7546 8708 7890
rect 8760 7880 8812 7886
rect 8758 7848 8760 7857
rect 8812 7848 8814 7857
rect 8758 7783 8814 7792
rect 8864 7698 8892 11183
rect 8772 7670 8892 7698
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8666 6216 8722 6225
rect 8666 6151 8722 6160
rect 8680 5778 8708 6151
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8680 5370 8708 5714
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8482 3224 8538 3233
rect 8482 3159 8538 3168
rect 8022 2544 8078 2553
rect 8022 2479 8078 2488
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7668 480 7696 2246
rect 8772 480 8800 7670
rect 8956 4298 8984 20454
rect 9048 19310 9076 21791
rect 9324 21554 9352 21927
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 9324 21078 9352 21490
rect 9968 21350 9996 22102
rect 9956 21344 10008 21350
rect 9402 21312 9458 21321
rect 9956 21286 10008 21292
rect 9402 21247 9458 21256
rect 9312 21072 9364 21078
rect 9312 21014 9364 21020
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9140 20058 9168 20402
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 9036 19304 9088 19310
rect 9036 19246 9088 19252
rect 9048 18766 9076 19246
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 9232 17542 9260 18158
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9232 16998 9260 17478
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 9048 15706 9076 15982
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9416 14906 9444 21247
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9692 20754 9720 20810
rect 9600 20726 9720 20754
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9600 19378 9628 20726
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9692 17762 9720 18906
rect 9508 17734 9720 17762
rect 9508 17649 9536 17734
rect 9680 17672 9732 17678
rect 9494 17640 9550 17649
rect 9680 17614 9732 17620
rect 9494 17575 9550 17584
rect 9508 17134 9536 17575
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9600 16794 9628 17070
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9692 16726 9720 17614
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9692 15706 9720 15914
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9692 15416 9720 15642
rect 9600 15388 9720 15416
rect 9600 15026 9628 15388
rect 9678 15056 9734 15065
rect 9588 15020 9640 15026
rect 9678 14991 9734 15000
rect 9588 14962 9640 14968
rect 9416 14878 9628 14906
rect 9034 14784 9090 14793
rect 9034 14719 9090 14728
rect 9048 14074 9076 14719
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 9048 12782 9076 14010
rect 9140 13802 9168 14214
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9140 13190 9168 13738
rect 9232 13258 9260 13806
rect 9220 13252 9272 13258
rect 9220 13194 9272 13200
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9048 12306 9076 12718
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 9140 12209 9168 13126
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9494 12744 9550 12753
rect 9126 12200 9182 12209
rect 9126 12135 9182 12144
rect 9036 11688 9088 11694
rect 9140 11676 9168 12135
rect 9088 11648 9168 11676
rect 9036 11630 9088 11636
rect 9048 11354 9076 11630
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9416 11098 9444 12718
rect 9494 12679 9550 12688
rect 9508 12646 9536 12679
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9600 12345 9628 14878
rect 9692 13938 9720 14991
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9586 12336 9642 12345
rect 9586 12271 9642 12280
rect 9680 12300 9732 12306
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9324 11070 9444 11098
rect 9324 9738 9352 11070
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10810 9444 10950
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9508 9761 9536 11562
rect 9600 11257 9628 12271
rect 9680 12242 9732 12248
rect 9692 11558 9720 12242
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9586 11248 9642 11257
rect 9692 11234 9720 11494
rect 9784 11393 9812 20742
rect 9876 19281 9904 20878
rect 9968 20534 9996 21286
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9968 20330 9996 20470
rect 9956 20324 10008 20330
rect 9956 20266 10008 20272
rect 9968 19990 9996 20266
rect 9956 19984 10008 19990
rect 9956 19926 10008 19932
rect 10060 19802 10088 24806
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 10704 24682 10732 25094
rect 10140 24676 10192 24682
rect 10140 24618 10192 24624
rect 10692 24676 10744 24682
rect 10692 24618 10744 24624
rect 10152 23322 10180 24618
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10692 24064 10744 24070
rect 10692 24006 10744 24012
rect 10704 23594 10732 24006
rect 10692 23588 10744 23594
rect 10692 23530 10744 23536
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10704 22778 10732 23530
rect 10692 22772 10744 22778
rect 10692 22714 10744 22720
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 10152 20874 10180 21966
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10140 20868 10192 20874
rect 10140 20810 10192 20816
rect 10428 20398 10456 20946
rect 10704 20942 10732 21422
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 9968 19774 10088 19802
rect 9862 19272 9918 19281
rect 9862 19207 9918 19216
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9876 14074 9904 14350
rect 9968 14249 9996 19774
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10060 19417 10088 19654
rect 10046 19408 10102 19417
rect 10046 19343 10102 19352
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10046 18184 10102 18193
rect 10152 18154 10180 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10704 18970 10732 19246
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 10704 18222 10732 18770
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10046 18119 10102 18128
rect 10140 18148 10192 18154
rect 9954 14240 10010 14249
rect 9954 14175 10010 14184
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9876 13530 9904 14010
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9770 11384 9826 11393
rect 9770 11319 9826 11328
rect 9864 11280 9916 11286
rect 9692 11206 9812 11234
rect 9864 11222 9916 11228
rect 9586 11183 9642 11192
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9494 9752 9550 9761
rect 9324 9710 9444 9738
rect 9416 9654 9444 9710
rect 9494 9687 9550 9696
rect 9404 9648 9456 9654
rect 9310 9616 9366 9625
rect 9404 9590 9456 9596
rect 9310 9551 9366 9560
rect 9324 9518 9352 9551
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9324 8430 9352 9046
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9324 7954 9352 8366
rect 9416 8362 9444 9590
rect 9600 8514 9628 11086
rect 9680 10464 9732 10470
rect 9678 10432 9680 10441
rect 9732 10432 9734 10441
rect 9678 10367 9734 10376
rect 9678 10160 9734 10169
rect 9678 10095 9680 10104
rect 9732 10095 9734 10104
rect 9680 10066 9732 10072
rect 9692 9722 9720 10066
rect 9784 10010 9812 11206
rect 9876 10849 9904 11222
rect 9862 10840 9918 10849
rect 9862 10775 9918 10784
rect 9876 10130 9904 10775
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9784 9982 9904 10010
rect 9876 9926 9904 9982
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9600 8486 9720 8514
rect 9692 8430 9720 8486
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9232 7410 9260 7686
rect 9600 7585 9628 8298
rect 9876 8265 9904 9862
rect 9862 8256 9918 8265
rect 9862 8191 9918 8200
rect 9770 7984 9826 7993
rect 9770 7919 9772 7928
rect 9824 7919 9826 7928
rect 9772 7890 9824 7896
rect 9586 7576 9642 7585
rect 9784 7546 9812 7890
rect 9586 7511 9642 7520
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9140 7002 9168 7142
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9048 6458 9076 6734
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9048 5914 9076 6394
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9140 5098 9168 6190
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9232 5234 9260 5850
rect 9416 5846 9444 6394
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 9140 4826 9168 5034
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 8956 4270 9076 4298
rect 9048 4185 9076 4270
rect 9232 4214 9260 5170
rect 9220 4208 9272 4214
rect 9034 4176 9090 4185
rect 8944 4140 8996 4146
rect 9220 4150 9272 4156
rect 9034 4111 9090 4120
rect 8944 4082 8996 4088
rect 8956 3738 8984 4082
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9232 3534 9260 4150
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9416 3194 9444 5238
rect 9508 3670 9536 6054
rect 9692 5642 9720 7346
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9876 6458 9904 6870
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9862 5944 9918 5953
rect 9862 5879 9918 5888
rect 9876 5846 9904 5879
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9588 5296 9640 5302
rect 9692 5284 9720 5578
rect 9640 5256 9720 5284
rect 9588 5238 9640 5244
rect 9784 5137 9812 5646
rect 9876 5370 9904 5782
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9770 5128 9826 5137
rect 9770 5063 9826 5072
rect 9784 4826 9812 5063
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9588 4140 9640 4146
rect 9692 4128 9720 4422
rect 9876 4282 9904 4626
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9640 4100 9720 4128
rect 9588 4082 9640 4088
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9784 3194 9812 3606
rect 9876 3233 9904 3606
rect 9862 3224 9918 3233
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9772 3188 9824 3194
rect 9862 3159 9918 3168
rect 9772 3130 9824 3136
rect 9876 3126 9904 3159
rect 9864 3120 9916 3126
rect 9770 3088 9826 3097
rect 9864 3062 9916 3068
rect 9770 3023 9826 3032
rect 9784 480 9812 3023
rect 9968 2650 9996 13874
rect 10060 13530 10088 18119
rect 10140 18090 10192 18096
rect 10152 17814 10180 18090
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10140 17808 10192 17814
rect 10140 17750 10192 17756
rect 10152 17338 10180 17750
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16697 10732 18158
rect 10690 16688 10746 16697
rect 10140 16652 10192 16658
rect 10690 16623 10692 16632
rect 10140 16594 10192 16600
rect 10744 16623 10746 16632
rect 10692 16594 10744 16600
rect 10152 16182 10180 16594
rect 10230 16280 10286 16289
rect 10230 16215 10232 16224
rect 10284 16215 10286 16224
rect 10232 16186 10284 16192
rect 10140 16176 10192 16182
rect 10140 16118 10192 16124
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10060 12782 10088 13466
rect 10152 12986 10180 15914
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 15706 10732 16594
rect 10796 16522 10824 27520
rect 10876 25424 10928 25430
rect 10876 25366 10928 25372
rect 10888 24682 10916 25366
rect 10876 24676 10928 24682
rect 10876 24618 10928 24624
rect 11428 24676 11480 24682
rect 11428 24618 11480 24624
rect 10888 17882 10916 24618
rect 11440 24342 11468 24618
rect 10968 24336 11020 24342
rect 10968 24278 11020 24284
rect 11428 24336 11480 24342
rect 11428 24278 11480 24284
rect 10980 23526 11008 24278
rect 11440 23882 11468 24278
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11256 23854 11468 23882
rect 11532 23866 11560 24142
rect 11520 23860 11572 23866
rect 11256 23798 11284 23854
rect 11520 23802 11572 23808
rect 11244 23792 11296 23798
rect 11808 23769 11836 27520
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 12162 23896 12218 23905
rect 12162 23831 12164 23840
rect 12216 23831 12218 23840
rect 12164 23802 12216 23808
rect 11244 23734 11296 23740
rect 11794 23760 11850 23769
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10980 23304 11008 23462
rect 10980 23276 11100 23304
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 10980 22574 11008 23122
rect 10968 22568 11020 22574
rect 10966 22536 10968 22545
rect 11020 22536 11022 22545
rect 10966 22471 11022 22480
rect 11072 22386 11100 23276
rect 11256 23118 11284 23734
rect 11794 23695 11850 23704
rect 12176 23594 12204 23802
rect 12544 23730 12572 25094
rect 12728 24954 12756 25298
rect 12716 24948 12768 24954
rect 12716 24890 12768 24896
rect 12728 24449 12756 24890
rect 12714 24440 12770 24449
rect 12714 24375 12770 24384
rect 12714 24304 12770 24313
rect 12714 24239 12770 24248
rect 12728 24206 12756 24239
rect 12716 24200 12768 24206
rect 12716 24142 12768 24148
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 11428 23588 11480 23594
rect 11428 23530 11480 23536
rect 12164 23588 12216 23594
rect 12164 23530 12216 23536
rect 11336 23248 11388 23254
rect 11336 23190 11388 23196
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11256 22710 11284 23054
rect 11348 22778 11376 23190
rect 11440 23118 11468 23530
rect 11428 23112 11480 23118
rect 11428 23054 11480 23060
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11244 22704 11296 22710
rect 11244 22646 11296 22652
rect 10980 22358 11100 22386
rect 10980 21162 11008 22358
rect 11348 22234 11376 22714
rect 11336 22228 11388 22234
rect 11336 22170 11388 22176
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11900 21690 11928 21966
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11334 21448 11390 21457
rect 11334 21383 11336 21392
rect 11388 21383 11390 21392
rect 11336 21354 11388 21360
rect 10980 21146 11100 21162
rect 10980 21140 11112 21146
rect 10980 21134 11060 21140
rect 11060 21082 11112 21088
rect 10966 20632 11022 20641
rect 11072 20602 11100 21082
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 10966 20567 11022 20576
rect 11060 20596 11112 20602
rect 10980 18902 11008 20567
rect 11060 20538 11112 20544
rect 11164 20466 11192 20878
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 11348 19310 11376 21354
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11624 19718 11652 20878
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 11888 20052 11940 20058
rect 11888 19994 11940 20000
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 11072 18970 11100 19246
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 11072 18834 11100 18906
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 10980 18086 11008 18702
rect 11164 18426 11192 18838
rect 11624 18766 11652 19654
rect 11900 19514 11928 19994
rect 11992 19961 12020 20198
rect 11978 19952 12034 19961
rect 11978 19887 12034 19896
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 12176 18902 12204 23530
rect 12544 23322 12572 23666
rect 12728 23322 12756 24142
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12716 23316 12768 23322
rect 12716 23258 12768 23264
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12636 22574 12664 23054
rect 12624 22568 12676 22574
rect 12624 22510 12676 22516
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 12268 21350 12296 22034
rect 12440 21412 12492 21418
rect 12440 21354 12492 21360
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12268 21078 12296 21286
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 12268 20534 12296 21014
rect 12256 20528 12308 20534
rect 12256 20470 12308 20476
rect 12268 20398 12296 20470
rect 12452 20398 12480 21354
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12268 19854 12296 20334
rect 12636 19990 12664 22510
rect 12808 20936 12860 20942
rect 12808 20878 12860 20884
rect 12820 20641 12848 20878
rect 12806 20632 12862 20641
rect 12806 20567 12862 20576
rect 12624 19984 12676 19990
rect 12624 19926 12676 19932
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12440 19236 12492 19242
rect 12440 19178 12492 19184
rect 12452 18970 12480 19178
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12164 18896 12216 18902
rect 12164 18838 12216 18844
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11886 18728 11942 18737
rect 11348 18426 11376 18702
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11336 18420 11388 18426
rect 11336 18362 11388 18368
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10888 17338 10916 17818
rect 10980 17626 11008 18022
rect 11348 17882 11376 18362
rect 11336 17876 11388 17882
rect 11336 17818 11388 17824
rect 10980 17598 11100 17626
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10888 17066 10916 17274
rect 10980 17202 11008 17478
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 11072 17082 11100 17598
rect 11624 17270 11652 18702
rect 11886 18663 11942 18672
rect 11900 18426 11928 18663
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11900 18222 11928 18362
rect 12452 18290 12480 18906
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12176 17814 12204 18022
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 10876 17060 10928 17066
rect 10876 17002 10928 17008
rect 10980 17054 11100 17082
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10692 15496 10744 15502
rect 10506 15464 10562 15473
rect 10692 15438 10744 15444
rect 10506 15399 10562 15408
rect 10520 15162 10548 15399
rect 10704 15337 10732 15438
rect 10690 15328 10746 15337
rect 10690 15263 10746 15272
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10244 14890 10272 15030
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 10520 14804 10548 15098
rect 10520 14776 10732 14804
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14618 10732 14776
rect 10692 14612 10744 14618
rect 10612 14572 10692 14600
rect 10612 14074 10640 14572
rect 10692 14554 10744 14560
rect 10796 14521 10824 15846
rect 10876 15632 10928 15638
rect 10876 15574 10928 15580
rect 10888 14890 10916 15574
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10782 14512 10838 14521
rect 10782 14447 10838 14456
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10612 13870 10640 14010
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10704 13705 10732 14350
rect 10874 14240 10930 14249
rect 10874 14175 10930 14184
rect 10690 13696 10746 13705
rect 10289 13628 10585 13648
rect 10690 13631 10746 13640
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10060 12306 10088 12582
rect 10152 12306 10180 12922
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10428 11898 10456 12242
rect 10796 12238 10824 13262
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10888 11778 10916 14175
rect 10980 12646 11008 17054
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11164 15094 11192 16730
rect 11808 16726 11836 17614
rect 12176 17338 12204 17750
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 11796 16720 11848 16726
rect 11980 16720 12032 16726
rect 11796 16662 11848 16668
rect 11978 16688 11980 16697
rect 12348 16720 12400 16726
rect 12032 16688 12034 16697
rect 12348 16662 12400 16668
rect 11978 16623 12034 16632
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 11348 15638 11376 16526
rect 11992 15706 12020 16623
rect 12360 15910 12388 16662
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12636 15978 12664 16390
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12360 15638 12388 15846
rect 11336 15632 11388 15638
rect 12348 15632 12400 15638
rect 11388 15592 11468 15620
rect 11336 15574 11388 15580
rect 11242 15328 11298 15337
rect 11242 15263 11298 15272
rect 11256 15162 11284 15263
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11072 14550 11100 15030
rect 11336 14952 11388 14958
rect 11334 14920 11336 14929
rect 11388 14920 11390 14929
rect 11334 14855 11390 14864
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11164 13938 11192 14214
rect 11440 14006 11468 15592
rect 12348 15574 12400 15580
rect 12360 15026 12388 15574
rect 12636 15473 12664 15914
rect 12622 15464 12678 15473
rect 12440 15428 12492 15434
rect 12622 15399 12678 15408
rect 12440 15370 12492 15376
rect 12452 15094 12480 15370
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11428 14000 11480 14006
rect 11428 13942 11480 13948
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11256 13462 11284 13670
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 11256 12646 11284 13398
rect 11440 13326 11468 13942
rect 11716 13734 11744 14486
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11992 13190 12020 14350
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12268 13462 12296 14214
rect 12452 13802 12480 15030
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12728 14618 12756 14758
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 13938 12848 14214
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12820 13802 12848 13874
rect 12440 13796 12492 13802
rect 12440 13738 12492 13744
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12452 13530 12480 13738
rect 12530 13696 12586 13705
rect 12530 13631 12586 13640
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11716 12986 11744 13126
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11992 12850 12020 13126
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 10704 11750 10916 11778
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10060 10810 10088 11154
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10060 10198 10088 10746
rect 10152 10674 10180 11290
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10152 10266 10180 10610
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10060 8498 10088 8910
rect 10152 8566 10180 9046
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10060 8090 10088 8434
rect 10152 8362 10180 8502
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10152 6882 10180 8298
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10508 7472 10560 7478
rect 10506 7440 10508 7449
rect 10560 7440 10562 7449
rect 10506 7375 10562 7384
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10152 6854 10272 6882
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5817 10088 6054
rect 10152 5914 10180 6734
rect 10244 6458 10272 6854
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10046 5808 10102 5817
rect 10046 5743 10102 5752
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10704 4706 10732 11750
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10980 9654 11008 11494
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11072 10713 11100 11154
rect 11058 10704 11114 10713
rect 11058 10639 11114 10648
rect 11072 10470 11100 10639
rect 11256 10538 11284 12582
rect 12084 12442 12112 13262
rect 12268 12918 12296 13398
rect 12544 13258 12572 13631
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 12438 13016 12494 13025
rect 12438 12951 12494 12960
rect 12256 12912 12308 12918
rect 12256 12854 12308 12860
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 11518 12336 11574 12345
rect 11518 12271 11520 12280
rect 11572 12271 11574 12280
rect 12164 12300 12216 12306
rect 11520 12242 11572 12248
rect 12164 12242 12216 12248
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11244 10532 11296 10538
rect 11244 10474 11296 10480
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10980 9450 11008 9590
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 10796 8906 10824 9318
rect 11348 9178 11376 9318
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10612 4690 10732 4706
rect 10600 4684 10732 4690
rect 10652 4678 10732 4684
rect 10600 4626 10652 4632
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10060 3913 10088 3946
rect 10152 3942 10180 4558
rect 10704 4049 10732 4678
rect 10690 4040 10746 4049
rect 10690 3975 10746 3984
rect 10140 3936 10192 3942
rect 10046 3904 10102 3913
rect 10140 3878 10192 3884
rect 10690 3904 10746 3913
rect 10046 3839 10102 3848
rect 10152 3641 10180 3878
rect 10289 3836 10585 3856
rect 10690 3839 10746 3848
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10138 3632 10194 3641
rect 10138 3567 10194 3576
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9876 2417 9904 2450
rect 9862 2408 9918 2417
rect 9862 2343 9918 2352
rect 10704 1034 10732 3839
rect 10796 2650 10824 8842
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 10888 8090 10916 8366
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10980 7970 11008 8230
rect 10888 7954 11008 7970
rect 10876 7948 11008 7954
rect 10928 7942 11008 7948
rect 10876 7890 10928 7896
rect 10888 7342 10916 7890
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10888 7002 10916 7278
rect 11256 7002 11284 7346
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11150 6896 11206 6905
rect 11150 6831 11152 6840
rect 11204 6831 11206 6840
rect 11152 6802 11204 6808
rect 11164 5914 11192 6802
rect 11256 6322 11284 6938
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10980 5234 11008 5646
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 11072 5098 11100 5578
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 11348 5030 11376 8366
rect 11440 8022 11468 12038
rect 11532 11898 11560 12242
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11716 11694 11744 12174
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 11716 10470 11744 11630
rect 12084 11354 12112 11630
rect 12176 11558 12204 12242
rect 12452 12102 12480 12951
rect 12544 12850 12572 13194
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12636 12714 12664 12922
rect 12728 12850 12756 13262
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11886 10568 11942 10577
rect 11886 10503 11942 10512
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11532 9450 11560 9998
rect 11520 9444 11572 9450
rect 11520 9386 11572 9392
rect 11532 9042 11560 9386
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11532 7886 11560 8978
rect 11716 8022 11744 10406
rect 11900 10198 11928 10503
rect 12084 10266 12112 11290
rect 12176 11218 12204 11494
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12176 10810 12204 11154
rect 12268 11082 12296 11222
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12268 10810 12296 11018
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12176 10606 12204 10746
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 12084 9722 12112 10202
rect 12452 10130 12480 11290
rect 12636 10538 12664 12038
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12636 10266 12664 10474
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12164 9920 12216 9926
rect 12162 9888 12164 9897
rect 12216 9888 12218 9897
rect 12162 9823 12218 9832
rect 12438 9752 12494 9761
rect 12072 9716 12124 9722
rect 12438 9687 12494 9696
rect 12072 9658 12124 9664
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12176 8430 12204 9046
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11716 7546 11744 7958
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11624 6934 11652 7142
rect 11612 6928 11664 6934
rect 11612 6870 11664 6876
rect 11624 6186 11652 6870
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11808 5642 11836 6394
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11808 5370 11836 5578
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 10888 4758 10916 4966
rect 11532 4758 11560 5034
rect 10876 4752 10928 4758
rect 10876 4694 10928 4700
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 10888 4282 10916 4694
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 11532 4146 11560 4694
rect 11794 4176 11850 4185
rect 11520 4140 11572 4146
rect 11794 4111 11850 4120
rect 11520 4082 11572 4088
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10888 3738 10916 3946
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10980 3602 11008 3946
rect 11808 3602 11836 4111
rect 11992 3738 12020 5034
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 12084 4078 12112 4694
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12176 4026 12204 6598
rect 12268 5216 12296 9318
rect 12346 9072 12402 9081
rect 12346 9007 12402 9016
rect 12360 8974 12388 9007
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12452 8430 12480 9687
rect 12530 9616 12586 9625
rect 12530 9551 12532 9560
rect 12584 9551 12586 9560
rect 12532 9522 12584 9528
rect 12544 8906 12572 9522
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12622 8392 12678 8401
rect 12622 8327 12678 8336
rect 12438 7848 12494 7857
rect 12438 7783 12440 7792
rect 12492 7783 12494 7792
rect 12440 7754 12492 7760
rect 12452 7410 12480 7754
rect 12530 7576 12586 7585
rect 12530 7511 12586 7520
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12544 6866 12572 7511
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12544 6322 12572 6802
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12636 5846 12664 8327
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12532 5228 12584 5234
rect 12268 5188 12388 5216
rect 12360 4758 12388 5188
rect 12532 5170 12584 5176
rect 12544 5098 12572 5170
rect 12636 5098 12664 5238
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12360 4282 12388 4558
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12176 3998 12480 4026
rect 12544 4010 12572 4082
rect 12452 3942 12480 3998
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 3738 12480 3878
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12544 3670 12572 3946
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 11808 3194 11836 3538
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 12728 2990 12756 12786
rect 12912 12050 12940 27520
rect 13450 24848 13506 24857
rect 13450 24783 13506 24792
rect 13268 24744 13320 24750
rect 13268 24686 13320 24692
rect 12992 24336 13044 24342
rect 12992 24278 13044 24284
rect 13004 23526 13032 24278
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 13004 21418 13032 23462
rect 13280 22778 13308 24686
rect 13464 24614 13492 24783
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13556 23730 13584 24142
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13726 23488 13782 23497
rect 13726 23423 13782 23432
rect 13740 23118 13768 23423
rect 13820 23248 13872 23254
rect 13820 23190 13872 23196
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13740 22778 13768 23054
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 13726 22536 13782 22545
rect 13726 22471 13782 22480
rect 13740 21690 13768 22471
rect 13832 22438 13860 23190
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 13004 21146 13032 21354
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 13004 19938 13032 21082
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 13740 20602 13768 20878
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 13832 20398 13860 22374
rect 13268 20392 13320 20398
rect 13268 20334 13320 20340
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 13280 20058 13308 20334
rect 13268 20052 13320 20058
rect 13268 19994 13320 20000
rect 13832 19990 13860 20334
rect 13820 19984 13872 19990
rect 13004 19910 13308 19938
rect 13820 19926 13872 19932
rect 13924 19938 13952 27520
rect 14936 25242 14964 27520
rect 14384 25214 14964 25242
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 14108 23633 14136 24006
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 14094 23624 14150 23633
rect 14094 23559 14096 23568
rect 14148 23559 14150 23568
rect 14096 23530 14148 23536
rect 14200 23118 14228 23666
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 14200 22642 14228 23054
rect 14188 22636 14240 22642
rect 14188 22578 14240 22584
rect 14004 22500 14056 22506
rect 14004 22442 14056 22448
rect 14016 22234 14044 22442
rect 14200 22234 14228 22578
rect 14004 22228 14056 22234
rect 14004 22170 14056 22176
rect 14188 22228 14240 22234
rect 14188 22170 14240 22176
rect 14280 21888 14332 21894
rect 14280 21830 14332 21836
rect 14292 21622 14320 21830
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14292 21418 14320 21558
rect 14280 21412 14332 21418
rect 14280 21354 14332 21360
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 14016 21146 14044 21286
rect 14004 21140 14056 21146
rect 14004 21082 14056 21088
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14108 19990 14136 20402
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14096 19984 14148 19990
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 13004 19514 13032 19790
rect 12992 19508 13044 19514
rect 12992 19450 13044 19456
rect 13004 19242 13032 19450
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 13096 18970 13124 19246
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13188 18193 13216 18702
rect 13280 18222 13308 19910
rect 13832 19446 13860 19926
rect 13924 19910 14044 19938
rect 14096 19926 14148 19932
rect 13912 19780 13964 19786
rect 13912 19722 13964 19728
rect 13820 19440 13872 19446
rect 13820 19382 13872 19388
rect 13924 18970 13952 19722
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13372 18426 13400 18770
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13268 18216 13320 18222
rect 13174 18184 13230 18193
rect 13268 18158 13320 18164
rect 13174 18119 13230 18128
rect 13820 18148 13872 18154
rect 13188 17882 13216 18119
rect 13820 18090 13872 18096
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 13634 17776 13690 17785
rect 13464 17338 13492 17750
rect 13634 17711 13690 17720
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13648 17134 13676 17711
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 13004 16833 13032 16934
rect 12990 16824 13046 16833
rect 13740 16794 13768 17614
rect 13832 17338 13860 18090
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 12990 16759 13046 16768
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 16250 13400 16390
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 13188 15094 13216 15914
rect 13464 15910 13492 16594
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 13464 14929 13492 15846
rect 13556 15706 13584 15846
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13556 15026 13584 15642
rect 13740 15570 13768 16458
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13740 15162 13768 15506
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13450 14920 13506 14929
rect 13506 14878 13584 14906
rect 13450 14855 13506 14864
rect 13452 14544 13504 14550
rect 13082 14512 13138 14521
rect 13452 14486 13504 14492
rect 13082 14447 13084 14456
rect 13136 14447 13138 14456
rect 13084 14418 13136 14424
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13004 13326 13032 13874
rect 13096 13530 13124 14418
rect 13464 13734 13492 14486
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 13450 12880 13506 12889
rect 13450 12815 13452 12824
rect 13504 12815 13506 12824
rect 13452 12786 13504 12792
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 12912 12022 13032 12050
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12912 11218 12940 11834
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12912 10849 12940 11154
rect 13004 11121 13032 12022
rect 13372 11898 13400 12242
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13556 11336 13584 14878
rect 13740 12918 13768 15098
rect 13728 12912 13780 12918
rect 13728 12854 13780 12860
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13832 12442 13860 12582
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13832 12073 13860 12378
rect 13818 12064 13874 12073
rect 13818 11999 13874 12008
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13464 11308 13584 11336
rect 12990 11112 13046 11121
rect 12990 11047 13046 11056
rect 12898 10840 12954 10849
rect 12898 10775 12900 10784
rect 12952 10775 12954 10784
rect 12900 10746 12952 10752
rect 12912 10715 12940 10746
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13096 10198 13124 10406
rect 13372 10198 13400 10542
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13360 10192 13412 10198
rect 13360 10134 13412 10140
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13004 9110 13032 9522
rect 13096 9382 13124 10134
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12992 9104 13044 9110
rect 12898 9072 12954 9081
rect 12992 9046 13044 9052
rect 12898 9007 12954 9016
rect 12912 8090 12940 9007
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 13004 6730 13032 9046
rect 13096 7546 13124 9318
rect 13280 9178 13308 10066
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13096 7274 13124 7482
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 13176 6928 13228 6934
rect 13176 6870 13228 6876
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 13188 6458 13216 6870
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13188 5914 13216 6394
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 12912 4826 12940 5850
rect 13280 5710 13308 6734
rect 13464 6225 13492 11308
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13556 9926 13584 11154
rect 13648 10266 13676 11630
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13556 9042 13584 9862
rect 13740 9602 13768 11562
rect 13820 9648 13872 9654
rect 13740 9596 13820 9602
rect 13740 9590 13872 9596
rect 13740 9574 13860 9590
rect 13832 9450 13860 9574
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13556 8634 13584 8978
rect 13740 8634 13768 9318
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13740 7478 13768 7822
rect 13728 7472 13780 7478
rect 13728 7414 13780 7420
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13450 6216 13506 6225
rect 13450 6151 13506 6160
rect 13268 5704 13320 5710
rect 13636 5704 13688 5710
rect 13268 5646 13320 5652
rect 13634 5672 13636 5681
rect 13688 5672 13690 5681
rect 13084 5636 13136 5642
rect 13634 5607 13690 5616
rect 13084 5578 13136 5584
rect 13096 5302 13124 5578
rect 13740 5522 13768 7278
rect 13832 7274 13860 7958
rect 13924 7342 13952 15982
rect 14016 13938 14044 19910
rect 14200 19514 14228 20198
rect 14384 19938 14412 25214
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15948 24818 15976 27520
rect 15936 24812 15988 24818
rect 15936 24754 15988 24760
rect 16212 24608 16264 24614
rect 16212 24550 16264 24556
rect 15384 24268 15436 24274
rect 15384 24210 15436 24216
rect 15292 24064 15344 24070
rect 15292 24006 15344 24012
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15108 23588 15160 23594
rect 15108 23530 15160 23536
rect 15120 23338 15148 23530
rect 15304 23497 15332 24006
rect 15396 23662 15424 24210
rect 15934 24032 15990 24041
rect 15934 23967 15990 23976
rect 15948 23866 15976 23967
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 15384 23656 15436 23662
rect 15382 23624 15384 23633
rect 15436 23624 15438 23633
rect 15382 23559 15438 23568
rect 15290 23488 15346 23497
rect 15290 23423 15346 23432
rect 15120 23310 15516 23338
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15304 22642 15332 23122
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15396 22545 15424 22918
rect 15382 22536 15438 22545
rect 14740 22500 14792 22506
rect 15382 22471 15438 22480
rect 14740 22442 14792 22448
rect 14648 22432 14700 22438
rect 14554 22400 14610 22409
rect 14648 22374 14700 22380
rect 14554 22335 14610 22344
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14476 20330 14504 20742
rect 14464 20324 14516 20330
rect 14464 20266 14516 20272
rect 14292 19910 14412 19938
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14292 18714 14320 19910
rect 14372 19848 14424 19854
rect 14476 19836 14504 20266
rect 14424 19808 14504 19836
rect 14372 19790 14424 19796
rect 14200 18686 14320 18714
rect 14096 17128 14148 17134
rect 14094 17096 14096 17105
rect 14148 17096 14150 17105
rect 14094 17031 14150 17040
rect 14200 16182 14228 18686
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14292 18154 14320 18566
rect 14384 18290 14412 19790
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 14384 17814 14412 18226
rect 14372 17808 14424 17814
rect 14372 17750 14424 17756
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14188 16176 14240 16182
rect 14188 16118 14240 16124
rect 14476 15337 14504 16934
rect 14462 15328 14518 15337
rect 14462 15263 14518 15272
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 14016 12306 14044 13262
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14016 10674 14044 10950
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10198 14044 10610
rect 14004 10192 14056 10198
rect 14004 10134 14056 10140
rect 14016 9178 14044 10134
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14108 8401 14136 14758
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14384 13530 14412 13670
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14384 12782 14412 13330
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14372 12776 14424 12782
rect 14186 12744 14242 12753
rect 14372 12718 14424 12724
rect 14186 12679 14242 12688
rect 14200 12646 14228 12679
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14200 11898 14228 12582
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14186 11112 14242 11121
rect 14186 11047 14242 11056
rect 14094 8392 14150 8401
rect 14094 8327 14150 8336
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 14016 5914 14044 6666
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 13740 5494 13860 5522
rect 13832 5370 13860 5494
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 13096 4758 13124 5238
rect 13832 5030 13860 5306
rect 14016 5302 14044 5850
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 14200 4690 14228 11047
rect 14292 8498 14320 12106
rect 14384 12102 14412 12718
rect 14476 12374 14504 13126
rect 14464 12368 14516 12374
rect 14464 12310 14516 12316
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14384 9178 14412 9522
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14292 8090 14320 8434
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14292 6322 14320 6598
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14292 5642 14320 6258
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14384 5234 14412 6258
rect 14568 5778 14596 22335
rect 14660 21894 14688 22374
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14752 21554 14780 22442
rect 15384 22432 15436 22438
rect 15384 22374 15436 22380
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14752 20466 14780 21490
rect 15014 21448 15070 21457
rect 15014 21383 15070 21392
rect 15028 21146 15056 21383
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 15304 21049 15332 21286
rect 15396 21078 15424 22374
rect 15488 21078 15516 23310
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15752 22092 15804 22098
rect 15752 22034 15804 22040
rect 15580 21350 15608 22034
rect 15764 21457 15792 22034
rect 16028 21616 16080 21622
rect 16028 21558 16080 21564
rect 15750 21448 15806 21457
rect 15750 21383 15806 21392
rect 15844 21412 15896 21418
rect 15844 21354 15896 21360
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15856 21146 15884 21354
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 15384 21072 15436 21078
rect 15290 21040 15346 21049
rect 15384 21014 15436 21020
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15290 20975 15346 20984
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15396 20602 15424 21014
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15488 20534 15516 21014
rect 15476 20528 15528 20534
rect 15476 20470 15528 20476
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14646 19952 14702 19961
rect 14646 19887 14702 19896
rect 14660 17338 14688 19887
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15198 19408 15254 19417
rect 15198 19343 15254 19352
rect 14924 19304 14976 19310
rect 14924 19246 14976 19252
rect 14936 18970 14964 19246
rect 15212 19174 15240 19343
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 14924 18964 14976 18970
rect 14924 18906 14976 18912
rect 14936 18766 14964 18906
rect 15382 18864 15438 18873
rect 15382 18799 15384 18808
rect 15436 18799 15438 18808
rect 15384 18770 15436 18776
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 15290 18728 15346 18737
rect 15290 18663 15346 18672
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14660 17134 14688 17274
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 15200 16720 15252 16726
rect 15198 16688 15200 16697
rect 15252 16688 15254 16697
rect 15304 16658 15332 18663
rect 15396 18426 15424 18770
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15488 17882 15516 20470
rect 15856 20466 15884 21082
rect 16040 21078 16068 21558
rect 16028 21072 16080 21078
rect 16028 21014 16080 21020
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 16040 19446 16068 19858
rect 16028 19440 16080 19446
rect 16026 19408 16028 19417
rect 16080 19408 16082 19417
rect 16026 19343 16082 19352
rect 15936 18624 15988 18630
rect 15936 18566 15988 18572
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15396 17513 15424 17682
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15382 17504 15438 17513
rect 15382 17439 15438 17448
rect 15396 17338 15424 17439
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15396 17241 15424 17274
rect 15382 17232 15438 17241
rect 15382 17167 15438 17176
rect 15764 16998 15792 17614
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15566 16688 15622 16697
rect 15198 16623 15254 16632
rect 15292 16652 15344 16658
rect 15566 16623 15622 16632
rect 15292 16594 15344 16600
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16182 15332 16594
rect 15580 16250 15608 16623
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15580 16046 15608 16186
rect 15672 16046 15700 16390
rect 15568 16040 15620 16046
rect 14830 16008 14886 16017
rect 15568 15982 15620 15988
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 14830 15943 14886 15952
rect 14844 15473 14872 15943
rect 15568 15496 15620 15502
rect 14830 15464 14886 15473
rect 15568 15438 15620 15444
rect 14830 15399 14886 15408
rect 14844 15162 14872 15399
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14844 14958 14872 15098
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14660 14249 14688 14418
rect 14740 14272 14792 14278
rect 14646 14240 14702 14249
rect 14740 14214 14792 14220
rect 14646 14175 14702 14184
rect 14660 14074 14688 14175
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14660 12186 14688 13874
rect 14752 13870 14780 14214
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15304 13938 15332 15302
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 14278 15516 14894
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 15304 13326 15332 13874
rect 15488 13870 15516 14214
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15488 13530 15516 13806
rect 15580 13802 15608 15438
rect 15672 14822 15700 15982
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15764 14618 15792 16934
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15856 14278 15884 14894
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15856 14006 15884 14214
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15856 13870 15884 13942
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15488 13394 15516 13466
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15580 12782 15608 13194
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15304 12442 15332 12718
rect 15844 12708 15896 12714
rect 15844 12650 15896 12656
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15292 12436 15344 12442
rect 15344 12396 15424 12424
rect 15292 12378 15344 12384
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15304 12209 15332 12242
rect 15290 12200 15346 12209
rect 14660 12158 14780 12186
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 11694 14688 12038
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14646 10568 14702 10577
rect 14646 10503 14702 10512
rect 14660 9654 14688 10503
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14752 6474 14780 12158
rect 15290 12135 15346 12144
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15396 11694 15424 12396
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15396 11354 15424 11630
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14844 10690 14872 11018
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10742 15332 11154
rect 15292 10736 15344 10742
rect 15290 10704 15292 10713
rect 15344 10704 15346 10713
rect 14844 10662 14964 10690
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 14844 9042 14872 10474
rect 14936 10266 14964 10662
rect 15290 10639 15346 10648
rect 15488 10606 15516 12174
rect 15580 11286 15608 12582
rect 15856 12345 15884 12650
rect 15842 12336 15898 12345
rect 15842 12271 15898 12280
rect 15752 11688 15804 11694
rect 15658 11656 15714 11665
rect 15752 11630 15804 11636
rect 15658 11591 15714 11600
rect 15672 11354 15700 11591
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9722 15332 9998
rect 15488 9722 15516 10542
rect 15764 10198 15792 11630
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15948 9625 15976 18566
rect 16224 17882 16252 24550
rect 16304 24268 16356 24274
rect 16304 24210 16356 24216
rect 16316 23866 16344 24210
rect 16486 24168 16542 24177
rect 16486 24103 16488 24112
rect 16540 24103 16542 24112
rect 16488 24074 16540 24080
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 16488 23860 16540 23866
rect 16488 23802 16540 23808
rect 16396 23520 16448 23526
rect 16396 23462 16448 23468
rect 16408 23322 16436 23462
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16304 23180 16356 23186
rect 16304 23122 16356 23128
rect 16316 22506 16344 23122
rect 16500 22778 16528 23802
rect 16856 23656 16908 23662
rect 16856 23598 16908 23604
rect 16488 22772 16540 22778
rect 16488 22714 16540 22720
rect 16304 22500 16356 22506
rect 16304 22442 16356 22448
rect 16316 22001 16344 22442
rect 16302 21992 16358 22001
rect 16302 21927 16358 21936
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16316 21418 16344 21830
rect 16868 21593 16896 23598
rect 17052 23186 17080 27520
rect 18064 24041 18092 27520
rect 18234 24712 18290 24721
rect 18234 24647 18290 24656
rect 18248 24410 18276 24647
rect 18236 24404 18288 24410
rect 18236 24346 18288 24352
rect 18420 24268 18472 24274
rect 18420 24210 18472 24216
rect 18050 24032 18106 24041
rect 18050 23967 18106 23976
rect 17130 23896 17186 23905
rect 17130 23831 17132 23840
rect 17184 23831 17186 23840
rect 17132 23802 17184 23808
rect 18050 23760 18106 23769
rect 17132 23724 17184 23730
rect 18050 23695 18106 23704
rect 17132 23666 17184 23672
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 17052 22778 17080 23122
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 17144 22438 17172 23666
rect 18064 23662 18092 23695
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18432 23526 18460 24210
rect 19076 23905 19104 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 20088 24721 20116 27520
rect 20074 24712 20130 24721
rect 20074 24647 20130 24656
rect 19430 24576 19486 24585
rect 19430 24511 19486 24520
rect 19062 23896 19118 23905
rect 19062 23831 19118 23840
rect 19246 23896 19302 23905
rect 19246 23831 19248 23840
rect 19300 23831 19302 23840
rect 19248 23802 19300 23808
rect 19444 23730 19472 24511
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20626 24304 20682 24313
rect 20626 24239 20682 24248
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 18512 23656 18564 23662
rect 20640 23633 20668 24239
rect 21192 23905 21220 27520
rect 22204 24857 22232 27520
rect 22190 24848 22246 24857
rect 22190 24783 22246 24792
rect 22374 24304 22430 24313
rect 22374 24239 22430 24248
rect 21270 24032 21326 24041
rect 21270 23967 21326 23976
rect 21178 23896 21234 23905
rect 21284 23866 21312 23967
rect 22388 23866 22416 24239
rect 23216 24041 23244 27520
rect 23662 27296 23718 27305
rect 23662 27231 23718 27240
rect 23202 24032 23258 24041
rect 23202 23967 23258 23976
rect 21178 23831 21234 23840
rect 21272 23860 21324 23866
rect 21272 23802 21324 23808
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22192 23656 22244 23662
rect 18512 23598 18564 23604
rect 20626 23624 20682 23633
rect 18420 23520 18472 23526
rect 18420 23462 18472 23468
rect 17868 22976 17920 22982
rect 17868 22918 17920 22924
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 17132 22432 17184 22438
rect 17132 22374 17184 22380
rect 17038 21992 17094 22001
rect 17038 21927 17040 21936
rect 17092 21927 17094 21936
rect 17040 21898 17092 21904
rect 16854 21584 16910 21593
rect 16854 21519 16910 21528
rect 16304 21412 16356 21418
rect 16304 21354 16356 21360
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16132 13818 16160 17478
rect 16224 17270 16252 17818
rect 16592 17814 16620 18158
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16580 17808 16632 17814
rect 16500 17768 16580 17796
rect 16212 17264 16264 17270
rect 16212 17206 16264 17212
rect 16500 16998 16528 17768
rect 16580 17750 16632 17756
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16224 15978 16252 16390
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 16224 15638 16252 15914
rect 16500 15706 16528 16934
rect 16684 16726 16712 17614
rect 16776 17066 16804 18022
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 16960 17066 16988 17546
rect 17040 17128 17092 17134
rect 17040 17070 17092 17076
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 16948 17060 17000 17066
rect 16948 17002 17000 17008
rect 16776 16726 16804 17002
rect 16672 16720 16724 16726
rect 16672 16662 16724 16668
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16684 15706 16712 16662
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16224 15162 16252 15574
rect 16960 15502 16988 17002
rect 17052 16250 17080 17070
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 17052 15638 17080 16186
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16212 15156 16264 15162
rect 16264 15116 16344 15144
rect 16212 15098 16264 15104
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16224 13938 16252 14894
rect 16316 14074 16344 15116
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16132 13790 16252 13818
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16040 12238 16068 12922
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16132 10606 16160 11562
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16132 10266 16160 10542
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 15934 9616 15990 9625
rect 15934 9551 15990 9560
rect 16224 9466 16252 13790
rect 16592 13394 16620 14418
rect 16684 14278 16712 14418
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16684 13870 16712 14214
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16684 13394 16712 13806
rect 16856 13796 16908 13802
rect 16856 13738 16908 13744
rect 16868 13682 16896 13738
rect 17052 13734 17080 14418
rect 17040 13728 17092 13734
rect 16868 13654 16988 13682
rect 17040 13670 17092 13676
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16592 12986 16620 13330
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16684 12646 16712 13330
rect 16868 12714 16896 13330
rect 16960 13326 16988 13654
rect 17052 13394 17080 13670
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16960 12782 16988 13262
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16856 12708 16908 12714
rect 16856 12650 16908 12656
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 11218 16436 12038
rect 16580 11552 16632 11558
rect 16684 11540 16712 12582
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16776 11694 16804 12242
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16632 11512 16712 11540
rect 16580 11494 16632 11500
rect 16592 11218 16620 11494
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16408 10538 16436 11154
rect 16592 10810 16620 11154
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16396 10532 16448 10538
rect 16396 10474 16448 10480
rect 16408 10130 16436 10474
rect 16592 10130 16620 10746
rect 16684 10606 16712 11290
rect 16960 11014 16988 12718
rect 17144 12424 17172 22374
rect 17236 22166 17264 22578
rect 17224 22160 17276 22166
rect 17224 22102 17276 22108
rect 17236 21350 17264 22102
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17236 15881 17264 21286
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17880 16674 17908 22918
rect 18432 22409 18460 23462
rect 18418 22400 18474 22409
rect 18418 22335 18474 22344
rect 18052 17060 18104 17066
rect 18052 17002 18104 17008
rect 17328 16250 17356 16662
rect 17880 16646 18000 16674
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17222 15872 17278 15881
rect 17222 15807 17278 15816
rect 17052 12396 17172 12424
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16960 10606 16988 10950
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16396 10124 16448 10130
rect 16580 10124 16632 10130
rect 16396 10066 16448 10072
rect 16500 10084 16580 10112
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 16132 9438 16252 9466
rect 16408 9466 16436 10066
rect 16500 9654 16528 10084
rect 16580 10066 16632 10072
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 16408 9438 16620 9466
rect 16040 9178 16068 9386
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 14844 8090 14872 8978
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15396 8634 15424 9046
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 15212 8022 15240 8366
rect 16040 8022 16068 9114
rect 16132 9081 16160 9438
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16224 9178 16252 9318
rect 16592 9178 16620 9438
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16684 9081 16712 9386
rect 16118 9072 16174 9081
rect 16118 9007 16174 9016
rect 16670 9072 16726 9081
rect 16670 9007 16726 9016
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16224 8498 16252 8910
rect 16684 8566 16712 9007
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16224 8362 16252 8434
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 15476 8016 15528 8022
rect 16028 8016 16080 8022
rect 15476 7958 15528 7964
rect 15948 7964 16028 7970
rect 15948 7958 16080 7964
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15396 7546 15424 7822
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 14922 7440 14978 7449
rect 14922 7375 14924 7384
rect 14976 7375 14978 7384
rect 15200 7404 15252 7410
rect 14924 7346 14976 7352
rect 15200 7346 15252 7352
rect 15212 7154 15240 7346
rect 15488 7206 15516 7958
rect 15948 7942 16068 7958
rect 15948 7410 15976 7942
rect 16132 7818 16160 8298
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 15120 7126 15240 7154
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15120 6730 15148 7126
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14660 6446 14780 6474
rect 14660 5817 14688 6446
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14646 5808 14702 5817
rect 14556 5772 14608 5778
rect 14646 5743 14702 5752
rect 14556 5714 14608 5720
rect 14568 5370 14596 5714
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 14200 4282 14228 4626
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14384 4214 14412 5170
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10980 2825 11008 2858
rect 10966 2816 11022 2825
rect 10966 2751 11022 2760
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 10704 1006 10824 1034
rect 10796 480 10824 1006
rect 11808 480 11836 2246
rect 12912 480 12940 3334
rect 13910 3224 13966 3233
rect 13910 3159 13966 3168
rect 13726 2952 13782 2961
rect 13726 2887 13728 2896
rect 13780 2887 13782 2896
rect 13728 2858 13780 2864
rect 13924 480 13952 3159
rect 14568 3097 14596 5306
rect 14752 3942 14780 6258
rect 14844 5914 14872 6598
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 15304 5846 15332 7142
rect 15488 6934 15516 7142
rect 16132 6934 16160 7754
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15396 6322 15424 6734
rect 15488 6458 15516 6870
rect 16868 6866 16896 10406
rect 16960 10198 16988 10542
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15488 5778 15516 6394
rect 16868 5914 16896 6802
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15488 5370 15516 5714
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 16776 5030 16804 5646
rect 17052 5250 17080 12396
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17144 11286 17172 12242
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17236 10792 17264 15807
rect 17972 15706 18000 16646
rect 18064 16250 18092 17002
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18340 16726 18368 16934
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18144 16516 18196 16522
rect 18144 16458 18196 16464
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 18064 15994 18092 16186
rect 18156 16114 18184 16458
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 18064 15978 18184 15994
rect 18064 15972 18196 15978
rect 18064 15966 18144 15972
rect 18144 15914 18196 15920
rect 18340 15706 18368 16662
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17512 15162 17540 15574
rect 17868 15496 17920 15502
rect 17920 15444 18000 15450
rect 17868 15438 18000 15444
rect 17880 15422 18000 15438
rect 17972 15162 18000 15422
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 17604 14482 17632 14758
rect 18432 14550 18460 14758
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17500 12300 17552 12306
rect 17604 12288 17632 14418
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17972 13394 18000 14350
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 13462 18092 13806
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 17972 12986 18000 13330
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17552 12260 17632 12288
rect 17500 12242 17552 12248
rect 17512 11830 17540 12242
rect 17684 12164 17736 12170
rect 17684 12106 17736 12112
rect 17500 11824 17552 11830
rect 17500 11766 17552 11772
rect 17512 11218 17540 11766
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17144 10764 17264 10792
rect 17144 9194 17172 10764
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17236 10130 17264 10610
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17236 9654 17264 10066
rect 17328 9722 17356 10134
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17144 9166 17264 9194
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 17144 8634 17172 8978
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17052 5234 17172 5250
rect 17052 5228 17184 5234
rect 17052 5222 17132 5228
rect 17132 5170 17184 5176
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 15764 4690 15792 4966
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15764 4282 15792 4626
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15948 4049 15976 4422
rect 16120 4208 16172 4214
rect 16120 4150 16172 4156
rect 15934 4040 15990 4049
rect 15934 3975 15990 3984
rect 14740 3936 14792 3942
rect 14924 3936 14976 3942
rect 14740 3878 14792 3884
rect 14922 3904 14924 3913
rect 16132 3913 16160 4150
rect 14976 3904 14978 3913
rect 14922 3839 14978 3848
rect 15934 3904 15990 3913
rect 15934 3839 15990 3848
rect 16118 3904 16174 3913
rect 16118 3839 16174 3848
rect 14830 3632 14886 3641
rect 14830 3567 14886 3576
rect 14554 3088 14610 3097
rect 14554 3023 14610 3032
rect 14844 1850 14872 3567
rect 15384 3392 15436 3398
rect 15382 3360 15384 3369
rect 15436 3360 15438 3369
rect 14956 3292 15252 3312
rect 15382 3295 15438 3304
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14844 1822 14964 1850
rect 14936 480 14964 1822
rect 15948 480 15976 3839
rect 16776 2650 16804 4966
rect 17144 3505 17172 5170
rect 17236 3641 17264 9166
rect 17696 7954 17724 12106
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 18064 10130 18092 11018
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17972 9586 18000 9998
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17880 8906 17908 9386
rect 17972 9178 18000 9522
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 18524 9110 18552 23598
rect 20626 23559 20682 23568
rect 22190 23624 22192 23633
rect 22244 23624 22246 23633
rect 22190 23559 22246 23568
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18800 15706 18828 16730
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 18880 15972 18932 15978
rect 18880 15914 18932 15920
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18892 15434 18920 15914
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 18972 15632 19024 15638
rect 18972 15574 19024 15580
rect 18880 15428 18932 15434
rect 18880 15370 18932 15376
rect 18892 15065 18920 15370
rect 18878 15056 18934 15065
rect 18878 14991 18934 15000
rect 18984 14618 19012 15574
rect 19076 14890 19104 15846
rect 19168 15638 19196 15914
rect 19444 15910 19472 16594
rect 19432 15904 19484 15910
rect 19430 15872 19432 15881
rect 19484 15872 19486 15881
rect 19430 15807 19486 15816
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19156 15632 19208 15638
rect 19156 15574 19208 15580
rect 19168 15162 19196 15574
rect 19524 15428 19576 15434
rect 19524 15370 19576 15376
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 19064 14884 19116 14890
rect 19064 14826 19116 14832
rect 18972 14612 19024 14618
rect 18972 14554 19024 14560
rect 19076 14074 19104 14826
rect 19168 14618 19196 15098
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19168 14074 19196 14554
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19352 14074 19380 14486
rect 19536 14385 19564 15370
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19996 15162 20024 15302
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 20640 15042 20668 23559
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21652 19378 21680 23462
rect 23478 23080 23534 23089
rect 23478 23015 23534 23024
rect 23492 19417 23520 23015
rect 23478 19408 23534 19417
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 21640 19372 21692 19378
rect 23478 19343 23534 19352
rect 21640 19314 21692 19320
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 20364 15014 20760 15042
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19996 14550 20024 14962
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19522 14376 19578 14385
rect 19522 14311 19578 14320
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19246 13832 19302 13841
rect 18880 13796 18932 13802
rect 19246 13767 19302 13776
rect 18880 13738 18932 13744
rect 18892 13462 18920 13738
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18788 12980 18840 12986
rect 18892 12968 18920 13398
rect 19260 12986 19288 13767
rect 19536 13530 19564 14311
rect 19996 13938 20024 14486
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19996 13530 20024 13874
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 18840 12940 18920 12968
rect 18788 12922 18840 12928
rect 18892 12374 18920 12940
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19536 12850 19564 13466
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 18880 12368 18932 12374
rect 18786 12336 18842 12345
rect 18880 12310 18932 12316
rect 18786 12271 18788 12280
rect 18840 12271 18842 12280
rect 18788 12242 18840 12248
rect 18800 11354 18828 12242
rect 18892 11898 18920 12310
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 18892 11626 18920 11834
rect 18880 11620 18932 11626
rect 18880 11562 18932 11568
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18892 10198 18920 11562
rect 19536 11218 19564 12038
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19536 10810 19564 11154
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 18880 10192 18932 10198
rect 18880 10134 18932 10140
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18616 9178 18644 10066
rect 18892 9586 18920 10134
rect 18984 9722 19012 10542
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 18972 9716 19024 9722
rect 18972 9658 19024 9664
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 19076 9110 19104 10406
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 19996 9450 20024 9590
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17880 8022 17908 8842
rect 18524 8634 18552 9046
rect 18786 8936 18842 8945
rect 18786 8871 18842 8880
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18800 8498 18828 8871
rect 19076 8634 19104 9046
rect 19536 8838 19564 9386
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 19536 8090 19564 8774
rect 19996 8650 20024 9386
rect 20180 9110 20208 9522
rect 20168 9104 20220 9110
rect 20168 9046 20220 9052
rect 19996 8634 20116 8650
rect 19984 8628 20116 8634
rect 20036 8622 20116 8628
rect 19984 8570 20036 8576
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 17868 8016 17920 8022
rect 19996 7970 20024 8434
rect 20088 8362 20116 8622
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 17868 7958 17920 7964
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17696 7546 17724 7890
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17880 7410 17908 7958
rect 19904 7942 20024 7970
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18892 7410 18920 7686
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 17880 6934 17908 7346
rect 17408 6928 17460 6934
rect 17408 6870 17460 6876
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 18788 6928 18840 6934
rect 18788 6870 18840 6876
rect 17420 6458 17448 6870
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17788 6254 17816 6598
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17788 6118 17816 6190
rect 17972 6186 18000 6598
rect 17960 6180 18012 6186
rect 17880 6140 17960 6168
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17788 5846 17816 6054
rect 17776 5840 17828 5846
rect 17590 5808 17646 5817
rect 17776 5782 17828 5788
rect 17590 5743 17646 5752
rect 17604 4690 17632 5743
rect 17788 5658 17816 5782
rect 17696 5630 17816 5658
rect 17696 5234 17724 5630
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17788 5370 17816 5510
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17880 4826 17908 6140
rect 17960 6122 18012 6128
rect 18708 5574 18736 6734
rect 18800 6458 18828 6870
rect 18892 6798 18920 7346
rect 18984 7313 19012 7754
rect 19904 7750 19932 7942
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19892 7744 19944 7750
rect 19890 7712 19892 7721
rect 19944 7712 19946 7721
rect 19890 7647 19946 7656
rect 18970 7304 19026 7313
rect 18970 7239 18972 7248
rect 19024 7239 19026 7248
rect 19524 7268 19576 7274
rect 18972 7210 19024 7216
rect 19524 7210 19576 7216
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18892 6322 18920 6734
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19248 5840 19300 5846
rect 19248 5782 19300 5788
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 19260 5370 19288 5782
rect 19352 5710 19380 6258
rect 19444 6254 19472 6598
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 5370 19380 5646
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19444 5234 19472 6190
rect 19536 5710 19564 7210
rect 19996 7206 20024 7822
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 19812 6186 19840 6326
rect 19800 6180 19852 6186
rect 19800 6122 19852 6128
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17592 4684 17644 4690
rect 17592 4626 17644 4632
rect 17604 4282 17632 4626
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17222 3632 17278 3641
rect 17222 3567 17278 3576
rect 17604 3505 17632 4218
rect 19996 4185 20024 7142
rect 18970 4176 19026 4185
rect 18970 4111 19026 4120
rect 19982 4176 20038 4185
rect 19982 4111 20038 4120
rect 18050 4040 18106 4049
rect 18050 3975 18106 3984
rect 17958 3768 18014 3777
rect 17958 3703 18014 3712
rect 17130 3496 17186 3505
rect 17130 3431 17186 3440
rect 17590 3496 17646 3505
rect 17590 3431 17646 3440
rect 17972 2990 18000 3703
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17052 2310 17080 2450
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 17052 480 17080 2246
rect 18064 480 18092 3975
rect 18984 2650 19012 4111
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19444 2825 19472 4014
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20076 3120 20128 3126
rect 20076 3062 20128 3068
rect 19430 2816 19486 2825
rect 19430 2751 19486 2760
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 19064 2372 19116 2378
rect 19064 2314 19116 2320
rect 19076 480 19104 2314
rect 20088 480 20116 3062
rect 20272 2650 20300 12854
rect 20364 3233 20392 15014
rect 20732 14958 20760 15014
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 21192 14550 21220 14826
rect 21180 14544 21232 14550
rect 21180 14486 21232 14492
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 20904 13864 20956 13870
rect 21008 13841 21036 14350
rect 21192 14074 21220 14486
rect 21272 14408 21324 14414
rect 21270 14376 21272 14385
rect 21324 14376 21326 14385
rect 21270 14311 21326 14320
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 20904 13806 20956 13812
rect 20994 13832 21050 13841
rect 20720 13796 20772 13802
rect 20720 13738 20772 13744
rect 20732 13462 20760 13738
rect 20720 13456 20772 13462
rect 20720 13398 20772 13404
rect 20916 12889 20944 13806
rect 20994 13767 21050 13776
rect 20996 13388 21048 13394
rect 20996 13330 21048 13336
rect 21008 12986 21036 13330
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20626 12880 20682 12889
rect 20626 12815 20628 12824
rect 20680 12815 20682 12824
rect 20902 12880 20958 12889
rect 20902 12815 20958 12824
rect 20628 12786 20680 12792
rect 21008 12714 21036 12922
rect 21376 12782 21404 19314
rect 23570 15056 23626 15065
rect 23570 14991 23626 15000
rect 23584 14958 23612 14991
rect 23572 14952 23624 14958
rect 23572 14894 23624 14900
rect 21548 13864 21600 13870
rect 21546 13832 21548 13841
rect 21600 13832 21602 13841
rect 21546 13767 21602 13776
rect 22466 12880 22522 12889
rect 22466 12815 22522 12824
rect 22480 12782 22508 12815
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 20996 12708 21048 12714
rect 20996 12650 21048 12656
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20916 11558 20944 12378
rect 21192 12322 21220 12582
rect 21008 12294 21220 12322
rect 21008 12238 21036 12294
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21008 11898 21036 12174
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21100 11626 21128 12174
rect 21376 11642 21404 12718
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22468 12300 22520 12306
rect 22468 12242 22520 12248
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 21088 11620 21140 11626
rect 21088 11562 21140 11568
rect 21192 11614 21404 11642
rect 22100 11620 22152 11626
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20916 11286 20944 11494
rect 20904 11280 20956 11286
rect 20904 11222 20956 11228
rect 20442 11112 20498 11121
rect 20442 11047 20498 11056
rect 20456 10674 20484 11047
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20456 10266 20484 10610
rect 20548 10538 20576 10746
rect 21100 10674 21128 11562
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20536 10532 20588 10538
rect 20536 10474 20588 10480
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20812 10192 20864 10198
rect 20812 10134 20864 10140
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20732 9722 20760 9998
rect 20824 9926 20852 10134
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20732 9586 20760 9658
rect 20824 9654 20852 9862
rect 20812 9648 20864 9654
rect 20812 9590 20864 9596
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20824 8430 20852 9590
rect 21088 9104 21140 9110
rect 21088 9046 21140 9052
rect 20996 8968 21048 8974
rect 20994 8936 20996 8945
rect 21048 8936 21050 8945
rect 20994 8871 21050 8880
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 21008 8090 21036 8871
rect 21100 8566 21128 9046
rect 21088 8560 21140 8566
rect 21088 8502 21140 8508
rect 21192 8106 21220 11614
rect 22100 11562 22152 11568
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21376 11354 21404 11494
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21376 10606 21404 11290
rect 22112 11286 22140 11562
rect 21916 11280 21968 11286
rect 21916 11222 21968 11228
rect 22100 11280 22152 11286
rect 22100 11222 22152 11228
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21468 10810 21496 11086
rect 21928 10810 21956 11222
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21916 10804 21968 10810
rect 21916 10746 21968 10752
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 22020 10266 22048 10542
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 22112 10130 22140 11222
rect 22204 11121 22232 12038
rect 22480 11558 22508 12242
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22480 11257 22508 11494
rect 22466 11248 22522 11257
rect 22466 11183 22522 11192
rect 22190 11112 22246 11121
rect 22190 11047 22246 11056
rect 22100 10124 22152 10130
rect 22100 10066 22152 10072
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 21744 9586 21772 9998
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21732 9580 21784 9586
rect 21732 9522 21784 9528
rect 21284 8974 21312 9522
rect 21548 9444 21600 9450
rect 21548 9386 21600 9392
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21284 8498 21312 8910
rect 21560 8634 21588 9386
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21100 8078 21220 8106
rect 21652 8090 21680 8366
rect 21640 8084 21692 8090
rect 20534 7848 20590 7857
rect 20534 7783 20590 7792
rect 20548 7546 20576 7783
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20994 7304 21050 7313
rect 20994 7239 21050 7248
rect 21008 6866 21036 7239
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20916 5846 20944 6734
rect 21008 6458 21036 6802
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 20904 5840 20956 5846
rect 20904 5782 20956 5788
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20350 3224 20406 3233
rect 20350 3159 20406 3168
rect 20456 3097 20484 3878
rect 21100 3369 21128 8078
rect 21640 8026 21692 8032
rect 21744 7954 21772 9522
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21732 7948 21784 7954
rect 21732 7890 21784 7896
rect 21192 7546 21220 7890
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21284 3602 21312 7686
rect 22664 6361 22692 12582
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 23124 9722 23152 10066
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23112 9716 23164 9722
rect 23112 9658 23164 9664
rect 23400 8514 23428 9862
rect 23570 9072 23626 9081
rect 23570 9007 23572 9016
rect 23624 9007 23626 9016
rect 23572 8978 23624 8984
rect 23584 8634 23612 8978
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23400 8486 23520 8514
rect 23492 8430 23520 8486
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23478 7712 23534 7721
rect 23478 7647 23534 7656
rect 23492 7546 23520 7647
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 22834 7440 22890 7449
rect 22834 7375 22890 7384
rect 22650 6352 22706 6361
rect 22650 6287 22706 6296
rect 21730 3632 21786 3641
rect 21272 3596 21324 3602
rect 21730 3567 21786 3576
rect 22100 3596 22152 3602
rect 21272 3538 21324 3544
rect 21638 3496 21694 3505
rect 21638 3431 21694 3440
rect 21086 3360 21142 3369
rect 21086 3295 21142 3304
rect 20442 3088 20498 3097
rect 20442 3023 20498 3032
rect 21652 2802 21680 3431
rect 21744 3194 21772 3567
rect 22100 3538 22152 3544
rect 21822 3496 21878 3505
rect 21822 3431 21824 3440
rect 21876 3431 21878 3440
rect 21824 3402 21876 3408
rect 22112 3194 22140 3538
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 21744 2990 21772 3130
rect 22190 3088 22246 3097
rect 22190 3023 22246 3032
rect 21732 2984 21784 2990
rect 21732 2926 21784 2932
rect 21914 2816 21970 2825
rect 21652 2774 21772 2802
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 21744 2514 21772 2774
rect 21914 2751 21970 2760
rect 21928 2650 21956 2751
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 21732 2508 21784 2514
rect 21732 2450 21784 2456
rect 21180 2372 21232 2378
rect 21180 2314 21232 2320
rect 21192 480 21220 2314
rect 22204 480 22232 3023
rect 22848 2514 22876 7375
rect 23478 5672 23534 5681
rect 23478 5607 23534 5616
rect 23492 5370 23520 5607
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 23216 480 23244 2790
rect 23676 2514 23704 27231
rect 23846 25936 23902 25945
rect 23846 25871 23902 25880
rect 23754 24576 23810 24585
rect 23754 24511 23810 24520
rect 23768 18873 23796 24511
rect 23860 19961 23888 25871
rect 24228 24313 24256 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24214 24304 24270 24313
rect 24214 24239 24270 24248
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 25332 22001 25360 27520
rect 26344 24313 26372 27520
rect 26330 24304 26386 24313
rect 26330 24239 26386 24248
rect 27356 23769 27384 27520
rect 27342 23760 27398 23769
rect 27342 23695 27398 23704
rect 25318 21992 25374 22001
rect 25318 21927 25374 21936
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24674 21720 24730 21729
rect 24674 21655 24730 21664
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24122 20360 24178 20369
rect 24122 20295 24178 20304
rect 23846 19952 23902 19961
rect 23846 19887 23902 19896
rect 23754 18864 23810 18873
rect 23754 18799 23810 18808
rect 24136 17513 24164 20295
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24688 18737 24716 21655
rect 24766 18864 24822 18873
rect 24766 18799 24822 18808
rect 24674 18728 24730 18737
rect 24674 18663 24730 18672
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24122 17504 24178 17513
rect 24122 17439 24178 17448
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24780 17105 24808 18799
rect 24766 17096 24822 17105
rect 24766 17031 24822 17040
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24216 14884 24268 14890
rect 24216 14826 24268 14832
rect 24124 11212 24176 11218
rect 24124 11154 24176 11160
rect 24136 10606 24164 11154
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24228 4690 24256 14826
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24766 13288 24822 13297
rect 24766 13223 24822 13232
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24780 12442 24808 13223
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24766 11928 24822 11937
rect 24766 11863 24822 11872
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10606 24716 10950
rect 24780 10810 24808 11863
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24308 10600 24360 10606
rect 24306 10568 24308 10577
rect 24676 10600 24728 10606
rect 24360 10568 24362 10577
rect 24676 10542 24728 10548
rect 24766 10568 24822 10577
rect 24306 10503 24362 10512
rect 24766 10503 24822 10512
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24780 9654 24808 10503
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24596 9178 24624 9454
rect 24584 9172 24636 9178
rect 24584 9114 24636 9120
rect 24766 9072 24822 9081
rect 24766 9007 24822 9016
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24584 7948 24636 7954
rect 24584 7890 24636 7896
rect 24596 7857 24624 7890
rect 24582 7848 24638 7857
rect 24582 7783 24638 7792
rect 24688 7721 24716 8230
rect 24780 8090 24808 9007
rect 24768 8084 24820 8090
rect 24768 8026 24820 8032
rect 25412 7948 25464 7954
rect 25412 7890 25464 7896
rect 24674 7712 24730 7721
rect 24289 7644 24585 7664
rect 24674 7647 24730 7656
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 25424 7546 25452 7890
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24582 6352 24638 6361
rect 24582 6287 24638 6296
rect 24596 6254 24624 6287
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24216 4684 24268 4690
rect 24216 4626 24268 4632
rect 24228 4282 24256 4626
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24216 4276 24268 4282
rect 24216 4218 24268 4224
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24308 2984 24360 2990
rect 24306 2952 24308 2961
rect 24360 2952 24362 2961
rect 24306 2887 24362 2896
rect 24492 2848 24544 2854
rect 24214 2816 24270 2825
rect 24214 2751 24270 2760
rect 24490 2816 24492 2825
rect 24544 2816 24546 2825
rect 24490 2751 24546 2760
rect 23664 2508 23716 2514
rect 23664 2450 23716 2456
rect 24228 480 24256 2751
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 785 24716 7278
rect 24768 6384 24820 6390
rect 24766 6352 24768 6361
rect 24820 6352 24822 6361
rect 24766 6287 24822 6296
rect 25136 5024 25188 5030
rect 25134 4992 25136 5001
rect 25188 4992 25190 5001
rect 25134 4927 25190 4936
rect 27342 4992 27398 5001
rect 27342 4927 27398 4936
rect 24766 4856 24822 4865
rect 24766 4791 24768 4800
rect 24820 4791 24822 4800
rect 24768 4762 24820 4768
rect 26330 2816 26386 2825
rect 26330 2751 26386 2760
rect 25320 2372 25372 2378
rect 25320 2314 25372 2320
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 24780 2145 24808 2246
rect 24766 2136 24822 2145
rect 24766 2071 24822 2080
rect 24674 776 24730 785
rect 24674 711 24730 720
rect 25332 480 25360 2314
rect 26344 480 26372 2751
rect 27356 480 27384 4927
rect 478 0 534 480
rect 1490 0 1546 480
rect 2502 0 2558 480
rect 3514 0 3570 480
rect 4618 0 4674 480
rect 5630 0 5686 480
rect 6642 0 6698 480
rect 7654 0 7710 480
rect 8758 0 8814 480
rect 9770 0 9826 480
rect 10782 0 10838 480
rect 11794 0 11850 480
rect 12898 0 12954 480
rect 13910 0 13966 480
rect 14922 0 14978 480
rect 15934 0 15990 480
rect 17038 0 17094 480
rect 18050 0 18106 480
rect 19062 0 19118 480
rect 20074 0 20130 480
rect 21178 0 21234 480
rect 22190 0 22246 480
rect 23202 0 23258 480
rect 24214 0 24270 480
rect 25318 0 25374 480
rect 26330 0 26386 480
rect 27342 0 27398 480
<< via2 >>
rect 2686 24132 2742 24168
rect 2686 24112 2688 24132
rect 2688 24112 2740 24132
rect 2740 24112 2742 24132
rect 4066 26424 4122 26480
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5446 24248 5502 24304
rect 2686 23568 2742 23624
rect 5354 23432 5410 23488
rect 3422 23296 3478 23352
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5078 22344 5134 22400
rect 8574 24812 8630 24848
rect 8574 24792 8576 24812
rect 8576 24792 8628 24812
rect 8628 24792 8630 24812
rect 7102 23468 7104 23488
rect 7104 23468 7156 23488
rect 7156 23468 7158 23488
rect 7102 23432 7158 23468
rect 5998 21836 6000 21856
rect 6000 21836 6052 21856
rect 6052 21836 6054 21856
rect 5998 21800 6054 21836
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 6182 21004 6238 21040
rect 6182 20984 6184 21004
rect 6184 20984 6236 21004
rect 6236 20984 6238 21004
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5722 20340 5724 20360
rect 5724 20340 5776 20360
rect 5776 20340 5778 20360
rect 5722 20304 5778 20340
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5722 19252 5724 19272
rect 5724 19252 5776 19272
rect 5776 19252 5778 19272
rect 5078 18808 5134 18864
rect 5722 19216 5778 19252
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5354 17584 5410 17640
rect 4066 17040 4122 17096
rect 3422 14864 3478 14920
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 6274 17720 6330 17776
rect 4342 16632 4398 16688
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 6274 16224 6330 16280
rect 5262 15988 5264 16008
rect 5264 15988 5316 16008
rect 5316 15988 5318 16008
rect 5262 15952 5318 15988
rect 4250 15000 4306 15056
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5538 14864 5594 14920
rect 4066 13912 4122 13968
rect 2502 13640 2558 13696
rect 4342 13640 4398 13696
rect 2870 12708 2926 12744
rect 2870 12688 2872 12708
rect 2872 12688 2924 12708
rect 2924 12688 2926 12708
rect 3606 12280 3662 12336
rect 2594 12144 2650 12200
rect 2226 11600 2282 11656
rect 2594 7656 2650 7712
rect 2686 3576 2742 3632
rect 1582 2644 1638 2680
rect 1582 2624 1584 2644
rect 1584 2624 1636 2644
rect 1636 2624 1638 2644
rect 1490 2488 1546 2544
rect 478 1808 534 1864
rect 1398 1808 1454 1864
rect 6458 18128 6514 18184
rect 7286 20168 7342 20224
rect 6550 17584 6606 17640
rect 6458 15816 6514 15872
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 3330 10784 3386 10840
rect 3146 10124 3202 10160
rect 3146 10104 3148 10124
rect 3148 10104 3200 10124
rect 3200 10104 3202 10124
rect 3698 10684 3700 10704
rect 3700 10684 3752 10704
rect 3752 10684 3754 10704
rect 3698 10648 3754 10684
rect 4066 10412 4068 10432
rect 4068 10412 4120 10432
rect 4120 10412 4122 10432
rect 4066 10376 4122 10412
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5998 10648 6054 10704
rect 5538 10376 5594 10432
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5446 9288 5502 9344
rect 3882 6840 3938 6896
rect 5170 7948 5226 7984
rect 5170 7928 5172 7948
rect 5172 7928 5224 7948
rect 5224 7928 5226 7948
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 6642 13640 6698 13696
rect 6550 12044 6552 12064
rect 6552 12044 6604 12064
rect 6604 12044 6606 12064
rect 6550 12008 6606 12044
rect 5998 8608 6054 8664
rect 5446 7384 5502 7440
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 6274 7928 6330 7984
rect 6642 10648 6698 10704
rect 6642 10412 6644 10432
rect 6644 10412 6696 10432
rect 6696 10412 6698 10432
rect 6642 10376 6698 10412
rect 8482 23840 8538 23896
rect 8206 21292 8208 21312
rect 8208 21292 8260 21312
rect 8260 21292 8262 21312
rect 8206 21256 8262 21292
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 9678 24112 9734 24168
rect 9862 24132 9918 24168
rect 9862 24112 9864 24132
rect 9864 24112 9916 24132
rect 9916 24112 9918 24132
rect 9126 22380 9128 22400
rect 9128 22380 9180 22400
rect 9180 22380 9182 22400
rect 9126 22344 9182 22380
rect 9310 21936 9366 21992
rect 9034 21800 9090 21856
rect 8850 20304 8906 20360
rect 8666 17212 8668 17232
rect 8668 17212 8720 17232
rect 8720 17212 8722 17232
rect 8666 17176 8722 17212
rect 8758 15852 8760 15872
rect 8760 15852 8812 15872
rect 8812 15852 8814 15872
rect 7194 12300 7250 12336
rect 7194 12280 7196 12300
rect 7196 12280 7248 12300
rect 7248 12280 7250 12300
rect 6826 9560 6882 9616
rect 7010 9324 7012 9344
rect 7012 9324 7064 9344
rect 7064 9324 7066 9344
rect 7010 9288 7066 9324
rect 6458 8200 6514 8256
rect 6366 7384 6422 7440
rect 5446 6296 5502 6352
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 6918 6860 6974 6896
rect 6918 6840 6920 6860
rect 6920 6840 6972 6860
rect 6972 6840 6974 6860
rect 7194 6840 7250 6896
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 4066 4528 4122 4584
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5446 3848 5502 3904
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 3514 2760 3570 2816
rect 2870 1536 2926 1592
rect 4618 2488 4674 2544
rect 6366 2796 6368 2816
rect 6368 2796 6420 2816
rect 6420 2796 6422 2816
rect 6366 2760 6422 2796
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 7562 12708 7618 12744
rect 7562 12688 7564 12708
rect 7564 12688 7616 12708
rect 7616 12688 7618 12708
rect 7838 12688 7894 12744
rect 8758 15816 8814 15852
rect 8206 14864 8262 14920
rect 7930 11348 7986 11384
rect 7930 11328 7932 11348
rect 7932 11328 7984 11348
rect 7984 11328 7986 11348
rect 7562 9868 7564 9888
rect 7564 9868 7616 9888
rect 7616 9868 7618 9888
rect 7562 9832 7618 9868
rect 7930 6296 7986 6352
rect 7838 5888 7894 5944
rect 7194 2624 7250 2680
rect 7746 3168 7802 3224
rect 8114 12824 8170 12880
rect 8298 13640 8354 13696
rect 8482 12960 8538 13016
rect 8758 12164 8814 12200
rect 8758 12144 8760 12164
rect 8760 12144 8812 12164
rect 8812 12144 8814 12164
rect 8574 12008 8630 12064
rect 8482 11328 8538 11384
rect 8850 11192 8906 11248
rect 8114 5092 8170 5128
rect 8114 5072 8116 5092
rect 8116 5072 8168 5092
rect 8168 5072 8170 5092
rect 8666 8628 8722 8664
rect 8666 8608 8668 8628
rect 8668 8608 8720 8628
rect 8720 8608 8722 8628
rect 8758 7828 8760 7848
rect 8760 7828 8812 7848
rect 8812 7828 8814 7848
rect 8758 7792 8814 7828
rect 8666 6160 8722 6216
rect 8482 3168 8538 3224
rect 8022 2488 8078 2544
rect 9402 21256 9458 21312
rect 9494 17584 9550 17640
rect 9678 15000 9734 15056
rect 9034 14728 9090 14784
rect 9126 12144 9182 12200
rect 9494 12688 9550 12744
rect 9586 12280 9642 12336
rect 9586 11192 9642 11248
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 9862 19216 9918 19272
rect 10046 19352 10102 19408
rect 10046 18128 10102 18184
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 9954 14184 10010 14240
rect 9770 11328 9826 11384
rect 9494 9696 9550 9752
rect 9310 9560 9366 9616
rect 9678 10412 9680 10432
rect 9680 10412 9732 10432
rect 9732 10412 9734 10432
rect 9678 10376 9734 10412
rect 9678 10124 9734 10160
rect 9678 10104 9680 10124
rect 9680 10104 9732 10124
rect 9732 10104 9734 10124
rect 9862 10784 9918 10840
rect 9862 8200 9918 8256
rect 9770 7948 9826 7984
rect 9770 7928 9772 7948
rect 9772 7928 9824 7948
rect 9824 7928 9826 7948
rect 9586 7520 9642 7576
rect 9034 4120 9090 4176
rect 9862 5888 9918 5944
rect 9770 5072 9826 5128
rect 9862 3168 9918 3224
rect 9770 3032 9826 3088
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10690 16652 10746 16688
rect 10690 16632 10692 16652
rect 10692 16632 10744 16652
rect 10744 16632 10746 16652
rect 10230 16244 10286 16280
rect 10230 16224 10232 16244
rect 10232 16224 10284 16244
rect 10284 16224 10286 16244
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 12162 23860 12218 23896
rect 12162 23840 12164 23860
rect 12164 23840 12216 23860
rect 12216 23840 12218 23860
rect 10966 22516 10968 22536
rect 10968 22516 11020 22536
rect 11020 22516 11022 22536
rect 10966 22480 11022 22516
rect 11794 23704 11850 23760
rect 12714 24384 12770 24440
rect 12714 24248 12770 24304
rect 11334 21412 11390 21448
rect 11334 21392 11336 21412
rect 11336 21392 11388 21412
rect 11388 21392 11390 21412
rect 10966 20576 11022 20632
rect 11978 19896 12034 19952
rect 12806 20576 12862 20632
rect 11886 18672 11942 18728
rect 10506 15408 10562 15464
rect 10690 15272 10746 15328
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10782 14456 10838 14512
rect 10874 14184 10930 14240
rect 10690 13640 10746 13696
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 11978 16668 11980 16688
rect 11980 16668 12032 16688
rect 12032 16668 12034 16688
rect 11978 16632 12034 16668
rect 11242 15272 11298 15328
rect 11334 14900 11336 14920
rect 11336 14900 11388 14920
rect 11388 14900 11390 14920
rect 11334 14864 11390 14900
rect 12622 15408 12678 15464
rect 12530 13640 12586 13696
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10506 7420 10508 7440
rect 10508 7420 10560 7440
rect 10560 7420 10562 7440
rect 10506 7384 10562 7420
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10046 5752 10102 5808
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 11058 10648 11114 10704
rect 12438 12960 12494 13016
rect 11518 12300 11574 12336
rect 11518 12280 11520 12300
rect 11520 12280 11572 12300
rect 11572 12280 11574 12300
rect 10690 3984 10746 4040
rect 10046 3848 10102 3904
rect 10690 3848 10746 3904
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10138 3576 10194 3632
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 9862 2352 9918 2408
rect 11150 6860 11206 6896
rect 11150 6840 11152 6860
rect 11152 6840 11204 6860
rect 11204 6840 11206 6860
rect 11886 10512 11942 10568
rect 12162 9868 12164 9888
rect 12164 9868 12216 9888
rect 12216 9868 12218 9888
rect 12162 9832 12218 9868
rect 12438 9696 12494 9752
rect 11794 4120 11850 4176
rect 12346 9016 12402 9072
rect 12530 9580 12586 9616
rect 12530 9560 12532 9580
rect 12532 9560 12584 9580
rect 12584 9560 12586 9580
rect 12622 8336 12678 8392
rect 12438 7812 12494 7848
rect 12438 7792 12440 7812
rect 12440 7792 12492 7812
rect 12492 7792 12494 7812
rect 12530 7520 12586 7576
rect 13450 24792 13506 24848
rect 13726 23432 13782 23488
rect 13726 22480 13782 22536
rect 14094 23588 14150 23624
rect 14094 23568 14096 23588
rect 14096 23568 14148 23588
rect 14148 23568 14150 23588
rect 13174 18128 13230 18184
rect 13634 17720 13690 17776
rect 12990 16768 13046 16824
rect 13450 14864 13506 14920
rect 13082 14476 13138 14512
rect 13082 14456 13084 14476
rect 13084 14456 13136 14476
rect 13136 14456 13138 14476
rect 13450 12844 13506 12880
rect 13450 12824 13452 12844
rect 13452 12824 13504 12844
rect 13504 12824 13506 12844
rect 13818 12008 13874 12064
rect 12990 11056 13046 11112
rect 12898 10804 12954 10840
rect 12898 10784 12900 10804
rect 12900 10784 12952 10804
rect 12952 10784 12954 10804
rect 12898 9016 12954 9072
rect 13450 6160 13506 6216
rect 13634 5652 13636 5672
rect 13636 5652 13688 5672
rect 13688 5652 13690 5672
rect 13634 5616 13690 5652
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15934 23976 15990 24032
rect 15382 23604 15384 23624
rect 15384 23604 15436 23624
rect 15436 23604 15438 23624
rect 15382 23568 15438 23604
rect 15290 23432 15346 23488
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15382 22480 15438 22536
rect 14554 22344 14610 22400
rect 14094 17076 14096 17096
rect 14096 17076 14148 17096
rect 14148 17076 14150 17096
rect 14094 17040 14150 17076
rect 14462 15272 14518 15328
rect 14186 12688 14242 12744
rect 14186 11056 14242 11112
rect 14094 8336 14150 8392
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15014 21392 15070 21448
rect 15750 21392 15806 21448
rect 15290 20984 15346 21040
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14646 19896 14702 19952
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15198 19352 15254 19408
rect 15382 18828 15438 18864
rect 15382 18808 15384 18828
rect 15384 18808 15436 18828
rect 15436 18808 15438 18828
rect 15290 18672 15346 18728
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15198 16668 15200 16688
rect 15200 16668 15252 16688
rect 15252 16668 15254 16688
rect 15198 16632 15254 16668
rect 16026 19388 16028 19408
rect 16028 19388 16080 19408
rect 16080 19388 16082 19408
rect 16026 19352 16082 19388
rect 15382 17448 15438 17504
rect 15382 17176 15438 17232
rect 15566 16632 15622 16688
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14830 15952 14886 16008
rect 14830 15408 14886 15464
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14646 14184 14702 14240
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14646 10512 14702 10568
rect 15290 12144 15346 12200
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15290 10684 15292 10704
rect 15292 10684 15344 10704
rect 15344 10684 15346 10704
rect 15290 10648 15346 10684
rect 15842 12280 15898 12336
rect 15658 11600 15714 11656
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 16486 24132 16542 24168
rect 16486 24112 16488 24132
rect 16488 24112 16540 24132
rect 16540 24112 16542 24132
rect 16302 21936 16358 21992
rect 18234 24656 18290 24712
rect 18050 23976 18106 24032
rect 17130 23860 17186 23896
rect 17130 23840 17132 23860
rect 17132 23840 17184 23860
rect 17184 23840 17186 23860
rect 18050 23704 18106 23760
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 20074 24656 20130 24712
rect 19430 24520 19486 24576
rect 19062 23840 19118 23896
rect 19246 23860 19302 23896
rect 19246 23840 19248 23860
rect 19248 23840 19300 23860
rect 19300 23840 19302 23860
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20626 24248 20682 24304
rect 22190 24792 22246 24848
rect 22374 24248 22430 24304
rect 21270 23976 21326 24032
rect 21178 23840 21234 23896
rect 23662 27240 23718 27296
rect 23202 23976 23258 24032
rect 17038 21956 17094 21992
rect 17038 21936 17040 21956
rect 17040 21936 17092 21956
rect 17092 21936 17094 21956
rect 16854 21528 16910 21584
rect 15934 9560 15990 9616
rect 18418 22344 18474 22400
rect 17222 15816 17278 15872
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 16118 9016 16174 9072
rect 16670 9016 16726 9072
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14922 7404 14978 7440
rect 14922 7384 14924 7404
rect 14924 7384 14976 7404
rect 14976 7384 14978 7404
rect 14646 5752 14702 5808
rect 10966 2760 11022 2816
rect 13910 3168 13966 3224
rect 13726 2916 13782 2952
rect 13726 2896 13728 2916
rect 13728 2896 13780 2916
rect 13780 2896 13782 2916
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15934 3984 15990 4040
rect 14922 3884 14924 3904
rect 14924 3884 14976 3904
rect 14976 3884 14978 3904
rect 14922 3848 14978 3884
rect 15934 3848 15990 3904
rect 16118 3848 16174 3904
rect 14830 3576 14886 3632
rect 14554 3032 14610 3088
rect 15382 3340 15384 3360
rect 15384 3340 15436 3360
rect 15436 3340 15438 3360
rect 15382 3304 15438 3340
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 20626 23568 20682 23624
rect 22190 23604 22192 23624
rect 22192 23604 22244 23624
rect 22244 23604 22246 23624
rect 22190 23568 22246 23604
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 18878 15000 18934 15056
rect 19430 15852 19432 15872
rect 19432 15852 19484 15872
rect 19484 15852 19486 15872
rect 19430 15816 19486 15852
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 23478 23024 23534 23080
rect 23478 19352 23534 19408
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19522 14320 19578 14376
rect 19246 13776 19302 13832
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 18786 12300 18842 12336
rect 18786 12280 18788 12300
rect 18788 12280 18840 12300
rect 18840 12280 18842 12300
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 18786 8880 18842 8936
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 17590 5752 17646 5808
rect 19890 7692 19892 7712
rect 19892 7692 19944 7712
rect 19944 7692 19946 7712
rect 19890 7656 19946 7692
rect 18970 7268 19026 7304
rect 18970 7248 18972 7268
rect 18972 7248 19024 7268
rect 19024 7248 19026 7268
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 17222 3576 17278 3632
rect 18970 4120 19026 4176
rect 19982 4120 20038 4176
rect 18050 3984 18106 4040
rect 17958 3712 18014 3768
rect 17130 3440 17186 3496
rect 17590 3440 17646 3496
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19430 2760 19486 2816
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 21270 14356 21272 14376
rect 21272 14356 21324 14376
rect 21324 14356 21326 14376
rect 21270 14320 21326 14356
rect 20994 13776 21050 13832
rect 20626 12844 20682 12880
rect 20626 12824 20628 12844
rect 20628 12824 20680 12844
rect 20680 12824 20682 12844
rect 20902 12824 20958 12880
rect 23570 15000 23626 15056
rect 21546 13812 21548 13832
rect 21548 13812 21600 13832
rect 21600 13812 21602 13832
rect 21546 13776 21602 13812
rect 22466 12824 22522 12880
rect 20442 11056 20498 11112
rect 20994 8916 20996 8936
rect 20996 8916 21048 8936
rect 21048 8916 21050 8936
rect 20994 8880 21050 8916
rect 22466 11192 22522 11248
rect 22190 11056 22246 11112
rect 20534 7792 20590 7848
rect 20994 7248 21050 7304
rect 20350 3168 20406 3224
rect 23570 9036 23626 9072
rect 23570 9016 23572 9036
rect 23572 9016 23624 9036
rect 23624 9016 23626 9036
rect 23478 7656 23534 7712
rect 22834 7384 22890 7440
rect 22650 6296 22706 6352
rect 21730 3576 21786 3632
rect 21638 3440 21694 3496
rect 21086 3304 21142 3360
rect 20442 3032 20498 3088
rect 21822 3460 21878 3496
rect 21822 3440 21824 3460
rect 21824 3440 21876 3460
rect 21876 3440 21878 3460
rect 22190 3032 22246 3088
rect 21914 2760 21970 2816
rect 23478 5616 23534 5672
rect 23846 25880 23902 25936
rect 23754 24520 23810 24576
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24214 24248 24270 24304
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 26330 24248 26386 24304
rect 27342 23704 27398 23760
rect 25318 21936 25374 21992
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24674 21664 24730 21720
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24122 20304 24178 20360
rect 23846 19896 23902 19952
rect 23754 18808 23810 18864
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24766 18808 24822 18864
rect 24674 18672 24730 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24122 17448 24178 17504
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24766 17040 24822 17096
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24766 13232 24822 13288
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24766 11872 24822 11928
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24306 10548 24308 10568
rect 24308 10548 24360 10568
rect 24360 10548 24362 10568
rect 24306 10512 24362 10548
rect 24766 10512 24822 10568
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24766 9016 24822 9072
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24582 7792 24638 7848
rect 24674 7656 24730 7712
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24582 6296 24638 6352
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24306 2932 24308 2952
rect 24308 2932 24360 2952
rect 24360 2932 24362 2952
rect 24306 2896 24362 2932
rect 24214 2760 24270 2816
rect 24490 2796 24492 2816
rect 24492 2796 24544 2816
rect 24544 2796 24546 2816
rect 24490 2760 24546 2796
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24766 6332 24768 6352
rect 24768 6332 24820 6352
rect 24820 6332 24822 6352
rect 24766 6296 24822 6332
rect 25134 4972 25136 4992
rect 25136 4972 25188 4992
rect 25188 4972 25190 4992
rect 25134 4936 25190 4972
rect 27342 4936 27398 4992
rect 24766 4820 24822 4856
rect 24766 4800 24768 4820
rect 24768 4800 24820 4820
rect 24820 4800 24822 4820
rect 26330 2760 26386 2816
rect 24766 2080 24822 2136
rect 24674 720 24730 776
<< metal3 >>
rect 23657 27298 23723 27301
rect 27520 27298 28000 27328
rect 23657 27296 28000 27298
rect 23657 27240 23662 27296
rect 23718 27240 28000 27296
rect 23657 27238 28000 27240
rect 23657 27235 23723 27238
rect 27520 27208 28000 27238
rect 0 26482 480 26512
rect 4061 26482 4127 26485
rect 0 26480 4127 26482
rect 0 26424 4066 26480
rect 4122 26424 4127 26480
rect 0 26422 4127 26424
rect 0 26392 480 26422
rect 4061 26419 4127 26422
rect 23841 25938 23907 25941
rect 27520 25938 28000 25968
rect 23841 25936 28000 25938
rect 23841 25880 23846 25936
rect 23902 25880 28000 25936
rect 23841 25878 28000 25880
rect 23841 25875 23907 25878
rect 27520 25848 28000 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 8569 24850 8635 24853
rect 13445 24850 13511 24853
rect 22185 24850 22251 24853
rect 8569 24848 10794 24850
rect 8569 24792 8574 24848
rect 8630 24792 10794 24848
rect 8569 24790 10794 24792
rect 8569 24787 8635 24790
rect 10734 24578 10794 24790
rect 13445 24848 22251 24850
rect 13445 24792 13450 24848
rect 13506 24792 22190 24848
rect 22246 24792 22251 24848
rect 13445 24790 22251 24792
rect 13445 24787 13511 24790
rect 22185 24787 22251 24790
rect 18229 24714 18295 24717
rect 20069 24714 20135 24717
rect 18229 24712 20135 24714
rect 18229 24656 18234 24712
rect 18290 24656 20074 24712
rect 20130 24656 20135 24712
rect 18229 24654 20135 24656
rect 18229 24651 18295 24654
rect 20069 24651 20135 24654
rect 19425 24578 19491 24581
rect 10734 24576 19491 24578
rect 10734 24520 19430 24576
rect 19486 24520 19491 24576
rect 10734 24518 19491 24520
rect 19425 24515 19491 24518
rect 23749 24578 23815 24581
rect 27520 24578 28000 24608
rect 23749 24576 28000 24578
rect 23749 24520 23754 24576
rect 23810 24520 28000 24576
rect 23749 24518 28000 24520
rect 23749 24515 23815 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 27520 24488 28000 24518
rect 19610 24447 19930 24448
rect 12709 24442 12775 24445
rect 12709 24440 19442 24442
rect 12709 24384 12714 24440
rect 12770 24384 19442 24440
rect 12709 24382 19442 24384
rect 12709 24379 12775 24382
rect 5441 24306 5507 24309
rect 12709 24306 12775 24309
rect 5441 24304 12775 24306
rect 5441 24248 5446 24304
rect 5502 24248 12714 24304
rect 12770 24248 12775 24304
rect 5441 24246 12775 24248
rect 19382 24306 19442 24382
rect 20621 24306 20687 24309
rect 19382 24304 20687 24306
rect 19382 24248 20626 24304
rect 20682 24248 20687 24304
rect 19382 24246 20687 24248
rect 5441 24243 5507 24246
rect 12709 24243 12775 24246
rect 20621 24243 20687 24246
rect 22369 24306 22435 24309
rect 24209 24306 24275 24309
rect 26325 24306 26391 24309
rect 22369 24304 24275 24306
rect 22369 24248 22374 24304
rect 22430 24248 24214 24304
rect 24270 24248 24275 24304
rect 22369 24246 24275 24248
rect 22369 24243 22435 24246
rect 24209 24243 24275 24246
rect 24350 24304 26391 24306
rect 24350 24248 26330 24304
rect 26386 24248 26391 24304
rect 24350 24246 26391 24248
rect 2681 24170 2747 24173
rect 9673 24170 9739 24173
rect 9857 24170 9923 24173
rect 2681 24168 9923 24170
rect 2681 24112 2686 24168
rect 2742 24112 9678 24168
rect 9734 24112 9862 24168
rect 9918 24112 9923 24168
rect 2681 24110 9923 24112
rect 2681 24107 2747 24110
rect 9673 24107 9739 24110
rect 9857 24107 9923 24110
rect 16481 24170 16547 24173
rect 24350 24170 24410 24246
rect 26325 24243 26391 24246
rect 16481 24168 24410 24170
rect 16481 24112 16486 24168
rect 16542 24112 24410 24168
rect 16481 24110 24410 24112
rect 16481 24107 16547 24110
rect 15929 24034 15995 24037
rect 18045 24034 18111 24037
rect 15929 24032 18111 24034
rect 15929 23976 15934 24032
rect 15990 23976 18050 24032
rect 18106 23976 18111 24032
rect 15929 23974 18111 23976
rect 15929 23971 15995 23974
rect 18045 23971 18111 23974
rect 21265 24034 21331 24037
rect 23197 24034 23263 24037
rect 21265 24032 23263 24034
rect 21265 23976 21270 24032
rect 21326 23976 23202 24032
rect 23258 23976 23263 24032
rect 21265 23974 23263 23976
rect 21265 23971 21331 23974
rect 23197 23971 23263 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 8477 23898 8543 23901
rect 12157 23898 12223 23901
rect 8477 23896 12223 23898
rect 8477 23840 8482 23896
rect 8538 23840 12162 23896
rect 12218 23840 12223 23896
rect 8477 23838 12223 23840
rect 8477 23835 8543 23838
rect 12157 23835 12223 23838
rect 17125 23898 17191 23901
rect 19057 23898 19123 23901
rect 17125 23896 19123 23898
rect 17125 23840 17130 23896
rect 17186 23840 19062 23896
rect 19118 23840 19123 23896
rect 17125 23838 19123 23840
rect 17125 23835 17191 23838
rect 19057 23835 19123 23838
rect 19241 23898 19307 23901
rect 21173 23898 21239 23901
rect 19241 23896 21239 23898
rect 19241 23840 19246 23896
rect 19302 23840 21178 23896
rect 21234 23840 21239 23896
rect 19241 23838 21239 23840
rect 19241 23835 19307 23838
rect 21173 23835 21239 23838
rect 11789 23762 11855 23765
rect 18045 23762 18111 23765
rect 27337 23762 27403 23765
rect 11789 23760 18111 23762
rect 11789 23704 11794 23760
rect 11850 23704 18050 23760
rect 18106 23704 18111 23760
rect 11789 23702 18111 23704
rect 11789 23699 11855 23702
rect 18045 23699 18111 23702
rect 18278 23760 27403 23762
rect 18278 23704 27342 23760
rect 27398 23704 27403 23760
rect 18278 23702 27403 23704
rect 2681 23626 2747 23629
rect 14089 23626 14155 23629
rect 2681 23624 14155 23626
rect 2681 23568 2686 23624
rect 2742 23568 14094 23624
rect 14150 23568 14155 23624
rect 2681 23566 14155 23568
rect 2681 23563 2747 23566
rect 14089 23563 14155 23566
rect 15377 23626 15443 23629
rect 18278 23626 18338 23702
rect 27337 23699 27403 23702
rect 15377 23624 18338 23626
rect 15377 23568 15382 23624
rect 15438 23568 18338 23624
rect 15377 23566 18338 23568
rect 20621 23626 20687 23629
rect 22185 23626 22251 23629
rect 20621 23624 22251 23626
rect 20621 23568 20626 23624
rect 20682 23568 22190 23624
rect 22246 23568 22251 23624
rect 20621 23566 22251 23568
rect 15377 23563 15443 23566
rect 20621 23563 20687 23566
rect 22185 23563 22251 23566
rect 5349 23490 5415 23493
rect 7097 23490 7163 23493
rect 5349 23488 7163 23490
rect 5349 23432 5354 23488
rect 5410 23432 7102 23488
rect 7158 23432 7163 23488
rect 5349 23430 7163 23432
rect 5349 23427 5415 23430
rect 7097 23427 7163 23430
rect 13721 23490 13787 23493
rect 15285 23490 15351 23493
rect 13721 23488 15351 23490
rect 13721 23432 13726 23488
rect 13782 23432 15290 23488
rect 15346 23432 15351 23488
rect 13721 23430 15351 23432
rect 13721 23427 13787 23430
rect 15285 23427 15351 23430
rect 10277 23424 10597 23425
rect 0 23354 480 23384
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 3417 23354 3483 23357
rect 0 23352 3483 23354
rect 0 23296 3422 23352
rect 3478 23296 3483 23352
rect 0 23294 3483 23296
rect 0 23264 480 23294
rect 3417 23291 3483 23294
rect 23473 23082 23539 23085
rect 27520 23082 28000 23112
rect 23473 23080 28000 23082
rect 23473 23024 23478 23080
rect 23534 23024 28000 23080
rect 23473 23022 28000 23024
rect 23473 23019 23539 23022
rect 27520 22992 28000 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 10961 22538 11027 22541
rect 13721 22538 13787 22541
rect 15377 22538 15443 22541
rect 10961 22536 13554 22538
rect 10961 22480 10966 22536
rect 11022 22480 13554 22536
rect 10961 22478 13554 22480
rect 10961 22475 11027 22478
rect 5073 22402 5139 22405
rect 9121 22402 9187 22405
rect 5073 22400 9187 22402
rect 5073 22344 5078 22400
rect 5134 22344 9126 22400
rect 9182 22344 9187 22400
rect 5073 22342 9187 22344
rect 13494 22402 13554 22478
rect 13721 22536 15443 22538
rect 13721 22480 13726 22536
rect 13782 22480 15382 22536
rect 15438 22480 15443 22536
rect 13721 22478 15443 22480
rect 13721 22475 13787 22478
rect 15377 22475 15443 22478
rect 14549 22402 14615 22405
rect 18413 22402 18479 22405
rect 13494 22400 18479 22402
rect 13494 22344 14554 22400
rect 14610 22344 18418 22400
rect 18474 22344 18479 22400
rect 13494 22342 18479 22344
rect 5073 22339 5139 22342
rect 9121 22339 9187 22342
rect 14549 22339 14615 22342
rect 18413 22339 18479 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 9305 21994 9371 21997
rect 16297 21994 16363 21997
rect 9305 21992 16363 21994
rect 9305 21936 9310 21992
rect 9366 21936 16302 21992
rect 16358 21936 16363 21992
rect 9305 21934 16363 21936
rect 9305 21931 9371 21934
rect 16297 21931 16363 21934
rect 17033 21994 17099 21997
rect 25313 21994 25379 21997
rect 17033 21992 25379 21994
rect 17033 21936 17038 21992
rect 17094 21936 25318 21992
rect 25374 21936 25379 21992
rect 17033 21934 25379 21936
rect 17033 21931 17099 21934
rect 25313 21931 25379 21934
rect 5993 21858 6059 21861
rect 9029 21858 9095 21861
rect 5993 21856 9095 21858
rect 5993 21800 5998 21856
rect 6054 21800 9034 21856
rect 9090 21800 9095 21856
rect 5993 21798 9095 21800
rect 5993 21795 6059 21798
rect 9029 21795 9095 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 24669 21722 24735 21725
rect 27520 21722 28000 21752
rect 24669 21720 28000 21722
rect 24669 21664 24674 21720
rect 24730 21664 28000 21720
rect 24669 21662 28000 21664
rect 24669 21659 24735 21662
rect 27520 21632 28000 21662
rect 16849 21586 16915 21589
rect 9630 21584 16915 21586
rect 9630 21528 16854 21584
rect 16910 21528 16915 21584
rect 9630 21526 16915 21528
rect 8201 21314 8267 21317
rect 9397 21314 9463 21317
rect 9630 21314 9690 21526
rect 16849 21523 16915 21526
rect 11329 21450 11395 21453
rect 15009 21450 15075 21453
rect 15745 21450 15811 21453
rect 11329 21448 15811 21450
rect 11329 21392 11334 21448
rect 11390 21392 15014 21448
rect 15070 21392 15750 21448
rect 15806 21392 15811 21448
rect 11329 21390 15811 21392
rect 11329 21387 11395 21390
rect 15009 21387 15075 21390
rect 15745 21387 15811 21390
rect 8201 21312 9690 21314
rect 8201 21256 8206 21312
rect 8262 21256 9402 21312
rect 9458 21256 9690 21312
rect 8201 21254 9690 21256
rect 8201 21251 8267 21254
rect 9397 21251 9463 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 6177 21042 6243 21045
rect 15285 21042 15351 21045
rect 6177 21040 15351 21042
rect 6177 20984 6182 21040
rect 6238 20984 15290 21040
rect 15346 20984 15351 21040
rect 6177 20982 15351 20984
rect 6177 20979 6243 20982
rect 15285 20979 15351 20982
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 10961 20634 11027 20637
rect 12801 20634 12867 20637
rect 10961 20632 12867 20634
rect 10961 20576 10966 20632
rect 11022 20576 12806 20632
rect 12862 20576 12867 20632
rect 10961 20574 12867 20576
rect 10961 20571 11027 20574
rect 12801 20571 12867 20574
rect 5717 20362 5783 20365
rect 8845 20362 8911 20365
rect 5717 20360 8911 20362
rect 5717 20304 5722 20360
rect 5778 20304 8850 20360
rect 8906 20304 8911 20360
rect 5717 20302 8911 20304
rect 5717 20299 5783 20302
rect 8845 20299 8911 20302
rect 24117 20362 24183 20365
rect 27520 20362 28000 20392
rect 24117 20360 28000 20362
rect 24117 20304 24122 20360
rect 24178 20304 28000 20360
rect 24117 20302 28000 20304
rect 24117 20299 24183 20302
rect 27520 20272 28000 20302
rect 0 20226 480 20256
rect 7281 20226 7347 20229
rect 0 20224 7347 20226
rect 0 20168 7286 20224
rect 7342 20168 7347 20224
rect 0 20166 7347 20168
rect 0 20136 480 20166
rect 7281 20163 7347 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 11973 19954 12039 19957
rect 14641 19954 14707 19957
rect 23841 19954 23907 19957
rect 11973 19952 23907 19954
rect 11973 19896 11978 19952
rect 12034 19896 14646 19952
rect 14702 19896 23846 19952
rect 23902 19896 23907 19952
rect 11973 19894 23907 19896
rect 11973 19891 12039 19894
rect 14641 19891 14707 19894
rect 23841 19891 23907 19894
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 10041 19410 10107 19413
rect 15193 19410 15259 19413
rect 10041 19408 15259 19410
rect 10041 19352 10046 19408
rect 10102 19352 15198 19408
rect 15254 19352 15259 19408
rect 10041 19350 15259 19352
rect 10041 19347 10107 19350
rect 15193 19347 15259 19350
rect 16021 19410 16087 19413
rect 23473 19410 23539 19413
rect 16021 19408 23539 19410
rect 16021 19352 16026 19408
rect 16082 19352 23478 19408
rect 23534 19352 23539 19408
rect 16021 19350 23539 19352
rect 16021 19347 16087 19350
rect 23473 19347 23539 19350
rect 5717 19274 5783 19277
rect 9857 19274 9923 19277
rect 5717 19272 9923 19274
rect 5717 19216 5722 19272
rect 5778 19216 9862 19272
rect 9918 19216 9923 19272
rect 5717 19214 9923 19216
rect 5717 19211 5783 19214
rect 9857 19211 9923 19214
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 5073 18866 5139 18869
rect 15377 18866 15443 18869
rect 23749 18866 23815 18869
rect 5073 18864 23815 18866
rect 5073 18808 5078 18864
rect 5134 18808 15382 18864
rect 15438 18808 23754 18864
rect 23810 18808 23815 18864
rect 5073 18806 23815 18808
rect 5073 18803 5139 18806
rect 15377 18803 15443 18806
rect 23749 18803 23815 18806
rect 24761 18866 24827 18869
rect 27520 18866 28000 18896
rect 24761 18864 28000 18866
rect 24761 18808 24766 18864
rect 24822 18808 28000 18864
rect 24761 18806 28000 18808
rect 24761 18803 24827 18806
rect 27520 18776 28000 18806
rect 11881 18730 11947 18733
rect 15285 18730 15351 18733
rect 24669 18730 24735 18733
rect 11881 18728 24735 18730
rect 11881 18672 11886 18728
rect 11942 18672 15290 18728
rect 15346 18672 24674 18728
rect 24730 18672 24735 18728
rect 11881 18670 24735 18672
rect 11881 18667 11947 18670
rect 15285 18667 15351 18670
rect 24669 18667 24735 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 6453 18186 6519 18189
rect 10041 18186 10107 18189
rect 13169 18186 13235 18189
rect 6453 18184 13235 18186
rect 6453 18128 6458 18184
rect 6514 18128 10046 18184
rect 10102 18128 13174 18184
rect 13230 18128 13235 18184
rect 6453 18126 13235 18128
rect 6453 18123 6519 18126
rect 10041 18123 10107 18126
rect 13169 18123 13235 18126
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 6269 17778 6335 17781
rect 13629 17778 13695 17781
rect 6269 17776 13695 17778
rect 6269 17720 6274 17776
rect 6330 17720 13634 17776
rect 13690 17720 13695 17776
rect 6269 17718 13695 17720
rect 6269 17715 6335 17718
rect 13629 17715 13695 17718
rect 5349 17642 5415 17645
rect 6545 17642 6611 17645
rect 9489 17642 9555 17645
rect 5349 17640 9555 17642
rect 5349 17584 5354 17640
rect 5410 17584 6550 17640
rect 6606 17584 9494 17640
rect 9550 17584 9555 17640
rect 5349 17582 9555 17584
rect 5349 17579 5415 17582
rect 6545 17579 6611 17582
rect 9489 17579 9555 17582
rect 15377 17506 15443 17509
rect 24117 17506 24183 17509
rect 27520 17506 28000 17536
rect 15377 17504 24183 17506
rect 15377 17448 15382 17504
rect 15438 17448 24122 17504
rect 24178 17448 24183 17504
rect 15377 17446 24183 17448
rect 15377 17443 15443 17446
rect 24117 17443 24183 17446
rect 24902 17446 28000 17506
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 8661 17234 8727 17237
rect 15377 17234 15443 17237
rect 8661 17232 15443 17234
rect 8661 17176 8666 17232
rect 8722 17176 15382 17232
rect 15438 17176 15443 17232
rect 8661 17174 15443 17176
rect 8661 17171 8727 17174
rect 15377 17171 15443 17174
rect 0 17098 480 17128
rect 4061 17098 4127 17101
rect 0 17096 4127 17098
rect 0 17040 4066 17096
rect 4122 17040 4127 17096
rect 0 17038 4127 17040
rect 0 17008 480 17038
rect 4061 17035 4127 17038
rect 14089 17098 14155 17101
rect 24761 17098 24827 17101
rect 14089 17096 24827 17098
rect 14089 17040 14094 17096
rect 14150 17040 24766 17096
rect 24822 17040 24827 17096
rect 14089 17038 24827 17040
rect 14089 17035 14155 17038
rect 24761 17035 24827 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 12985 16826 13051 16829
rect 12985 16824 15394 16826
rect 12985 16768 12990 16824
rect 13046 16768 15394 16824
rect 12985 16766 15394 16768
rect 12985 16763 13051 16766
rect 4337 16690 4403 16693
rect 10685 16690 10751 16693
rect 4337 16688 10751 16690
rect 4337 16632 4342 16688
rect 4398 16632 10690 16688
rect 10746 16632 10751 16688
rect 4337 16630 10751 16632
rect 4337 16627 4403 16630
rect 10685 16627 10751 16630
rect 11973 16690 12039 16693
rect 15193 16690 15259 16693
rect 11973 16688 15259 16690
rect 11973 16632 11978 16688
rect 12034 16632 15198 16688
rect 15254 16632 15259 16688
rect 11973 16630 15259 16632
rect 15334 16690 15394 16766
rect 15561 16690 15627 16693
rect 24902 16690 24962 17446
rect 27520 17416 28000 17446
rect 15334 16688 24962 16690
rect 15334 16632 15566 16688
rect 15622 16632 24962 16688
rect 15334 16630 24962 16632
rect 11973 16627 12039 16630
rect 15193 16627 15259 16630
rect 15561 16627 15627 16630
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 6269 16282 6335 16285
rect 10225 16282 10291 16285
rect 6269 16280 10291 16282
rect 6269 16224 6274 16280
rect 6330 16224 10230 16280
rect 10286 16224 10291 16280
rect 6269 16222 10291 16224
rect 6269 16219 6335 16222
rect 10225 16219 10291 16222
rect 27520 16146 28000 16176
rect 27478 16056 28000 16146
rect 5257 16010 5323 16013
rect 14825 16010 14891 16013
rect 5257 16008 14891 16010
rect 5257 15952 5262 16008
rect 5318 15952 14830 16008
rect 14886 15952 14891 16008
rect 5257 15950 14891 15952
rect 5257 15947 5323 15950
rect 14825 15947 14891 15950
rect 6453 15874 6519 15877
rect 8753 15874 8819 15877
rect 6453 15872 8819 15874
rect 6453 15816 6458 15872
rect 6514 15816 8758 15872
rect 8814 15816 8819 15872
rect 6453 15814 8819 15816
rect 6453 15811 6519 15814
rect 8753 15811 8819 15814
rect 17217 15874 17283 15877
rect 19425 15874 19491 15877
rect 17217 15872 19491 15874
rect 17217 15816 17222 15872
rect 17278 15816 19430 15872
rect 19486 15816 19491 15872
rect 17217 15814 19491 15816
rect 17217 15811 17283 15814
rect 19425 15811 19491 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 10501 15466 10567 15469
rect 12617 15466 12683 15469
rect 10501 15464 12683 15466
rect 10501 15408 10506 15464
rect 10562 15408 12622 15464
rect 12678 15408 12683 15464
rect 10501 15406 12683 15408
rect 10501 15403 10567 15406
rect 12617 15403 12683 15406
rect 14825 15466 14891 15469
rect 27478 15466 27538 16056
rect 14825 15464 27538 15466
rect 14825 15408 14830 15464
rect 14886 15408 27538 15464
rect 14825 15406 27538 15408
rect 14825 15403 14891 15406
rect 10685 15330 10751 15333
rect 11237 15330 11303 15333
rect 14457 15330 14523 15333
rect 10685 15328 14523 15330
rect 10685 15272 10690 15328
rect 10746 15272 11242 15328
rect 11298 15272 14462 15328
rect 14518 15272 14523 15328
rect 10685 15270 14523 15272
rect 10685 15267 10751 15270
rect 11237 15267 11303 15270
rect 14457 15267 14523 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 4245 15058 4311 15061
rect 9673 15058 9739 15061
rect 4245 15056 9739 15058
rect 4245 15000 4250 15056
rect 4306 15000 9678 15056
rect 9734 15000 9739 15056
rect 4245 14998 9739 15000
rect 4245 14995 4311 14998
rect 9673 14995 9739 14998
rect 18873 15058 18939 15061
rect 23565 15058 23631 15061
rect 18873 15056 23631 15058
rect 18873 15000 18878 15056
rect 18934 15000 23570 15056
rect 23626 15000 23631 15056
rect 18873 14998 23631 15000
rect 18873 14995 18939 14998
rect 23565 14995 23631 14998
rect 3417 14922 3483 14925
rect 5533 14922 5599 14925
rect 8201 14922 8267 14925
rect 11329 14922 11395 14925
rect 3417 14920 8034 14922
rect 3417 14864 3422 14920
rect 3478 14864 5538 14920
rect 5594 14864 8034 14920
rect 3417 14862 8034 14864
rect 3417 14859 3483 14862
rect 5533 14859 5599 14862
rect 7974 14786 8034 14862
rect 8201 14920 11395 14922
rect 8201 14864 8206 14920
rect 8262 14864 11334 14920
rect 11390 14864 11395 14920
rect 8201 14862 11395 14864
rect 8201 14859 8267 14862
rect 11329 14859 11395 14862
rect 13445 14922 13511 14925
rect 13445 14920 27538 14922
rect 13445 14864 13450 14920
rect 13506 14864 27538 14920
rect 13445 14862 27538 14864
rect 13445 14859 13511 14862
rect 27478 14816 27538 14862
rect 9029 14786 9095 14789
rect 7974 14784 9095 14786
rect 7974 14728 9034 14784
rect 9090 14728 9095 14784
rect 7974 14726 9095 14728
rect 27478 14726 28000 14816
rect 9029 14723 9095 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 27520 14696 28000 14726
rect 19610 14655 19930 14656
rect 10777 14514 10843 14517
rect 13077 14514 13143 14517
rect 10777 14512 13143 14514
rect 10777 14456 10782 14512
rect 10838 14456 13082 14512
rect 13138 14456 13143 14512
rect 10777 14454 13143 14456
rect 10777 14451 10843 14454
rect 13077 14451 13143 14454
rect 19517 14378 19583 14381
rect 21265 14378 21331 14381
rect 19517 14376 21331 14378
rect 19517 14320 19522 14376
rect 19578 14320 21270 14376
rect 21326 14320 21331 14376
rect 19517 14318 21331 14320
rect 19517 14315 19583 14318
rect 21265 14315 21331 14318
rect 9949 14242 10015 14245
rect 10869 14242 10935 14245
rect 14641 14242 14707 14245
rect 9949 14240 14707 14242
rect 9949 14184 9954 14240
rect 10010 14184 10874 14240
rect 10930 14184 14646 14240
rect 14702 14184 14707 14240
rect 9949 14182 14707 14184
rect 9949 14179 10015 14182
rect 10869 14179 10935 14182
rect 14641 14179 14707 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13970 480 14000
rect 4061 13970 4127 13973
rect 0 13968 4127 13970
rect 0 13912 4066 13968
rect 4122 13912 4127 13968
rect 0 13910 4127 13912
rect 0 13880 480 13910
rect 4061 13907 4127 13910
rect 19241 13834 19307 13837
rect 20989 13834 21055 13837
rect 21541 13834 21607 13837
rect 19241 13832 21607 13834
rect 19241 13776 19246 13832
rect 19302 13776 20994 13832
rect 21050 13776 21546 13832
rect 21602 13776 21607 13832
rect 19241 13774 21607 13776
rect 19241 13771 19307 13774
rect 20989 13771 21055 13774
rect 21541 13771 21607 13774
rect 2497 13698 2563 13701
rect 4337 13698 4403 13701
rect 2497 13696 4403 13698
rect 2497 13640 2502 13696
rect 2558 13640 4342 13696
rect 4398 13640 4403 13696
rect 2497 13638 4403 13640
rect 2497 13635 2563 13638
rect 4337 13635 4403 13638
rect 6637 13698 6703 13701
rect 8293 13698 8359 13701
rect 6637 13696 8359 13698
rect 6637 13640 6642 13696
rect 6698 13640 8298 13696
rect 8354 13640 8359 13696
rect 6637 13638 8359 13640
rect 6637 13635 6703 13638
rect 8293 13635 8359 13638
rect 10685 13698 10751 13701
rect 12525 13698 12591 13701
rect 10685 13696 12591 13698
rect 10685 13640 10690 13696
rect 10746 13640 12530 13696
rect 12586 13640 12591 13696
rect 10685 13638 12591 13640
rect 10685 13635 10751 13638
rect 12525 13635 12591 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 24761 13290 24827 13293
rect 27520 13290 28000 13320
rect 24761 13288 28000 13290
rect 24761 13232 24766 13288
rect 24822 13232 28000 13288
rect 24761 13230 28000 13232
rect 24761 13227 24827 13230
rect 27520 13200 28000 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 8477 13018 8543 13021
rect 12433 13018 12499 13021
rect 8477 13016 12499 13018
rect 8477 12960 8482 13016
rect 8538 12960 12438 13016
rect 12494 12960 12499 13016
rect 8477 12958 12499 12960
rect 8477 12955 8543 12958
rect 12433 12955 12499 12958
rect 8109 12882 8175 12885
rect 13445 12882 13511 12885
rect 8109 12880 13511 12882
rect 8109 12824 8114 12880
rect 8170 12824 13450 12880
rect 13506 12824 13511 12880
rect 8109 12822 13511 12824
rect 8109 12819 8175 12822
rect 13445 12819 13511 12822
rect 20621 12882 20687 12885
rect 20897 12882 20963 12885
rect 22461 12882 22527 12885
rect 20621 12880 22527 12882
rect 20621 12824 20626 12880
rect 20682 12824 20902 12880
rect 20958 12824 22466 12880
rect 22522 12824 22527 12880
rect 20621 12822 22527 12824
rect 20621 12819 20687 12822
rect 20897 12819 20963 12822
rect 22461 12819 22527 12822
rect 2865 12746 2931 12749
rect 7557 12746 7623 12749
rect 2865 12744 7623 12746
rect 2865 12688 2870 12744
rect 2926 12688 7562 12744
rect 7618 12688 7623 12744
rect 2865 12686 7623 12688
rect 2865 12683 2931 12686
rect 7557 12683 7623 12686
rect 7833 12746 7899 12749
rect 9489 12746 9555 12749
rect 14181 12746 14247 12749
rect 7833 12744 14247 12746
rect 7833 12688 7838 12744
rect 7894 12688 9494 12744
rect 9550 12688 14186 12744
rect 14242 12688 14247 12744
rect 7833 12686 14247 12688
rect 7833 12683 7899 12686
rect 9489 12683 9555 12686
rect 14181 12683 14247 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 3601 12338 3667 12341
rect 7189 12338 7255 12341
rect 3601 12336 7255 12338
rect 3601 12280 3606 12336
rect 3662 12280 7194 12336
rect 7250 12280 7255 12336
rect 3601 12278 7255 12280
rect 3601 12275 3667 12278
rect 7189 12275 7255 12278
rect 9581 12338 9647 12341
rect 11513 12338 11579 12341
rect 9581 12336 11579 12338
rect 9581 12280 9586 12336
rect 9642 12280 11518 12336
rect 11574 12280 11579 12336
rect 9581 12278 11579 12280
rect 9581 12275 9647 12278
rect 11513 12275 11579 12278
rect 15837 12338 15903 12341
rect 18781 12338 18847 12341
rect 15837 12336 18847 12338
rect 15837 12280 15842 12336
rect 15898 12280 18786 12336
rect 18842 12280 18847 12336
rect 15837 12278 18847 12280
rect 15837 12275 15903 12278
rect 18781 12275 18847 12278
rect 2589 12202 2655 12205
rect 8753 12202 8819 12205
rect 2589 12200 8819 12202
rect 2589 12144 2594 12200
rect 2650 12144 8758 12200
rect 8814 12144 8819 12200
rect 2589 12142 8819 12144
rect 2589 12139 2655 12142
rect 8753 12139 8819 12142
rect 9121 12202 9187 12205
rect 15285 12202 15351 12205
rect 9121 12200 15351 12202
rect 9121 12144 9126 12200
rect 9182 12144 15290 12200
rect 15346 12144 15351 12200
rect 9121 12142 15351 12144
rect 9121 12139 9187 12142
rect 15285 12139 15351 12142
rect 6545 12066 6611 12069
rect 8569 12066 8635 12069
rect 13813 12066 13879 12069
rect 6545 12064 13879 12066
rect 6545 12008 6550 12064
rect 6606 12008 8574 12064
rect 8630 12008 13818 12064
rect 13874 12008 13879 12064
rect 6545 12006 13879 12008
rect 6545 12003 6611 12006
rect 8569 12003 8635 12006
rect 13813 12003 13879 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 24761 11930 24827 11933
rect 27520 11930 28000 11960
rect 24761 11928 28000 11930
rect 24761 11872 24766 11928
rect 24822 11872 28000 11928
rect 24761 11870 28000 11872
rect 24761 11867 24827 11870
rect 27520 11840 28000 11870
rect 2221 11658 2287 11661
rect 15653 11658 15719 11661
rect 2221 11656 15719 11658
rect 2221 11600 2226 11656
rect 2282 11600 15658 11656
rect 15714 11600 15719 11656
rect 2221 11598 15719 11600
rect 2221 11595 2287 11598
rect 15653 11595 15719 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 7925 11386 7991 11389
rect 8477 11386 8543 11389
rect 9765 11386 9831 11389
rect 7925 11384 9831 11386
rect 7925 11328 7930 11384
rect 7986 11328 8482 11384
rect 8538 11328 9770 11384
rect 9826 11328 9831 11384
rect 7925 11326 9831 11328
rect 7925 11323 7991 11326
rect 8477 11323 8543 11326
rect 9765 11323 9831 11326
rect 8845 11250 8911 11253
rect 9581 11250 9647 11253
rect 22461 11250 22527 11253
rect 8845 11248 9647 11250
rect 8845 11192 8850 11248
rect 8906 11192 9586 11248
rect 9642 11192 9647 11248
rect 8845 11190 9647 11192
rect 8845 11187 8911 11190
rect 9581 11187 9647 11190
rect 14184 11248 22527 11250
rect 14184 11192 22466 11248
rect 22522 11192 22527 11248
rect 14184 11190 22527 11192
rect 14184 11117 14244 11190
rect 22461 11187 22527 11190
rect 12985 11114 13051 11117
rect 14181 11114 14247 11117
rect 12985 11112 14247 11114
rect 12985 11056 12990 11112
rect 13046 11056 14186 11112
rect 14242 11056 14247 11112
rect 12985 11054 14247 11056
rect 12985 11051 13051 11054
rect 14181 11051 14247 11054
rect 20437 11114 20503 11117
rect 22185 11114 22251 11117
rect 20437 11112 22251 11114
rect 20437 11056 20442 11112
rect 20498 11056 22190 11112
rect 22246 11056 22251 11112
rect 20437 11054 22251 11056
rect 20437 11051 20503 11054
rect 22185 11051 22251 11054
rect 5610 10912 5930 10913
rect 0 10842 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 3325 10842 3391 10845
rect 0 10840 3391 10842
rect 0 10784 3330 10840
rect 3386 10784 3391 10840
rect 0 10782 3391 10784
rect 0 10752 480 10782
rect 3325 10779 3391 10782
rect 9857 10842 9923 10845
rect 12893 10842 12959 10845
rect 9857 10840 12959 10842
rect 9857 10784 9862 10840
rect 9918 10784 12898 10840
rect 12954 10784 12959 10840
rect 9857 10782 12959 10784
rect 9857 10779 9923 10782
rect 12893 10779 12959 10782
rect 3693 10706 3759 10709
rect 5993 10706 6059 10709
rect 6637 10706 6703 10709
rect 3693 10704 6703 10706
rect 3693 10648 3698 10704
rect 3754 10648 5998 10704
rect 6054 10648 6642 10704
rect 6698 10648 6703 10704
rect 3693 10646 6703 10648
rect 3693 10643 3759 10646
rect 5993 10643 6059 10646
rect 6637 10643 6703 10646
rect 11053 10706 11119 10709
rect 15285 10706 15351 10709
rect 11053 10704 15351 10706
rect 11053 10648 11058 10704
rect 11114 10648 15290 10704
rect 15346 10648 15351 10704
rect 11053 10646 15351 10648
rect 11053 10643 11119 10646
rect 15285 10643 15351 10646
rect 11881 10570 11947 10573
rect 14641 10570 14707 10573
rect 24301 10570 24367 10573
rect 11881 10568 24367 10570
rect 11881 10512 11886 10568
rect 11942 10512 14646 10568
rect 14702 10512 24306 10568
rect 24362 10512 24367 10568
rect 11881 10510 24367 10512
rect 11881 10507 11947 10510
rect 14641 10507 14707 10510
rect 24301 10507 24367 10510
rect 24761 10570 24827 10573
rect 27520 10570 28000 10600
rect 24761 10568 28000 10570
rect 24761 10512 24766 10568
rect 24822 10512 28000 10568
rect 24761 10510 28000 10512
rect 24761 10507 24827 10510
rect 27520 10480 28000 10510
rect 4061 10434 4127 10437
rect 5533 10434 5599 10437
rect 4061 10432 5599 10434
rect 4061 10376 4066 10432
rect 4122 10376 5538 10432
rect 5594 10376 5599 10432
rect 4061 10374 5599 10376
rect 4061 10371 4127 10374
rect 5533 10371 5599 10374
rect 6637 10434 6703 10437
rect 9673 10434 9739 10437
rect 6637 10432 9739 10434
rect 6637 10376 6642 10432
rect 6698 10376 9678 10432
rect 9734 10376 9739 10432
rect 6637 10374 9739 10376
rect 6637 10371 6703 10374
rect 9673 10371 9739 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 3141 10162 3207 10165
rect 9673 10162 9739 10165
rect 3141 10160 9739 10162
rect 3141 10104 3146 10160
rect 3202 10104 9678 10160
rect 9734 10104 9739 10160
rect 3141 10102 9739 10104
rect 3141 10099 3207 10102
rect 9673 10099 9739 10102
rect 7557 9890 7623 9893
rect 12157 9890 12223 9893
rect 7557 9888 12223 9890
rect 7557 9832 7562 9888
rect 7618 9832 12162 9888
rect 12218 9832 12223 9888
rect 7557 9830 12223 9832
rect 7557 9827 7623 9830
rect 12157 9827 12223 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 9489 9754 9555 9757
rect 12433 9754 12499 9757
rect 9489 9752 12499 9754
rect 9489 9696 9494 9752
rect 9550 9696 12438 9752
rect 12494 9696 12499 9752
rect 9489 9694 12499 9696
rect 9489 9691 9555 9694
rect 12433 9691 12499 9694
rect 6821 9618 6887 9621
rect 9305 9618 9371 9621
rect 6821 9616 9371 9618
rect 6821 9560 6826 9616
rect 6882 9560 9310 9616
rect 9366 9560 9371 9616
rect 6821 9558 9371 9560
rect 6821 9555 6887 9558
rect 9305 9555 9371 9558
rect 12525 9618 12591 9621
rect 15929 9618 15995 9621
rect 12525 9616 15995 9618
rect 12525 9560 12530 9616
rect 12586 9560 15934 9616
rect 15990 9560 15995 9616
rect 12525 9558 15995 9560
rect 12525 9555 12591 9558
rect 15929 9555 15995 9558
rect 5441 9346 5507 9349
rect 7005 9346 7071 9349
rect 5441 9344 7071 9346
rect 5441 9288 5446 9344
rect 5502 9288 7010 9344
rect 7066 9288 7071 9344
rect 5441 9286 7071 9288
rect 5441 9283 5507 9286
rect 7005 9283 7071 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 12341 9074 12407 9077
rect 12893 9074 12959 9077
rect 16113 9074 16179 9077
rect 12341 9072 16179 9074
rect 12341 9016 12346 9072
rect 12402 9016 12898 9072
rect 12954 9016 16118 9072
rect 16174 9016 16179 9072
rect 12341 9014 16179 9016
rect 12341 9011 12407 9014
rect 12893 9011 12959 9014
rect 16113 9011 16179 9014
rect 16665 9074 16731 9077
rect 23565 9074 23631 9077
rect 16665 9072 23631 9074
rect 16665 9016 16670 9072
rect 16726 9016 23570 9072
rect 23626 9016 23631 9072
rect 16665 9014 23631 9016
rect 16665 9011 16731 9014
rect 23565 9011 23631 9014
rect 24761 9074 24827 9077
rect 27520 9074 28000 9104
rect 24761 9072 28000 9074
rect 24761 9016 24766 9072
rect 24822 9016 28000 9072
rect 24761 9014 28000 9016
rect 24761 9011 24827 9014
rect 27520 8984 28000 9014
rect 18781 8938 18847 8941
rect 20989 8938 21055 8941
rect 18781 8936 21055 8938
rect 18781 8880 18786 8936
rect 18842 8880 20994 8936
rect 21050 8880 21055 8936
rect 18781 8878 21055 8880
rect 18781 8875 18847 8878
rect 20989 8875 21055 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 5993 8666 6059 8669
rect 8661 8666 8727 8669
rect 5993 8664 8727 8666
rect 5993 8608 5998 8664
rect 6054 8608 8666 8664
rect 8722 8608 8727 8664
rect 5993 8606 8727 8608
rect 5993 8603 6059 8606
rect 8661 8603 8727 8606
rect 12617 8394 12683 8397
rect 14089 8394 14155 8397
rect 12617 8392 14155 8394
rect 12617 8336 12622 8392
rect 12678 8336 14094 8392
rect 14150 8336 14155 8392
rect 12617 8334 14155 8336
rect 12617 8331 12683 8334
rect 14089 8331 14155 8334
rect 6453 8258 6519 8261
rect 9857 8258 9923 8261
rect 6453 8256 9923 8258
rect 6453 8200 6458 8256
rect 6514 8200 9862 8256
rect 9918 8200 9923 8256
rect 6453 8198 9923 8200
rect 6453 8195 6519 8198
rect 9857 8195 9923 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 5165 7986 5231 7989
rect 6269 7986 6335 7989
rect 9765 7986 9831 7989
rect 5165 7984 9831 7986
rect 5165 7928 5170 7984
rect 5226 7928 6274 7984
rect 6330 7928 9770 7984
rect 9826 7928 9831 7984
rect 5165 7926 9831 7928
rect 5165 7923 5231 7926
rect 6269 7923 6335 7926
rect 9765 7923 9831 7926
rect 8753 7850 8819 7853
rect 12433 7850 12499 7853
rect 8753 7848 12499 7850
rect 8753 7792 8758 7848
rect 8814 7792 12438 7848
rect 12494 7792 12499 7848
rect 8753 7790 12499 7792
rect 8753 7787 8819 7790
rect 12433 7787 12499 7790
rect 20529 7850 20595 7853
rect 24577 7850 24643 7853
rect 20529 7848 24643 7850
rect 20529 7792 20534 7848
rect 20590 7792 24582 7848
rect 24638 7792 24643 7848
rect 20529 7790 24643 7792
rect 20529 7787 20595 7790
rect 24577 7787 24643 7790
rect 0 7714 480 7744
rect 2589 7714 2655 7717
rect 0 7712 2655 7714
rect 0 7656 2594 7712
rect 2650 7656 2655 7712
rect 0 7654 2655 7656
rect 0 7624 480 7654
rect 2589 7651 2655 7654
rect 19885 7714 19951 7717
rect 23473 7714 23539 7717
rect 19885 7712 23539 7714
rect 19885 7656 19890 7712
rect 19946 7656 23478 7712
rect 23534 7656 23539 7712
rect 19885 7654 23539 7656
rect 19885 7651 19951 7654
rect 23473 7651 23539 7654
rect 24669 7714 24735 7717
rect 27520 7714 28000 7744
rect 24669 7712 28000 7714
rect 24669 7656 24674 7712
rect 24730 7656 28000 7712
rect 24669 7654 28000 7656
rect 24669 7651 24735 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7654
rect 24277 7583 24597 7584
rect 9581 7578 9647 7581
rect 12525 7578 12591 7581
rect 9581 7576 12591 7578
rect 9581 7520 9586 7576
rect 9642 7520 12530 7576
rect 12586 7520 12591 7576
rect 9581 7518 12591 7520
rect 9581 7515 9647 7518
rect 12525 7515 12591 7518
rect 5441 7442 5507 7445
rect 6361 7442 6427 7445
rect 10501 7442 10567 7445
rect 5441 7440 10567 7442
rect 5441 7384 5446 7440
rect 5502 7384 6366 7440
rect 6422 7384 10506 7440
rect 10562 7384 10567 7440
rect 5441 7382 10567 7384
rect 5441 7379 5507 7382
rect 6361 7379 6427 7382
rect 10501 7379 10567 7382
rect 14917 7442 14983 7445
rect 22829 7442 22895 7445
rect 14917 7440 22895 7442
rect 14917 7384 14922 7440
rect 14978 7384 22834 7440
rect 22890 7384 22895 7440
rect 14917 7382 22895 7384
rect 14917 7379 14983 7382
rect 22829 7379 22895 7382
rect 18965 7306 19031 7309
rect 20989 7306 21055 7309
rect 18965 7304 21055 7306
rect 18965 7248 18970 7304
rect 19026 7248 20994 7304
rect 21050 7248 21055 7304
rect 18965 7246 21055 7248
rect 18965 7243 19031 7246
rect 20989 7243 21055 7246
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 3877 6898 3943 6901
rect 6913 6898 6979 6901
rect 3877 6896 6979 6898
rect 3877 6840 3882 6896
rect 3938 6840 6918 6896
rect 6974 6840 6979 6896
rect 3877 6838 6979 6840
rect 3877 6835 3943 6838
rect 6913 6835 6979 6838
rect 7189 6898 7255 6901
rect 11145 6898 11211 6901
rect 7189 6896 11211 6898
rect 7189 6840 7194 6896
rect 7250 6840 11150 6896
rect 11206 6840 11211 6896
rect 7189 6838 11211 6840
rect 7189 6835 7255 6838
rect 11145 6835 11211 6838
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 5441 6354 5507 6357
rect 7925 6354 7991 6357
rect 5441 6352 7991 6354
rect 5441 6296 5446 6352
rect 5502 6296 7930 6352
rect 7986 6296 7991 6352
rect 5441 6294 7991 6296
rect 5441 6291 5507 6294
rect 7925 6291 7991 6294
rect 22645 6354 22711 6357
rect 24577 6354 24643 6357
rect 22645 6352 24643 6354
rect 22645 6296 22650 6352
rect 22706 6296 24582 6352
rect 24638 6296 24643 6352
rect 22645 6294 24643 6296
rect 22645 6291 22711 6294
rect 24577 6291 24643 6294
rect 24761 6354 24827 6357
rect 27520 6354 28000 6384
rect 24761 6352 28000 6354
rect 24761 6296 24766 6352
rect 24822 6296 28000 6352
rect 24761 6294 28000 6296
rect 24761 6291 24827 6294
rect 27520 6264 28000 6294
rect 8661 6218 8727 6221
rect 13445 6218 13511 6221
rect 8661 6216 13511 6218
rect 8661 6160 8666 6216
rect 8722 6160 13450 6216
rect 13506 6160 13511 6216
rect 8661 6158 13511 6160
rect 8661 6155 8727 6158
rect 13445 6155 13511 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 7833 5946 7899 5949
rect 9857 5946 9923 5949
rect 7833 5944 9923 5946
rect 7833 5888 7838 5944
rect 7894 5888 9862 5944
rect 9918 5888 9923 5944
rect 7833 5886 9923 5888
rect 7833 5883 7899 5886
rect 9857 5883 9923 5886
rect 10041 5810 10107 5813
rect 14641 5810 14707 5813
rect 17585 5810 17651 5813
rect 10041 5808 17651 5810
rect 10041 5752 10046 5808
rect 10102 5752 14646 5808
rect 14702 5752 17590 5808
rect 17646 5752 17651 5808
rect 10041 5750 17651 5752
rect 10041 5747 10107 5750
rect 14641 5747 14707 5750
rect 17585 5747 17651 5750
rect 13629 5674 13695 5677
rect 23473 5674 23539 5677
rect 13629 5672 23539 5674
rect 13629 5616 13634 5672
rect 13690 5616 23478 5672
rect 23534 5616 23539 5672
rect 13629 5614 23539 5616
rect 13629 5611 13695 5614
rect 23473 5611 23539 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 8109 5130 8175 5133
rect 9765 5130 9831 5133
rect 8109 5128 9831 5130
rect 8109 5072 8114 5128
rect 8170 5072 9770 5128
rect 9826 5072 9831 5128
rect 8109 5070 9831 5072
rect 8109 5067 8175 5070
rect 9765 5067 9831 5070
rect 25129 4994 25195 4997
rect 27337 4994 27403 4997
rect 25129 4992 27403 4994
rect 25129 4936 25134 4992
rect 25190 4936 27342 4992
rect 27398 4936 27403 4992
rect 25129 4934 27403 4936
rect 25129 4931 25195 4934
rect 27337 4931 27403 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 24761 4858 24827 4861
rect 27520 4858 28000 4888
rect 24761 4856 28000 4858
rect 24761 4800 24766 4856
rect 24822 4800 28000 4856
rect 24761 4798 28000 4800
rect 24761 4795 24827 4798
rect 27520 4768 28000 4798
rect 0 4586 480 4616
rect 4061 4586 4127 4589
rect 0 4584 4127 4586
rect 0 4528 4066 4584
rect 4122 4528 4127 4584
rect 0 4526 4127 4528
rect 0 4496 480 4526
rect 4061 4523 4127 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 9029 4178 9095 4181
rect 11789 4178 11855 4181
rect 18965 4178 19031 4181
rect 19977 4178 20043 4181
rect 9029 4176 20043 4178
rect 9029 4120 9034 4176
rect 9090 4120 11794 4176
rect 11850 4120 18970 4176
rect 19026 4120 19982 4176
rect 20038 4120 20043 4176
rect 9029 4118 20043 4120
rect 9029 4115 9095 4118
rect 11789 4115 11855 4118
rect 18965 4115 19031 4118
rect 19977 4115 20043 4118
rect 10685 4042 10751 4045
rect 15929 4042 15995 4045
rect 18045 4042 18111 4045
rect 10685 4040 14842 4042
rect 10685 3984 10690 4040
rect 10746 3984 14842 4040
rect 10685 3982 14842 3984
rect 10685 3979 10751 3982
rect 5441 3906 5507 3909
rect 10041 3906 10107 3909
rect 5441 3904 10107 3906
rect 5441 3848 5446 3904
rect 5502 3848 10046 3904
rect 10102 3848 10107 3904
rect 5441 3846 10107 3848
rect 5441 3843 5507 3846
rect 10041 3843 10107 3846
rect 10685 3906 10751 3909
rect 10685 3904 14658 3906
rect 10685 3848 10690 3904
rect 10746 3848 14658 3904
rect 10685 3846 14658 3848
rect 10685 3843 10751 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 2681 3634 2747 3637
rect 10133 3634 10199 3637
rect 2681 3632 10199 3634
rect 2681 3576 2686 3632
rect 2742 3576 10138 3632
rect 10194 3576 10199 3632
rect 2681 3574 10199 3576
rect 2681 3571 2747 3574
rect 10133 3571 10199 3574
rect 14598 3498 14658 3846
rect 14782 3770 14842 3982
rect 15929 4040 18111 4042
rect 15929 3984 15934 4040
rect 15990 3984 18050 4040
rect 18106 3984 18111 4040
rect 15929 3982 18111 3984
rect 15929 3979 15995 3982
rect 18045 3979 18111 3982
rect 14917 3906 14983 3909
rect 15929 3906 15995 3909
rect 14917 3904 15995 3906
rect 14917 3848 14922 3904
rect 14978 3848 15934 3904
rect 15990 3848 15995 3904
rect 14917 3846 15995 3848
rect 14917 3843 14983 3846
rect 15929 3843 15995 3846
rect 16113 3906 16179 3909
rect 16113 3904 19442 3906
rect 16113 3848 16118 3904
rect 16174 3848 19442 3904
rect 16113 3846 19442 3848
rect 16113 3843 16179 3846
rect 17953 3770 18019 3773
rect 14782 3768 18019 3770
rect 14782 3712 17958 3768
rect 18014 3712 18019 3768
rect 14782 3710 18019 3712
rect 17953 3707 18019 3710
rect 14825 3634 14891 3637
rect 17217 3634 17283 3637
rect 14825 3632 17283 3634
rect 14825 3576 14830 3632
rect 14886 3576 17222 3632
rect 17278 3576 17283 3632
rect 14825 3574 17283 3576
rect 19382 3634 19442 3846
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 21725 3634 21791 3637
rect 19382 3632 21791 3634
rect 19382 3576 21730 3632
rect 21786 3576 21791 3632
rect 19382 3574 21791 3576
rect 14825 3571 14891 3574
rect 17217 3571 17283 3574
rect 21725 3571 21791 3574
rect 17125 3498 17191 3501
rect 14598 3496 17191 3498
rect 14598 3440 17130 3496
rect 17186 3440 17191 3496
rect 14598 3438 17191 3440
rect 17125 3435 17191 3438
rect 17585 3498 17651 3501
rect 21633 3498 21699 3501
rect 17585 3496 21699 3498
rect 17585 3440 17590 3496
rect 17646 3440 21638 3496
rect 21694 3440 21699 3496
rect 17585 3438 21699 3440
rect 17585 3435 17651 3438
rect 21633 3435 21699 3438
rect 21817 3498 21883 3501
rect 27520 3498 28000 3528
rect 21817 3496 28000 3498
rect 21817 3440 21822 3496
rect 21878 3440 28000 3496
rect 21817 3438 28000 3440
rect 21817 3435 21883 3438
rect 27520 3408 28000 3438
rect 15377 3362 15443 3365
rect 21081 3362 21147 3365
rect 15377 3360 21147 3362
rect 15377 3304 15382 3360
rect 15438 3304 21086 3360
rect 21142 3304 21147 3360
rect 15377 3302 21147 3304
rect 15377 3299 15443 3302
rect 21081 3299 21147 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 7741 3226 7807 3229
rect 8477 3226 8543 3229
rect 9857 3226 9923 3229
rect 7741 3224 9923 3226
rect 7741 3168 7746 3224
rect 7802 3168 8482 3224
rect 8538 3168 9862 3224
rect 9918 3168 9923 3224
rect 7741 3166 9923 3168
rect 7741 3163 7807 3166
rect 8477 3163 8543 3166
rect 9857 3163 9923 3166
rect 13905 3226 13971 3229
rect 20345 3226 20411 3229
rect 13905 3224 14842 3226
rect 13905 3168 13910 3224
rect 13966 3168 14842 3224
rect 13905 3166 14842 3168
rect 13905 3163 13971 3166
rect 9765 3090 9831 3093
rect 14549 3090 14615 3093
rect 9765 3088 14615 3090
rect 9765 3032 9770 3088
rect 9826 3032 14554 3088
rect 14610 3032 14615 3088
rect 9765 3030 14615 3032
rect 14782 3090 14842 3166
rect 15334 3224 20411 3226
rect 15334 3168 20350 3224
rect 20406 3168 20411 3224
rect 15334 3166 20411 3168
rect 15334 3090 15394 3166
rect 20345 3163 20411 3166
rect 14782 3030 15394 3090
rect 20437 3090 20503 3093
rect 22185 3090 22251 3093
rect 20437 3088 22251 3090
rect 20437 3032 20442 3088
rect 20498 3032 22190 3088
rect 22246 3032 22251 3088
rect 20437 3030 22251 3032
rect 9765 3027 9831 3030
rect 14549 3027 14615 3030
rect 20437 3027 20503 3030
rect 22185 3027 22251 3030
rect 13721 2954 13787 2957
rect 24301 2954 24367 2957
rect 13721 2952 24367 2954
rect 13721 2896 13726 2952
rect 13782 2896 24306 2952
rect 24362 2896 24367 2952
rect 13721 2894 24367 2896
rect 13721 2891 13787 2894
rect 24301 2891 24367 2894
rect 3509 2818 3575 2821
rect 6361 2818 6427 2821
rect 3509 2816 6427 2818
rect 3509 2760 3514 2816
rect 3570 2760 6366 2816
rect 6422 2760 6427 2816
rect 3509 2758 6427 2760
rect 3509 2755 3575 2758
rect 6361 2755 6427 2758
rect 10961 2818 11027 2821
rect 19425 2818 19491 2821
rect 10961 2816 19491 2818
rect 10961 2760 10966 2816
rect 11022 2760 19430 2816
rect 19486 2760 19491 2816
rect 10961 2758 19491 2760
rect 10961 2755 11027 2758
rect 19425 2755 19491 2758
rect 21909 2818 21975 2821
rect 24209 2818 24275 2821
rect 21909 2816 24275 2818
rect 21909 2760 21914 2816
rect 21970 2760 24214 2816
rect 24270 2760 24275 2816
rect 21909 2758 24275 2760
rect 21909 2755 21975 2758
rect 24209 2755 24275 2758
rect 24485 2818 24551 2821
rect 26325 2818 26391 2821
rect 24485 2816 26391 2818
rect 24485 2760 24490 2816
rect 24546 2760 26330 2816
rect 26386 2760 26391 2816
rect 24485 2758 26391 2760
rect 24485 2755 24551 2758
rect 26325 2755 26391 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 1577 2682 1643 2685
rect 7189 2682 7255 2685
rect 1577 2680 7255 2682
rect 1577 2624 1582 2680
rect 1638 2624 7194 2680
rect 7250 2624 7255 2680
rect 1577 2622 7255 2624
rect 1577 2619 1643 2622
rect 7189 2619 7255 2622
rect 1485 2546 1551 2549
rect 4613 2546 4679 2549
rect 8017 2546 8083 2549
rect 1485 2544 4538 2546
rect 1485 2488 1490 2544
rect 1546 2488 4538 2544
rect 1485 2486 4538 2488
rect 1485 2483 1551 2486
rect 4478 2410 4538 2486
rect 4613 2544 8083 2546
rect 4613 2488 4618 2544
rect 4674 2488 8022 2544
rect 8078 2488 8083 2544
rect 4613 2486 8083 2488
rect 4613 2483 4679 2486
rect 8017 2483 8083 2486
rect 9857 2410 9923 2413
rect 4478 2408 9923 2410
rect 4478 2352 9862 2408
rect 9918 2352 9923 2408
rect 4478 2350 9923 2352
rect 9857 2347 9923 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 24761 2138 24827 2141
rect 27520 2138 28000 2168
rect 24761 2136 28000 2138
rect 24761 2080 24766 2136
rect 24822 2080 28000 2136
rect 24761 2078 28000 2080
rect 24761 2075 24827 2078
rect 27520 2048 28000 2078
rect 473 1866 539 1869
rect 1393 1866 1459 1869
rect 473 1864 1459 1866
rect 473 1808 478 1864
rect 534 1808 1398 1864
rect 1454 1808 1459 1864
rect 473 1806 1459 1808
rect 473 1803 539 1806
rect 1393 1803 1459 1806
rect 0 1594 480 1624
rect 2865 1594 2931 1597
rect 0 1592 2931 1594
rect 0 1536 2870 1592
rect 2926 1536 2931 1592
rect 0 1534 2931 1536
rect 0 1504 480 1534
rect 2865 1531 2931 1534
rect 24669 778 24735 781
rect 27520 778 28000 808
rect 24669 776 28000 778
rect 24669 720 24674 776
rect 24730 720 28000 776
rect 24669 718 28000 720
rect 24669 715 24735 718
rect 27520 688 28000 718
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_8  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_11 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_14 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_22
timestamp 1586364061
transform 1 0 3128 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_0_30
timestamp 1586364061
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_39
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_43
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 774 592
use scs8hd_decap_8  FILLER_1_48
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_56
timestamp 1586364061
transform 1 0 6256 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_61
timestamp 1586364061
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_55 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6164 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_69
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_65
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_83
timestamp 1586364061
transform 1 0 8740 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_73
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_77
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_89
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_96
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_91
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_104
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_100
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_109
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_121
timestamp 1586364061
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_121
timestamp 1586364061
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_154
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_171
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_166
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_182
timestamp 1586364061
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_183
timestamp 1586364061
transform 1 0 17940 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _216_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _215_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_188
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_195
timestamp 1586364061
transform 1 0 19044 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_191
timestamp 1586364061
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__215__A
timestamp 1586364061
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__A
timestamp 1586364061
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_192
timestamp 1586364061
transform 1 0 18768 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _214_
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__214__A
timestamp 1586364061
transform 1 0 19964 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_203
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_207
timestamp 1586364061
transform 1 0 20148 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_204
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_222
timestamp 1586364061
transform 1 0 21528 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_216
timestamp 1586364061
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_215
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _212_
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_226
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_228
timestamp 1586364061
transform 1 0 22080 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__212__A
timestamp 1586364061
transform 1 0 21712 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _211_
timestamp 1586364061
transform 1 0 21712 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_230
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_232
timestamp 1586364061
transform 1 0 22448 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_242
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 24288 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_251
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_256
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_260
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_272
timestamp 1586364061
transform 1 0 26128 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_276
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_11
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_49
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_77
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_86
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_107
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11684 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_111
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_2_118
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 21620 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_76
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_80
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_93
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 590 592
use scs8hd_decap_4  FILLER_3_140
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__217__A
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_151
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_3_161
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_182
timestamp 1586364061
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _213_
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__213__A
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_212
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_216
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_228
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_253
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_conb_1  _189_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_77
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_4  FILLER_4_87
timestamp 1586364061
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_96
timestamp 1586364061
transform 1 0 9936 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_100
timestamp 1586364061
transform 1 0 10304 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_113
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_130
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_134
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _217_
timestamp 1586364061
transform 1 0 15732 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_175
timestamp 1586364061
transform 1 0 17204 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_179
timestamp 1586364061
transform 1 0 17572 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_183
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_195
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_207
timestamp 1586364061
transform 1 0 20148 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_259
timestamp 1586364061
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_271
timestamp 1586364061
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_77
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_83
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_102
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_149
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_164
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_187
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_198
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_202
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_226
timestamp 1586364061
transform 1 0 21896 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_5_238
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 590 592
use scs8hd_decap_8  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_253
timestamp 1586364061
transform 1 0 24380 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_262
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_274
timestamp 1586364061
transform 1 0 26312 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_35
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 314 592
use scs8hd_nor2_4  _140_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_46
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_58
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_76
timestamp 1586364061
transform 1 0 8096 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_72
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_83
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_107
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_115
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_6_133
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_137
timestamp 1586364061
transform 1 0 13708 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _182_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_160
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 406 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_6  FILLER_6_173
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_192
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_188
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_210
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_214
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_229
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_241
timestamp 1586364061
transform 1 0 23276 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 774 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 24564 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_253
timestamp 1586364061
transform 1 0 24380 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_259
timestamp 1586364061
transform 1 0 24932 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_263
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_29
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_40
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_43
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_55
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_60
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_74
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_78
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_82
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_86
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_4  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_182
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_199
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_203
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_236
timestamp 1586364061
transform 1 0 22816 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_248
timestamp 1586364061
transform 1 0 23920 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_260
timestamp 1586364061
transform 1 0 25024 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_272
timestamp 1586364061
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_36
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_40
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7360 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_96
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_138
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_142
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_151
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_164
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_168
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_181
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_188
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_201
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_205
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_212
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_216
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_253
timestamp 1586364061
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_262
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_266
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_274
timestamp 1586364061
transform 1 0 26312 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_40
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_54
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_89
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 9752 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_103
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_135
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_194
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_201
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_205
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_218
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_222
timestamp 1586364061
transform 1 0 21528 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_226
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_238
timestamp 1586364061
transform 1 0 23000 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 24564 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_4  FILLER_10_250
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_254
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_259
timestamp 1586364061
transform 1 0 24932 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_271
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_31
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_or3_4  _099_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_38
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_78
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_97
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _128_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_116
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_126
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_130
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_149
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_153
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 774 592
use scs8hd_conb_1  _193_
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_195
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_199
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_212
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 314 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_229
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_241
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_249
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 406 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 24380 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_261
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_273
timestamp 1586364061
transform 1 0 26220 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_50
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 6072 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_81
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_12_86
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_112
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_116
timestamp 1586364061
transform 1 0 11776 0 -1 9248
box -38 -48 314 592
use scs8hd_buf_1  _156_
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_130
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_134
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 590 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_169
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_201
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_228
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_240
timestamp 1586364061
transform 1 0 23184 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_247
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_259
timestamp 1586364061
transform 1 0 24932 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_271
timestamp 1586364061
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_6  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_11
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_9
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__C
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_or3_4  _077_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_8  _075_
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_20
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_35
timestamp 1586364061
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_38
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__C
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__C
timestamp 1586364061
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_51
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_52
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_or3_4  _093_
timestamp 1586364061
transform 1 0 4968 0 -1 10336
box -38 -48 866 592
use scs8hd_or3_4  _090_
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_62
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_56
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_70
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_66
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__C
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7544 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_85
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_81
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_96
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_96
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 10120 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _078_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_100
timestamp 1586364061
transform 1 0 10304 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_100
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_122
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__D
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_137
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_149
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_conb_1  _192_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_157
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_157
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _159_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1602 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__C
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__D
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_161
timestamp 1586364061
transform 1 0 15916 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_195
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_183
timestamp 1586364061
transform 1 0 17940 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_6  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_199
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_208
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_216
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_229
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_228
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23092 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_233
timestamp 1586364061
transform 1 0 22540 0 1 9248
box -38 -48 590 592
use scs8hd_decap_3  FILLER_13_241
timestamp 1586364061
transform 1 0 23276 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_236
timestamp 1586364061
transform 1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_242
timestamp 1586364061
transform 1 0 23368 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_253
timestamp 1586364061
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_263
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_254
timestamp 1586364061
transform 1 0 24472 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_266
timestamp 1586364061
transform 1 0 25576 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_275
timestamp 1586364061
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _091_
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_18
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_29
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_33
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _076_
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_46
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_50
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 222 592
use scs8hd_or3_4  _096_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_54
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_88
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__172__D
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__C
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_93
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_97
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _167_
timestamp 1586364061
transform 1 0 13340 0 1 10336
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 406 592
use scs8hd_nor4_4  _166_
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_150
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 18768 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_188
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20332 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_201
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_205
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 21896 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_218
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_222
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_235
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_243
timestamp 1586364061
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 590 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24288 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_251
timestamp 1586364061
transform 1 0 24196 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_259
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use scs8hd_or3_4  _137_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_9
timestamp 1586364061
transform 1 0 1932 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_12
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_6  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 4968 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_40
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_51
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_62
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use scs8hd_nor4_4  _172_
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _171_
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_112
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__167__D
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_137
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_1  _158_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__D
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_146
timestamp 1586364061
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_157
timestamp 1586364061
transform 1 0 15548 0 -1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _157_
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__165__C
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_161
timestamp 1586364061
transform 1 0 15916 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_184
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_194
timestamp 1586364061
transform 1 0 18952 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_219
timestamp 1586364061
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_222
timestamp 1586364061
transform 1 0 21528 0 -1 11424
box -38 -48 222 592
use scs8hd_conb_1  _196_
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_233
timestamp 1586364061
transform 1 0 22540 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_244
timestamp 1586364061
transform 1 0 23552 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_255
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_267
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_13
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_17
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_30
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _081_
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_47
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _106_
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_55
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _127_
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_92
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_102
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _169_
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 1602 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 16652 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__D
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_161
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_167
timestamp 1586364061
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_180
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_189
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_204
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_213
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_229
timestamp 1586364061
transform 1 0 22172 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_234
timestamp 1586364061
transform 1 0 22632 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_242
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_or3_4  _135_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_6  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 590 592
use scs8hd_or3_4  _104_
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__C
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_49
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_1  _116_
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_8  _125_
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_79
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_18_85
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 590 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 9936 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_109
timestamp 1586364061
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_116
timestamp 1586364061
transform 1 0 11776 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_120
timestamp 1586364061
transform 1 0 12144 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_124
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _168_
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__168__D
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _154_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_157
timestamp 1586364061
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _165_
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_161
timestamp 1586364061
transform 1 0 15916 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_18_182
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_203
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_211
timestamp 1586364061
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_228
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_235
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_247
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 24564 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_259
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_271
timestamp 1586364061
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_1  _126_
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_17
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_19_21
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _105_
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_32
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_28
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_8  _103_
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 866 592
use scs8hd_or3_4  _115_
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_45
timestamp 1586364061
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_49
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_61
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_66
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_77
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_73
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_85
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__C
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 314 592
use scs8hd_buf_1  _079_
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use scs8hd_or3_4  _146_
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_97
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_90
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_96
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 10304 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1050 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_19_113
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_109
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_120
timestamp 1586364061
transform 1 0 12144 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_116
timestamp 1586364061
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_133
timestamp 1586364061
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _160_
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 314 592
use scs8hd_nor4_4  _170_
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__D
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__C
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_162
timestamp 1586364061
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_167
timestamp 1586364061
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_161
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__D
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _164_
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 1602 592
use scs8hd_decap_4  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_188
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18768 0 1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_20_201
timestamp 1586364061
transform 1 0 19596 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_213
timestamp 1586364061
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21896 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_224
timestamp 1586364061
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_228
timestamp 1586364061
transform 1 0 22080 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_235
timestamp 1586364061
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_239
timestamp 1586364061
transform 1 0 23092 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_243
timestamp 1586364061
transform 1 0 23460 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_236
timestamp 1586364061
transform 1 0 22816 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_248
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_260
timestamp 1586364061
transform 1 0 25024 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_20_272
timestamp 1586364061
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_inv_8  _114_
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_44
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_48
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 6256 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_58
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 314 592
use scs8hd_or3_4  _117_
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_80
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_84
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_101
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_134
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 130 592
use scs8hd_nor4_4  _162_
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_149
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_170
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_174
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_178
timestamp 1586364061
transform 1 0 17480 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_195
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20148 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_199
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_203
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_216
timestamp 1586364061
transform 1 0 20976 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_224
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 774 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_1  _082_
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_48
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_54
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_65
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_86
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_90
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_103
timestamp 1586364061
transform 1 0 10580 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_107
timestamp 1586364061
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_122
timestamp 1586364061
transform 1 0 12328 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_128
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_158
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 222 592
use scs8hd_nor4_4  _163_
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 16192 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_162
timestamp 1586364061
transform 1 0 16008 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_191
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_195
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_236
timestamp 1586364061
transform 1 0 22816 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_248
timestamp 1586364061
transform 1 0 23920 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_260
timestamp 1586364061
transform 1 0 25024 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_272
timestamp 1586364061
transform 1 0 26128 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_buf_1  _147_
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_47
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7360 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_83
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_87
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_103
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_107
timestamp 1586364061
transform 1 0 10948 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _107_
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_139
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 406 592
use scs8hd_nor4_4  _161_
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 1602 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_146
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__161__D
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_172
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_176
timestamp 1586364061
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _195_
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_180
timestamp 1586364061
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_191
timestamp 1586364061
transform 1 0 18676 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_195
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20976 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_219
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_223
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_235
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_243
timestamp 1586364061
transform 1 0 23460 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_248
timestamp 1586364061
transform 1 0 23920 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_252
timestamp 1586364061
transform 1 0 24288 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_264
timestamp 1586364061
transform 1 0 25392 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_23_276
timestamp 1586364061
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_61
timestamp 1586364061
transform 1 0 6716 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_87
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 10304 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12144 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_112
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_116
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13708 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_133
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_140
timestamp 1586364061
transform 1 0 13984 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_148
timestamp 1586364061
transform 1 0 14720 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17296 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_172
timestamp 1586364061
transform 1 0 16928 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_185
timestamp 1586364061
transform 1 0 18124 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_189
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 590 592
use scs8hd_decap_8  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 774 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_43
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_46
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_73
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_81
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_94
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_111
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_143
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_154
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_174
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_178
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_210
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_222
timestamp 1586364061
transform 1 0 21528 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_234
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_242
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_1  _118_
timestamp 1586364061
transform 1 0 4140 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_43
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_36
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_47
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 6164 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_83
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_97
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_100
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 10304 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11868 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_109
timestamp 1586364061
transform 1 0 11132 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_119
timestamp 1586364061
transform 1 0 12052 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_130
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_126
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_130
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_126
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_142
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_138
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_137
timestamp 1586364061
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_149
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_153
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_157
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_160
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_165
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_161
timestamp 1586364061
transform 1 0 15916 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_177
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_173
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_177
timestamp 1586364061
transform 1 0 17388 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 866 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17940 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_194
timestamp 1586364061
transform 1 0 18952 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_205
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_205
timestamp 1586364061
transform 1 0 19964 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_217
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_229
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_241
timestamp 1586364061
transform 1 0 23276 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_1  FILLER_28_40
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_50
timestamp 1586364061
transform 1 0 5704 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_73
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_6  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_89
timestamp 1586364061
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_104
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_108
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_112
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_116
timestamp 1586364061
transform 1 0 11776 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_128
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_132
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_6  FILLER_28_157
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_176
timestamp 1586364061
transform 1 0 17296 0 -1 17952
box -38 -48 774 592
use scs8hd_conb_1  _194_
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_187
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_199
timestamp 1586364061
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_28_211
timestamp 1586364061
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_50
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_54
timestamp 1586364061
transform 1 0 6072 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_58
timestamp 1586364061
transform 1 0 6440 0 1 17952
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_73
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_77
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_102
timestamp 1586364061
transform 1 0 10488 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_106
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_134
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_138
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_151
timestamp 1586364061
transform 1 0 14996 0 1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_29_156
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 590 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_173
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_181
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 5888 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_46
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_61
timestamp 1586364061
transform 1 0 6716 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_65
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_78
timestamp 1586364061
transform 1 0 8280 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_87
timestamp 1586364061
transform 1 0 9108 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_119
timestamp 1586364061
transform 1 0 12052 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_136
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_140
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_144
timestamp 1586364061
transform 1 0 14352 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_157
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_169
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_181
timestamp 1586364061
transform 1 0 17756 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_193
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_205
timestamp 1586364061
transform 1 0 19964 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_213
timestamp 1586364061
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_35
timestamp 1586364061
transform 1 0 4324 0 1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 8924 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_73
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_77
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_81
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 10488 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_100
timestamp 1586364061
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_111
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_115
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_119
timestamp 1586364061
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13156 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12972 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_127
timestamp 1586364061
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_142
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_146
timestamp 1586364061
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_47
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_51
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6164 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_66
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_72
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_83
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  FILLER_32_89
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10120 0 -1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_109
timestamp 1586364061
transform 1 0 11132 0 -1 20128
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_126
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_130
timestamp 1586364061
transform 1 0 13064 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_134
timestamp 1586364061
transform 1 0 13432 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_157
timestamp 1586364061
transform 1 0 15548 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_169
timestamp 1586364061
transform 1 0 16652 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_181
timestamp 1586364061
transform 1 0 17756 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_193
timestamp 1586364061
transform 1 0 18860 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_205
timestamp 1586364061
transform 1 0 19964 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 774 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 5612 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 4784 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_42
timestamp 1586364061
transform 1 0 4968 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_46
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_62
timestamp 1586364061
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_58
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6624 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_68
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_79
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_83
timestamp 1586364061
transform 1 0 8740 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_75
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_8  FILLER_34_83
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_91
timestamp 1586364061
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_96
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_102
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_102
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10304 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_107
timestamp 1586364061
transform 1 0 10948 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_106
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12604 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_136
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_140
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_138
timestamp 1586364061
transform 1 0 13800 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_150
timestamp 1586364061
transform 1 0 14904 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_146
timestamp 1586364061
transform 1 0 14536 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_157
timestamp 1586364061
transform 1 0 15548 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_153
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use scs8hd_conb_1  _198_
timestamp 1586364061
transform 1 0 15916 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_164
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_176
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_163
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_167
timestamp 1586364061
transform 1 0 16468 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_182
timestamp 1586364061
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_179
timestamp 1586364061
transform 1 0 17572 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_191
timestamp 1586364061
transform 1 0 18676 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_203
timestamp 1586364061
transform 1 0 19780 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_211
timestamp 1586364061
transform 1 0 20516 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_35_35
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 130 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_38
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_42
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_73
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_78
timestamp 1586364061
transform 1 0 8280 0 1 21216
box -38 -48 314 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_90
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_102
timestamp 1586364061
transform 1 0 10488 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_134
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_138
timestamp 1586364061
transform 1 0 13800 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 15272 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_151
timestamp 1586364061
transform 1 0 14996 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__219__A
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_173
timestamp 1586364061
transform 1 0 17020 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_181
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 774 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 4784 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 5796 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_49
timestamp 1586364061
transform 1 0 5612 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_53
timestamp 1586364061
transform 1 0 5980 0 -1 22304
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_72
timestamp 1586364061
transform 1 0 7728 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_79
timestamp 1586364061
transform 1 0 8372 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_83
timestamp 1586364061
transform 1 0 8740 0 -1 22304
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10304 0 -1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_91
timestamp 1586364061
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_99
timestamp 1586364061
transform 1 0 10212 0 -1 22304
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12512 0 -1 22304
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_36_111
timestamp 1586364061
transform 1 0 11316 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_123
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_135
timestamp 1586364061
transform 1 0 13524 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_140
timestamp 1586364061
transform 1 0 13984 0 -1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_144
timestamp 1586364061
transform 1 0 14352 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_148
timestamp 1586364061
transform 1 0 14720 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_152
timestamp 1586364061
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_2  _219_
timestamp 1586364061
transform 1 0 16836 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_163
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_167
timestamp 1586364061
transform 1 0 16468 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_175
timestamp 1586364061
transform 1 0 17204 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_187
timestamp 1586364061
transform 1 0 18308 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_199
timestamp 1586364061
transform 1 0 19412 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_36_211
timestamp 1586364061
transform 1 0 20516 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_37_47
timestamp 1586364061
transform 1 0 5428 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_50
timestamp 1586364061
transform 1 0 5704 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_54
timestamp 1586364061
transform 1 0 6072 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_58
timestamp 1586364061
transform 1 0 6440 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_67
timestamp 1586364061
transform 1 0 7268 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_79
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_89
timestamp 1586364061
transform 1 0 9292 0 1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9476 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_104
timestamp 1586364061
transform 1 0 10672 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_108
timestamp 1586364061
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_112
timestamp 1586364061
transform 1 0 11408 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_116
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13800 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_126
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_134
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_37_158
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16376 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_162
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_169
timestamp 1586364061
transform 1 0 16652 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_173
timestamp 1586364061
transform 1 0 17020 0 1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_37_178
timestamp 1586364061
transform 1 0 17480 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_182
timestamp 1586364061
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5520 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_46
timestamp 1586364061
transform 1 0 5336 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_57
timestamp 1586364061
transform 1 0 6348 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_61
timestamp 1586364061
transform 1 0 6716 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_74
timestamp 1586364061
transform 1 0 7912 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_38_86
timestamp 1586364061
transform 1 0 9016 0 -1 23392
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10120 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_97
timestamp 1586364061
transform 1 0 10028 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_101
timestamp 1586364061
transform 1 0 10396 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11132 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_118
timestamp 1586364061
transform 1 0 11960 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_122
timestamp 1586364061
transform 1 0 12328 0 -1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_125
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_135
timestamp 1586364061
transform 1 0 13524 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_38_157
timestamp 1586364061
transform 1 0 15548 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_168
timestamp 1586364061
transform 1 0 16560 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_179
timestamp 1586364061
transform 1 0 17572 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_191
timestamp 1586364061
transform 1 0 18676 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_203
timestamp 1586364061
transform 1 0 19780 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_211
timestamp 1586364061
transform 1 0 20516 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_17
timestamp 1586364061
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_6
timestamp 1586364061
transform 1 0 1656 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_21
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_18
timestamp 1586364061
transform 1 0 2760 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_30
timestamp 1586364061
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_6  FILLER_40_38
timestamp 1586364061
transform 1 0 4600 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_40
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_36
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_49
timestamp 1586364061
transform 1 0 5612 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 23392
box -38 -48 866 592
use scs8hd_decap_4  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_71
timestamp 1586364061
transform 1 0 7636 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_40_66
timestamp 1586364061
transform 1 0 7176 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_78
timestamp 1586364061
transform 1 0 8280 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8464 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_88
timestamp 1586364061
transform 1 0 9200 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_89
timestamp 1586364061
transform 1 0 9292 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_82
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_96
timestamp 1586364061
transform 1 0 9936 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_93
timestamp 1586364061
transform 1 0 9660 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_conb_1  _199_
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_100
timestamp 1586364061
transform 1 0 10304 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_119
timestamp 1586364061
transform 1 0 12052 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_113
timestamp 1586364061
transform 1 0 11500 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_40_125
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_142
timestamp 1586364061
transform 1 0 14168 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_40_136
timestamp 1586364061
transform 1 0 13616 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_136
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 23392
box -38 -48 866 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_149
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_153
timestamp 1586364061
transform 1 0 15180 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_156
timestamp 1586364061
transform 1 0 15456 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_150
timestamp 1586364061
transform 1 0 14904 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_157
timestamp 1586364061
transform 1 0 15548 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _218_
timestamp 1586364061
transform 1 0 16284 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _225_
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 16284 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__218__A
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_163
timestamp 1586364061
transform 1 0 16100 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_167
timestamp 1586364061
transform 1 0 16468 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_169
timestamp 1586364061
transform 1 0 16652 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_40_181
timestamp 1586364061
transform 1 0 17756 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_187
timestamp 1586364061
transform 1 0 18308 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 314 592
use scs8hd_buf_2  _224_
timestamp 1586364061
transform 1 0 18032 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_191
timestamp 1586364061
transform 1 0 18676 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 18492 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _223_
timestamp 1586364061
transform 1 0 19044 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_188
timestamp 1586364061
transform 1 0 18400 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 19596 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_199
timestamp 1586364061
transform 1 0 19412 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_203
timestamp 1586364061
transform 1 0 19780 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_200
timestamp 1586364061
transform 1 0 19504 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_40_212
timestamp 1586364061
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use scs8hd_buf_2  _220_
timestamp 1586364061
transform 1 0 22172 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _221_
timestamp 1586364061
transform 1 0 21068 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__221__A
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_215
timestamp 1586364061
transform 1 0 20884 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_221
timestamp 1586364061
transform 1 0 21436 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_225
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__220__A
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_233
timestamp 1586364061
transform 1 0 22540 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_237
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5244 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_41_48
timestamp 1586364061
transform 1 0 5520 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_52
timestamp 1586364061
transform 1 0 5888 0 1 24480
box -38 -48 774 592
use scs8hd_conb_1  _197_
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_60
timestamp 1586364061
transform 1 0 6624 0 1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_41_65
timestamp 1586364061
transform 1 0 7084 0 1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8004 0 1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_73
timestamp 1586364061
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_78
timestamp 1586364061
transform 1 0 8280 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_82
timestamp 1586364061
transform 1 0 8648 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_95
timestamp 1586364061
transform 1 0 9844 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_99
timestamp 1586364061
transform 1 0 10212 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_41_112
timestamp 1586364061
transform 1 0 11408 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_120
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _222_
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_127
timestamp 1586364061
transform 1 0 12788 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_131
timestamp 1586364061
transform 1 0 13156 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_136
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_140
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_152
timestamp 1586364061
transform 1 0 15088 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_158
timestamp 1586364061
transform 1 0 15640 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_162
timestamp 1586364061
transform 1 0 16008 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_174
timestamp 1586364061
transform 1 0 17112 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_182
timestamp 1586364061
transform 1 0 17848 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_103
timestamp 1586364061
transform 1 0 10580 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_107
timestamp 1586364061
transform 1 0 10948 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_119
timestamp 1586364061
transform 1 0 12052 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_123
timestamp 1586364061
transform 1 0 12420 0 -1 25568
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_128
timestamp 1586364061
transform 1 0 12880 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_140
timestamp 1586364061
transform 1 0 13984 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_42_152
timestamp 1586364061
transform 1 0 15088 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 4496 480 4616 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 7624 480 7744 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 10752 480 10872 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 13880 480 14000 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 17008 480 17128 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 20136 480 20256 6 address[5]
port 5 nsew default input
rlabel metal3 s 0 23264 480 23384 6 address[6]
port 6 nsew default input
rlabel metal2 s 5630 0 5686 480 6 bottom_left_grid_pin_11_
port 7 nsew default input
rlabel metal2 s 6642 0 6698 480 6 bottom_left_grid_pin_13_
port 8 nsew default input
rlabel metal2 s 7654 0 7710 480 6 bottom_left_grid_pin_15_
port 9 nsew default input
rlabel metal2 s 478 0 534 480 6 bottom_left_grid_pin_1_
port 10 nsew default input
rlabel metal2 s 1490 0 1546 480 6 bottom_left_grid_pin_3_
port 11 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_5_
port 12 nsew default input
rlabel metal2 s 3514 0 3570 480 6 bottom_left_grid_pin_7_
port 13 nsew default input
rlabel metal2 s 4618 0 4674 480 6 bottom_left_grid_pin_9_
port 14 nsew default input
rlabel metal2 s 27342 0 27398 480 6 bottom_right_grid_pin_11_
port 15 nsew default input
rlabel metal3 s 27520 14696 28000 14816 6 chanx_right_in[0]
port 16 nsew default input
rlabel metal3 s 27520 16056 28000 16176 6 chanx_right_in[1]
port 17 nsew default input
rlabel metal3 s 27520 17416 28000 17536 6 chanx_right_in[2]
port 18 nsew default input
rlabel metal3 s 27520 18776 28000 18896 6 chanx_right_in[3]
port 19 nsew default input
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_in[4]
port 20 nsew default input
rlabel metal3 s 27520 21632 28000 21752 6 chanx_right_in[5]
port 21 nsew default input
rlabel metal3 s 27520 22992 28000 23112 6 chanx_right_in[6]
port 22 nsew default input
rlabel metal3 s 27520 24488 28000 24608 6 chanx_right_in[7]
port 23 nsew default input
rlabel metal3 s 27520 25848 28000 25968 6 chanx_right_in[8]
port 24 nsew default input
rlabel metal3 s 27520 2048 28000 2168 6 chanx_right_out[0]
port 25 nsew default tristate
rlabel metal3 s 27520 3408 28000 3528 6 chanx_right_out[1]
port 26 nsew default tristate
rlabel metal3 s 27520 4768 28000 4888 6 chanx_right_out[2]
port 27 nsew default tristate
rlabel metal3 s 27520 6264 28000 6384 6 chanx_right_out[3]
port 28 nsew default tristate
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_out[4]
port 29 nsew default tristate
rlabel metal3 s 27520 8984 28000 9104 6 chanx_right_out[5]
port 30 nsew default tristate
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_out[6]
port 31 nsew default tristate
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_out[7]
port 32 nsew default tristate
rlabel metal3 s 27520 13200 28000 13320 6 chanx_right_out[8]
port 33 nsew default tristate
rlabel metal2 s 8758 0 8814 480 6 chany_bottom_in[0]
port 34 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[1]
port 35 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[2]
port 36 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[3]
port 37 nsew default input
rlabel metal2 s 12898 0 12954 480 6 chany_bottom_in[4]
port 38 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[5]
port 39 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[6]
port 40 nsew default input
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_in[7]
port 41 nsew default input
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_in[8]
port 42 nsew default input
rlabel metal2 s 18050 0 18106 480 6 chany_bottom_out[0]
port 43 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 chany_bottom_out[1]
port 44 nsew default tristate
rlabel metal2 s 20074 0 20130 480 6 chany_bottom_out[2]
port 45 nsew default tristate
rlabel metal2 s 21178 0 21234 480 6 chany_bottom_out[3]
port 46 nsew default tristate
rlabel metal2 s 22190 0 22246 480 6 chany_bottom_out[4]
port 47 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_bottom_out[5]
port 48 nsew default tristate
rlabel metal2 s 24214 0 24270 480 6 chany_bottom_out[6]
port 49 nsew default tristate
rlabel metal2 s 25318 0 25374 480 6 chany_bottom_out[7]
port 50 nsew default tristate
rlabel metal2 s 26330 0 26386 480 6 chany_bottom_out[8]
port 51 nsew default tristate
rlabel metal2 s 8758 27520 8814 28000 6 chany_top_in[0]
port 52 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 10782 27520 10838 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 11794 27520 11850 28000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 12898 27520 12954 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 14922 27520 14978 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 17038 27520 17094 28000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 18050 27520 18106 28000 6 chany_top_out[0]
port 61 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[1]
port 62 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[2]
port 63 nsew default tristate
rlabel metal2 s 21178 27520 21234 28000 6 chany_top_out[3]
port 64 nsew default tristate
rlabel metal2 s 22190 27520 22246 28000 6 chany_top_out[4]
port 65 nsew default tristate
rlabel metal2 s 23202 27520 23258 28000 6 chany_top_out[5]
port 66 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[6]
port 67 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[7]
port 68 nsew default tristate
rlabel metal2 s 26330 27520 26386 28000 6 chany_top_out[8]
port 69 nsew default tristate
rlabel metal3 s 0 26392 480 26512 6 data_in
port 70 nsew default input
rlabel metal3 s 0 1504 480 1624 6 enable
port 71 nsew default input
rlabel metal3 s 27520 688 28000 808 6 right_bottom_grid_pin_12_
port 72 nsew default input
rlabel metal3 s 27520 27208 28000 27328 6 right_top_grid_pin_10_
port 73 nsew default input
rlabel metal2 s 5630 27520 5686 28000 6 top_left_grid_pin_11_
port 74 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 top_left_grid_pin_13_
port 75 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 top_left_grid_pin_15_
port 76 nsew default input
rlabel metal2 s 478 27520 534 28000 6 top_left_grid_pin_1_
port 77 nsew default input
rlabel metal2 s 1490 27520 1546 28000 6 top_left_grid_pin_3_
port 78 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_5_
port 79 nsew default input
rlabel metal2 s 3514 27520 3570 28000 6 top_left_grid_pin_7_
port 80 nsew default input
rlabel metal2 s 4618 27520 4674 28000 6 top_left_grid_pin_9_
port 81 nsew default input
rlabel metal2 s 27342 27520 27398 28000 6 top_right_grid_pin_11_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
