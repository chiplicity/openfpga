magic
tech sky130A
magscale 1 2
timestamp 1605198538
<< locali >>
rect 6929 20247 6963 20349
rect 10517 16575 10551 16745
rect 12265 12631 12299 12801
rect 12265 12087 12299 12393
rect 9137 7327 9171 7497
rect 9689 5763 9723 5865
rect 9631 3553 9815 3587
rect 9781 3519 9815 3553
rect 12633 2295 12667 2465
rect 13737 1683 13771 2057
<< viali >>
rect 14473 20553 14507 20587
rect 15761 20553 15795 20587
rect 7205 20485 7239 20519
rect 1409 20417 1443 20451
rect 2973 20417 3007 20451
rect 5641 20417 5675 20451
rect 8677 20417 8711 20451
rect 11253 20417 11287 20451
rect 13277 20417 13311 20451
rect 17141 20417 17175 20451
rect 17325 20417 17359 20451
rect 19625 20417 19659 20451
rect 2881 20349 2915 20383
rect 6929 20349 6963 20383
rect 7027 20349 7061 20383
rect 13093 20349 13127 20383
rect 14289 20349 14323 20383
rect 15577 20349 15611 20383
rect 19441 20349 19475 20383
rect 5549 20281 5583 20315
rect 11161 20281 11195 20315
rect 17049 20281 17083 20315
rect 2421 20213 2455 20247
rect 2789 20213 2823 20247
rect 4077 20213 4111 20247
rect 5089 20213 5123 20247
rect 5457 20213 5491 20247
rect 6929 20213 6963 20247
rect 8125 20213 8159 20247
rect 8493 20213 8527 20247
rect 8585 20213 8619 20247
rect 10701 20213 10735 20247
rect 11069 20213 11103 20247
rect 12633 20213 12667 20247
rect 13001 20213 13035 20247
rect 16681 20213 16715 20247
rect 18981 20213 19015 20247
rect 19349 20213 19383 20247
rect 4353 20009 4387 20043
rect 4721 20009 4755 20043
rect 6285 20009 6319 20043
rect 8033 20009 8067 20043
rect 12265 20009 12299 20043
rect 13461 20009 13495 20043
rect 17049 20009 17083 20043
rect 2789 19941 2823 19975
rect 8401 19941 8435 19975
rect 12357 19941 12391 19975
rect 15577 19941 15611 19975
rect 2881 19873 2915 19907
rect 9956 19873 9990 19907
rect 13829 19873 13863 19907
rect 15301 19873 15335 19907
rect 18245 19873 18279 19907
rect 19625 19873 19659 19907
rect 1409 19805 1443 19839
rect 3065 19805 3099 19839
rect 4813 19805 4847 19839
rect 4905 19805 4939 19839
rect 6377 19805 6411 19839
rect 6561 19805 6595 19839
rect 8493 19805 8527 19839
rect 8677 19805 8711 19839
rect 9689 19805 9723 19839
rect 12449 19805 12483 19839
rect 13921 19805 13955 19839
rect 14013 19805 14047 19839
rect 17141 19805 17175 19839
rect 17325 19805 17359 19839
rect 19717 19805 19751 19839
rect 19901 19805 19935 19839
rect 2421 19737 2455 19771
rect 5917 19669 5951 19703
rect 11069 19669 11103 19703
rect 11897 19669 11931 19703
rect 16681 19669 16715 19703
rect 19257 19669 19291 19703
rect 16957 19465 16991 19499
rect 8585 19397 8619 19431
rect 2421 19329 2455 19363
rect 3341 19329 3375 19363
rect 7389 19329 7423 19363
rect 19349 19329 19383 19363
rect 19533 19329 19567 19363
rect 5641 19261 5675 19295
rect 7297 19261 7331 19295
rect 8401 19261 8435 19295
rect 9505 19261 9539 19295
rect 13369 19261 13403 19295
rect 15577 19261 15611 19295
rect 19257 19261 19291 19295
rect 20545 19261 20579 19295
rect 3586 19193 3620 19227
rect 9772 19193 9806 19227
rect 13636 19193 13670 19227
rect 15822 19193 15856 19227
rect 1777 19125 1811 19159
rect 2145 19125 2179 19159
rect 2237 19125 2271 19159
rect 4721 19125 4755 19159
rect 5825 19125 5859 19159
rect 6837 19125 6871 19159
rect 7205 19125 7239 19159
rect 10885 19125 10919 19159
rect 14749 19125 14783 19159
rect 18889 19125 18923 19159
rect 20729 19125 20763 19159
rect 1409 18921 1443 18955
rect 2789 18921 2823 18955
rect 4537 18921 4571 18955
rect 6745 18921 6779 18955
rect 7849 18921 7883 18955
rect 8309 18921 8343 18955
rect 10701 18921 10735 18955
rect 15301 18921 15335 18955
rect 17693 18921 17727 18955
rect 6653 18853 6687 18887
rect 10609 18853 10643 18887
rect 18766 18853 18800 18887
rect 2881 18785 2915 18819
rect 4445 18785 4479 18819
rect 8217 18785 8251 18819
rect 12061 18785 12095 18819
rect 14105 18785 14139 18819
rect 16313 18785 16347 18819
rect 16580 18785 16614 18819
rect 18521 18785 18555 18819
rect 3065 18717 3099 18751
rect 4721 18717 4755 18751
rect 6837 18717 6871 18751
rect 8401 18717 8435 18751
rect 10793 18717 10827 18751
rect 11805 18717 11839 18751
rect 2421 18649 2455 18683
rect 13185 18649 13219 18683
rect 4077 18581 4111 18615
rect 6285 18581 6319 18615
rect 10241 18581 10275 18615
rect 14289 18581 14323 18615
rect 19901 18581 19935 18615
rect 4721 18377 4755 18411
rect 12449 18377 12483 18411
rect 16405 18377 16439 18411
rect 14013 18309 14047 18343
rect 2237 18241 2271 18275
rect 2421 18241 2455 18275
rect 3341 18241 3375 18275
rect 6837 18241 6871 18275
rect 13093 18241 13127 18275
rect 14657 18241 14691 18275
rect 16957 18241 16991 18275
rect 18797 18241 18831 18275
rect 2145 18173 2179 18207
rect 5549 18173 5583 18207
rect 9413 18173 9447 18207
rect 9680 18173 9714 18207
rect 19064 18173 19098 18207
rect 3586 18105 3620 18139
rect 7093 18105 7127 18139
rect 12817 18105 12851 18139
rect 14473 18105 14507 18139
rect 16773 18105 16807 18139
rect 1777 18037 1811 18071
rect 5733 18037 5767 18071
rect 8217 18037 8251 18071
rect 10793 18037 10827 18071
rect 12909 18037 12943 18071
rect 14381 18037 14415 18071
rect 16865 18037 16899 18071
rect 20177 18037 20211 18071
rect 2421 17833 2455 17867
rect 5825 17833 5859 17867
rect 9689 17833 9723 17867
rect 10149 17833 10183 17867
rect 13001 17833 13035 17867
rect 15669 17833 15703 17867
rect 19717 17833 19751 17867
rect 4712 17765 4746 17799
rect 6920 17765 6954 17799
rect 14105 17765 14139 17799
rect 15761 17765 15795 17799
rect 18153 17765 18187 17799
rect 2789 17697 2823 17731
rect 10057 17697 10091 17731
rect 11888 17697 11922 17731
rect 13829 17697 13863 17731
rect 18061 17697 18095 17731
rect 19625 17697 19659 17731
rect 1409 17629 1443 17663
rect 2881 17629 2915 17663
rect 3065 17629 3099 17663
rect 4445 17629 4479 17663
rect 6653 17629 6687 17663
rect 10241 17629 10275 17663
rect 11621 17629 11655 17663
rect 15853 17629 15887 17663
rect 18337 17629 18371 17663
rect 19809 17629 19843 17663
rect 15301 17561 15335 17595
rect 8033 17493 8067 17527
rect 17693 17493 17727 17527
rect 19257 17493 19291 17527
rect 3709 17289 3743 17323
rect 4537 17289 4571 17323
rect 20453 17289 20487 17323
rect 8309 17221 8343 17255
rect 16221 17221 16255 17255
rect 2329 17153 2363 17187
rect 5089 17153 5123 17187
rect 8769 17153 8803 17187
rect 8953 17153 8987 17187
rect 10701 17153 10735 17187
rect 13093 17153 13127 17187
rect 16681 17153 16715 17187
rect 16773 17153 16807 17187
rect 18061 17153 18095 17187
rect 19073 17153 19107 17187
rect 4905 17085 4939 17119
rect 7021 17085 7055 17119
rect 14013 17085 14047 17119
rect 19340 17085 19374 17119
rect 2596 17017 2630 17051
rect 7297 17017 7331 17051
rect 8677 17017 8711 17051
rect 10517 17017 10551 17051
rect 12909 17017 12943 17051
rect 14258 17017 14292 17051
rect 4997 16949 5031 16983
rect 10057 16949 10091 16983
rect 10425 16949 10459 16983
rect 12449 16949 12483 16983
rect 12817 16949 12851 16983
rect 15393 16949 15427 16983
rect 16589 16949 16623 16983
rect 2421 16745 2455 16779
rect 8677 16745 8711 16779
rect 10517 16745 10551 16779
rect 11989 16745 12023 16779
rect 12817 16745 12851 16779
rect 13277 16745 13311 16779
rect 18797 16745 18831 16779
rect 19165 16745 19199 16779
rect 2789 16677 2823 16711
rect 5733 16677 5767 16711
rect 1409 16609 1443 16643
rect 1685 16609 1719 16643
rect 4077 16609 4111 16643
rect 4353 16609 4387 16643
rect 7297 16609 7331 16643
rect 8493 16609 8527 16643
rect 19257 16677 19291 16711
rect 10865 16609 10899 16643
rect 13185 16609 13219 16643
rect 16037 16609 16071 16643
rect 16304 16609 16338 16643
rect 2881 16541 2915 16575
rect 3065 16541 3099 16575
rect 5825 16541 5859 16575
rect 6009 16541 6043 16575
rect 7389 16541 7423 16575
rect 7481 16541 7515 16575
rect 10517 16541 10551 16575
rect 10609 16541 10643 16575
rect 13369 16541 13403 16575
rect 19349 16541 19383 16575
rect 17417 16473 17451 16507
rect 5365 16405 5399 16439
rect 6929 16405 6963 16439
rect 3065 16201 3099 16235
rect 10425 16201 10459 16235
rect 9597 16133 9631 16167
rect 5181 16065 5215 16099
rect 10885 16065 10919 16099
rect 10977 16065 11011 16099
rect 15761 16065 15795 16099
rect 1685 15997 1719 16031
rect 4997 15997 5031 16031
rect 6929 15997 6963 16031
rect 8217 15997 8251 16031
rect 8484 15997 8518 16031
rect 13369 15997 13403 16031
rect 13636 15997 13670 16031
rect 18521 15997 18555 16031
rect 18788 15997 18822 16031
rect 1952 15929 1986 15963
rect 5089 15929 5123 15963
rect 7205 15929 7239 15963
rect 10793 15929 10827 15963
rect 16028 15929 16062 15963
rect 4629 15861 4663 15895
rect 14749 15861 14783 15895
rect 17141 15861 17175 15895
rect 19901 15861 19935 15895
rect 2881 15657 2915 15691
rect 8677 15657 8711 15691
rect 9689 15657 9723 15691
rect 10057 15657 10091 15691
rect 11253 15657 11287 15691
rect 11713 15657 11747 15691
rect 14381 15657 14415 15691
rect 19717 15657 19751 15691
rect 1409 15589 1443 15623
rect 1777 15589 1811 15623
rect 6736 15589 6770 15623
rect 13277 15589 13311 15623
rect 2789 15521 2823 15555
rect 4077 15521 4111 15555
rect 4344 15521 4378 15555
rect 6469 15521 6503 15555
rect 8861 15521 8895 15555
rect 11621 15521 11655 15555
rect 13185 15521 13219 15555
rect 14565 15521 14599 15555
rect 16488 15521 16522 15555
rect 19625 15521 19659 15555
rect 3065 15453 3099 15487
rect 10149 15453 10183 15487
rect 10333 15453 10367 15487
rect 11805 15453 11839 15487
rect 13461 15453 13495 15487
rect 16221 15453 16255 15487
rect 19901 15453 19935 15487
rect 7849 15385 7883 15419
rect 2421 15317 2455 15351
rect 5457 15317 5491 15351
rect 12817 15317 12851 15351
rect 17601 15317 17635 15351
rect 19257 15317 19291 15351
rect 3341 15113 3375 15147
rect 6469 15113 6503 15147
rect 14749 15113 14783 15147
rect 16313 15113 16347 15147
rect 10333 15045 10367 15079
rect 13921 15045 13955 15079
rect 2421 14977 2455 15011
rect 3893 14977 3927 15011
rect 5457 14977 5491 15011
rect 7389 14977 7423 15011
rect 8953 14977 8987 15011
rect 12541 14977 12575 15011
rect 15301 14977 15335 15011
rect 16865 14977 16899 15011
rect 2145 14909 2179 14943
rect 6653 14909 6687 14943
rect 7297 14909 7331 14943
rect 9220 14909 9254 14943
rect 11253 14909 11287 14943
rect 15209 14909 15243 14943
rect 18889 14909 18923 14943
rect 19156 14909 19190 14943
rect 2237 14841 2271 14875
rect 7205 14841 7239 14875
rect 12808 14841 12842 14875
rect 15117 14841 15151 14875
rect 16681 14841 16715 14875
rect 1777 14773 1811 14807
rect 3709 14773 3743 14807
rect 3801 14773 3835 14807
rect 4905 14773 4939 14807
rect 5273 14773 5307 14807
rect 5365 14773 5399 14807
rect 6837 14773 6871 14807
rect 11437 14773 11471 14807
rect 16773 14773 16807 14807
rect 20269 14773 20303 14807
rect 2881 14569 2915 14603
rect 4077 14569 4111 14603
rect 14289 14569 14323 14603
rect 15301 14569 15335 14603
rect 19625 14569 19659 14603
rect 6368 14501 6402 14535
rect 2789 14433 2823 14467
rect 4445 14433 4479 14467
rect 4537 14433 4571 14467
rect 6101 14433 6135 14467
rect 8309 14433 8343 14467
rect 9689 14433 9723 14467
rect 9956 14433 9990 14467
rect 12164 14433 12198 14467
rect 14105 14433 14139 14467
rect 16313 14433 16347 14467
rect 16580 14433 16614 14467
rect 18705 14433 18739 14467
rect 1409 14365 1443 14399
rect 3065 14365 3099 14399
rect 4721 14365 4755 14399
rect 8585 14365 8619 14399
rect 11897 14365 11931 14399
rect 19717 14365 19751 14399
rect 19901 14365 19935 14399
rect 13277 14297 13311 14331
rect 17693 14297 17727 14331
rect 2421 14229 2455 14263
rect 7481 14229 7515 14263
rect 11069 14229 11103 14263
rect 18521 14229 18555 14263
rect 19257 14229 19291 14263
rect 1777 14025 1811 14059
rect 8217 14025 8251 14059
rect 9045 14025 9079 14059
rect 14013 14025 14047 14059
rect 15577 14025 15611 14059
rect 4721 13957 4755 13991
rect 5733 13957 5767 13991
rect 10793 13957 10827 13991
rect 12449 13957 12483 13991
rect 2421 13889 2455 13923
rect 6837 13889 6871 13923
rect 9505 13889 9539 13923
rect 9689 13889 9723 13923
rect 11345 13889 11379 13923
rect 13093 13889 13127 13923
rect 14565 13889 14599 13923
rect 17049 13889 17083 13923
rect 2237 13821 2271 13855
rect 3341 13821 3375 13855
rect 5549 13821 5583 13855
rect 7104 13821 7138 13855
rect 12909 13821 12943 13855
rect 15761 13821 15795 13855
rect 16865 13821 16899 13855
rect 18797 13821 18831 13855
rect 19064 13821 19098 13855
rect 2145 13753 2179 13787
rect 3586 13753 3620 13787
rect 9413 13753 9447 13787
rect 11161 13753 11195 13787
rect 11253 13753 11287 13787
rect 14473 13753 14507 13787
rect 12817 13685 12851 13719
rect 14381 13685 14415 13719
rect 16405 13685 16439 13719
rect 16773 13685 16807 13719
rect 20177 13685 20211 13719
rect 4445 13481 4479 13515
rect 5641 13481 5675 13515
rect 6101 13481 6135 13515
rect 7481 13481 7515 13515
rect 8033 13481 8067 13515
rect 10149 13481 10183 13515
rect 16589 13481 16623 13515
rect 6009 13413 6043 13447
rect 11520 13413 11554 13447
rect 13829 13413 13863 13447
rect 1777 13345 1811 13379
rect 2044 13345 2078 13379
rect 4537 13345 4571 13379
rect 7665 13345 7699 13379
rect 8401 13345 8435 13379
rect 10057 13345 10091 13379
rect 13921 13345 13955 13379
rect 16497 13345 16531 13379
rect 17693 13345 17727 13379
rect 17960 13345 17994 13379
rect 4629 13277 4663 13311
rect 6285 13277 6319 13311
rect 8493 13277 8527 13311
rect 8677 13277 8711 13311
rect 10241 13277 10275 13311
rect 11253 13277 11287 13311
rect 14013 13277 14047 13311
rect 16773 13277 16807 13311
rect 3157 13141 3191 13175
rect 4077 13141 4111 13175
rect 9689 13141 9723 13175
rect 12633 13141 12667 13175
rect 13461 13141 13495 13175
rect 16129 13141 16163 13175
rect 19073 13141 19107 13175
rect 6837 12937 6871 12971
rect 9873 12937 9907 12971
rect 10701 12937 10735 12971
rect 17141 12937 17175 12971
rect 20729 12937 20763 12971
rect 2881 12801 2915 12835
rect 5641 12801 5675 12835
rect 7297 12801 7331 12835
rect 7389 12801 7423 12835
rect 11253 12801 11287 12835
rect 12265 12801 12299 12835
rect 13001 12801 13035 12835
rect 14565 12801 14599 12835
rect 15761 12801 15795 12835
rect 1593 12733 1627 12767
rect 3148 12733 3182 12767
rect 5457 12733 5491 12767
rect 5549 12733 5583 12767
rect 8493 12733 8527 12767
rect 8760 12733 8794 12767
rect 11069 12733 11103 12767
rect 1869 12665 1903 12699
rect 7205 12665 7239 12699
rect 16028 12733 16062 12767
rect 18061 12733 18095 12767
rect 19349 12733 19383 12767
rect 12909 12665 12943 12699
rect 14473 12665 14507 12699
rect 18337 12665 18371 12699
rect 19616 12665 19650 12699
rect 4261 12597 4295 12631
rect 5089 12597 5123 12631
rect 11161 12597 11195 12631
rect 12265 12597 12299 12631
rect 12449 12597 12483 12631
rect 12817 12597 12851 12631
rect 14013 12597 14047 12631
rect 14381 12597 14415 12631
rect 2697 12393 2731 12427
rect 6285 12393 6319 12427
rect 8033 12393 8067 12427
rect 12265 12393 12299 12427
rect 5172 12325 5206 12359
rect 8401 12325 8435 12359
rect 9956 12325 9990 12359
rect 2605 12257 2639 12291
rect 4905 12257 4939 12291
rect 7941 12257 7975 12291
rect 9689 12257 9723 12291
rect 2881 12189 2915 12223
rect 8493 12189 8527 12223
rect 8585 12189 8619 12223
rect 2237 12121 2271 12155
rect 7757 12121 7791 12155
rect 15761 12325 15795 12359
rect 17509 12325 17543 12359
rect 12633 12257 12667 12291
rect 13084 12257 13118 12291
rect 15669 12257 15703 12291
rect 16129 12257 16163 12291
rect 17417 12257 17451 12291
rect 18613 12257 18647 12291
rect 18869 12257 18903 12291
rect 12817 12189 12851 12223
rect 15853 12189 15887 12223
rect 17693 12189 17727 12223
rect 12449 12121 12483 12155
rect 11069 12053 11103 12087
rect 12265 12053 12299 12087
rect 14197 12053 14231 12087
rect 14841 12053 14875 12087
rect 15301 12053 15335 12087
rect 17049 12053 17083 12087
rect 19993 12053 20027 12087
rect 2237 11849 2271 11883
rect 3801 11849 3835 11883
rect 9321 11849 9355 11883
rect 13829 11849 13863 11883
rect 16405 11849 16439 11883
rect 19625 11849 19659 11883
rect 11529 11781 11563 11815
rect 2697 11713 2731 11747
rect 2881 11713 2915 11747
rect 4353 11713 4387 11747
rect 5733 11713 5767 11747
rect 9965 11713 9999 11747
rect 15209 11713 15243 11747
rect 16957 11713 16991 11747
rect 18705 11713 18739 11747
rect 20269 11713 20303 11747
rect 2605 11645 2639 11679
rect 5457 11645 5491 11679
rect 7021 11645 7055 11679
rect 7288 11645 7322 11679
rect 10149 11645 10183 11679
rect 10416 11645 10450 11679
rect 12449 11645 12483 11679
rect 15025 11645 15059 11679
rect 18429 11645 18463 11679
rect 4169 11577 4203 11611
rect 9689 11577 9723 11611
rect 12716 11577 12750 11611
rect 15117 11577 15151 11611
rect 16773 11577 16807 11611
rect 19993 11577 20027 11611
rect 4261 11509 4295 11543
rect 8401 11509 8435 11543
rect 9781 11509 9815 11543
rect 11621 11509 11655 11543
rect 14657 11509 14691 11543
rect 16865 11509 16899 11543
rect 18061 11509 18095 11543
rect 18521 11509 18555 11543
rect 19533 11509 19567 11543
rect 20085 11509 20119 11543
rect 6745 11305 6779 11339
rect 7941 11305 7975 11339
rect 11805 11305 11839 11339
rect 15669 11305 15703 11339
rect 18705 11305 18739 11339
rect 12725 11237 12759 11271
rect 14197 11237 14231 11271
rect 15761 11237 15795 11271
rect 17570 11237 17604 11271
rect 1409 11169 1443 11203
rect 2789 11169 2823 11203
rect 4077 11169 4111 11203
rect 4353 11169 4387 11203
rect 5632 11169 5666 11203
rect 9321 11169 9355 11203
rect 10517 11169 10551 11203
rect 12817 11169 12851 11203
rect 13921 11169 13955 11203
rect 19533 11169 19567 11203
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 5365 11101 5399 11135
rect 8033 11101 8067 11135
rect 8125 11101 8159 11135
rect 13001 11101 13035 11135
rect 15853 11101 15887 11135
rect 17325 11101 17359 11135
rect 19809 11101 19843 11135
rect 12357 11033 12391 11067
rect 15301 11033 15335 11067
rect 2421 10965 2455 10999
rect 7573 10965 7607 10999
rect 9137 10965 9171 10999
rect 5181 10761 5215 10795
rect 10241 10761 10275 10795
rect 12449 10761 12483 10795
rect 20821 10761 20855 10795
rect 15577 10693 15611 10727
rect 2329 10625 2363 10659
rect 3893 10625 3927 10659
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 7757 10625 7791 10659
rect 7941 10625 7975 10659
rect 13001 10625 13035 10659
rect 14473 10625 14507 10659
rect 14657 10625 14691 10659
rect 16129 10625 16163 10659
rect 2053 10557 2087 10591
rect 3617 10557 3651 10591
rect 5089 10557 5123 10591
rect 7665 10557 7699 10591
rect 8861 10557 8895 10591
rect 11069 10557 11103 10591
rect 17325 10557 17359 10591
rect 18061 10557 18095 10591
rect 19441 10557 19475 10591
rect 2145 10489 2179 10523
rect 9106 10489 9140 10523
rect 11345 10489 11379 10523
rect 14381 10489 14415 10523
rect 16037 10489 16071 10523
rect 18337 10489 18371 10523
rect 19708 10489 19742 10523
rect 1685 10421 1719 10455
rect 3249 10421 3283 10455
rect 3709 10421 3743 10455
rect 4905 10421 4939 10455
rect 5549 10421 5583 10455
rect 7297 10421 7331 10455
rect 12817 10421 12851 10455
rect 12909 10421 12943 10455
rect 14013 10421 14047 10455
rect 15945 10421 15979 10455
rect 17141 10421 17175 10455
rect 2605 10217 2639 10251
rect 8493 10217 8527 10251
rect 12357 10217 12391 10251
rect 14197 10217 14231 10251
rect 17509 10217 17543 10251
rect 7380 10149 7414 10183
rect 13001 10149 13035 10183
rect 16396 10149 16430 10183
rect 18858 10149 18892 10183
rect 2697 10081 2731 10115
rect 4813 10081 4847 10115
rect 5080 10081 5114 10115
rect 7113 10081 7147 10115
rect 10793 10081 10827 10115
rect 12541 10081 12575 10115
rect 13093 10081 13127 10115
rect 18613 10081 18647 10115
rect 2881 10013 2915 10047
rect 10885 10013 10919 10047
rect 10977 10013 11011 10047
rect 13185 10013 13219 10047
rect 16129 10013 16163 10047
rect 2237 9877 2271 9911
rect 6193 9877 6227 9911
rect 10425 9877 10459 9911
rect 12633 9877 12667 9911
rect 19993 9877 20027 9911
rect 3709 9673 3743 9707
rect 9137 9673 9171 9707
rect 2881 9605 2915 9639
rect 10609 9605 10643 9639
rect 15301 9605 15335 9639
rect 19441 9605 19475 9639
rect 4261 9537 4295 9571
rect 11069 9537 11103 9571
rect 11161 9537 11195 9571
rect 16589 9537 16623 9571
rect 16681 9537 16715 9571
rect 18061 9537 18095 9571
rect 1501 9469 1535 9503
rect 4077 9469 4111 9503
rect 5273 9469 5307 9503
rect 7757 9469 7791 9503
rect 8024 9469 8058 9503
rect 12633 9469 12667 9503
rect 13921 9469 13955 9503
rect 16497 9469 16531 9503
rect 20269 9469 20303 9503
rect 1768 9401 1802 9435
rect 5549 9401 5583 9435
rect 12909 9401 12943 9435
rect 14188 9401 14222 9435
rect 18306 9401 18340 9435
rect 20545 9401 20579 9435
rect 4169 9333 4203 9367
rect 10977 9333 11011 9367
rect 16129 9333 16163 9367
rect 3157 9129 3191 9163
rect 4261 9129 4295 9163
rect 6561 9129 6595 9163
rect 8033 9129 8067 9163
rect 11069 9129 11103 9163
rect 11897 9129 11931 9163
rect 12265 9129 12299 9163
rect 13461 9129 13495 9163
rect 15485 9129 15519 9163
rect 19257 9129 19291 9163
rect 19625 9129 19659 9163
rect 5448 9061 5482 9095
rect 12357 9061 12391 9095
rect 13829 9061 13863 9095
rect 2044 8993 2078 9027
rect 4077 8993 4111 9027
rect 7941 8993 7975 9027
rect 8401 8993 8435 9027
rect 9689 8993 9723 9027
rect 9956 8993 9990 9027
rect 13921 8993 13955 9027
rect 15301 8993 15335 9027
rect 16764 8993 16798 9027
rect 1777 8925 1811 8959
rect 5181 8925 5215 8959
rect 8493 8925 8527 8959
rect 8677 8925 8711 8959
rect 12449 8925 12483 8959
rect 14013 8925 14047 8959
rect 16497 8925 16531 8959
rect 19717 8925 19751 8959
rect 19901 8925 19935 8959
rect 7757 8789 7791 8823
rect 17877 8789 17911 8823
rect 4537 8585 4571 8619
rect 6837 8585 6871 8619
rect 10793 8585 10827 8619
rect 16037 8585 16071 8619
rect 18245 8585 18279 8619
rect 15209 8517 15243 8551
rect 2053 8449 2087 8483
rect 3157 8449 3191 8483
rect 5641 8449 5675 8483
rect 7389 8449 7423 8483
rect 8401 8449 8435 8483
rect 12725 8449 12759 8483
rect 16497 8449 16531 8483
rect 16589 8449 16623 8483
rect 19165 8449 19199 8483
rect 1777 8381 1811 8415
rect 5365 8381 5399 8415
rect 7205 8381 7239 8415
rect 7297 8381 7331 8415
rect 9413 8381 9447 8415
rect 12265 8381 12299 8415
rect 12449 8381 12483 8415
rect 13829 8381 13863 8415
rect 14096 8381 14130 8415
rect 18061 8381 18095 8415
rect 19432 8381 19466 8415
rect 3402 8313 3436 8347
rect 9658 8313 9692 8347
rect 16405 8313 16439 8347
rect 12081 8245 12115 8279
rect 20545 8245 20579 8279
rect 5457 8041 5491 8075
rect 6561 8041 6595 8075
rect 9873 8041 9907 8075
rect 10793 8041 10827 8075
rect 17509 8041 17543 8075
rect 19257 8041 19291 8075
rect 11161 7973 11195 8007
rect 12624 7973 12658 8007
rect 15568 7973 15602 8007
rect 2145 7905 2179 7939
rect 5365 7905 5399 7939
rect 6929 7905 6963 7939
rect 8309 7905 8343 7939
rect 9689 7905 9723 7939
rect 11253 7905 11287 7939
rect 15301 7905 15335 7939
rect 17877 7905 17911 7939
rect 19165 7905 19199 7939
rect 19625 7905 19659 7939
rect 2329 7837 2363 7871
rect 5641 7837 5675 7871
rect 7021 7837 7055 7871
rect 7113 7837 7147 7871
rect 8585 7837 8619 7871
rect 11345 7837 11379 7871
rect 12357 7837 12391 7871
rect 17969 7837 18003 7871
rect 18061 7837 18095 7871
rect 19717 7837 19751 7871
rect 19901 7837 19935 7871
rect 13737 7769 13771 7803
rect 4997 7701 5031 7735
rect 16681 7701 16715 7735
rect 3065 7497 3099 7531
rect 4905 7497 4939 7531
rect 6837 7497 6871 7531
rect 9137 7497 9171 7531
rect 14289 7497 14323 7531
rect 16405 7497 16439 7531
rect 20729 7497 20763 7531
rect 3617 7361 3651 7395
rect 5457 7361 5491 7395
rect 7389 7361 7423 7395
rect 9873 7361 9907 7395
rect 11345 7361 11379 7395
rect 13369 7361 13403 7395
rect 14841 7361 14875 7395
rect 16957 7361 16991 7395
rect 19349 7361 19383 7395
rect 1777 7293 1811 7327
rect 7297 7293 7331 7327
rect 9137 7293 9171 7327
rect 9689 7293 9723 7327
rect 13093 7293 13127 7327
rect 14657 7293 14691 7327
rect 16865 7293 16899 7327
rect 18071 7293 18105 7327
rect 19616 7293 19650 7327
rect 2053 7225 2087 7259
rect 3525 7225 3559 7259
rect 11253 7225 11287 7259
rect 16773 7225 16807 7259
rect 18337 7225 18371 7259
rect 3433 7157 3467 7191
rect 5273 7157 5307 7191
rect 5365 7157 5399 7191
rect 7205 7157 7239 7191
rect 9229 7157 9263 7191
rect 9597 7157 9631 7191
rect 10793 7157 10827 7191
rect 11161 7157 11195 7191
rect 12725 7157 12759 7191
rect 13185 7157 13219 7191
rect 14749 7157 14783 7191
rect 4721 6953 4755 6987
rect 7021 6953 7055 6987
rect 7389 6953 7423 6987
rect 11069 6953 11103 6987
rect 18797 6953 18831 6987
rect 5089 6885 5123 6919
rect 16466 6885 16500 6919
rect 2237 6817 2271 6851
rect 7481 6817 7515 6851
rect 9956 6817 9990 6851
rect 12817 6817 12851 6851
rect 13073 6817 13107 6851
rect 16221 6817 16255 6851
rect 2513 6749 2547 6783
rect 5181 6749 5215 6783
rect 5365 6749 5399 6783
rect 7573 6749 7607 6783
rect 8585 6749 8619 6783
rect 9689 6749 9723 6783
rect 18889 6749 18923 6783
rect 18981 6749 19015 6783
rect 14197 6681 14231 6715
rect 17601 6681 17635 6715
rect 18429 6681 18463 6715
rect 18245 6613 18279 6647
rect 3433 6409 3467 6443
rect 4997 6409 5031 6443
rect 7849 6409 7883 6443
rect 12449 6409 12483 6443
rect 14381 6409 14415 6443
rect 16405 6409 16439 6443
rect 18429 6409 18463 6443
rect 2237 6273 2271 6307
rect 5457 6273 5491 6307
rect 5641 6273 5675 6307
rect 13001 6273 13035 6307
rect 15025 6273 15059 6307
rect 17049 6273 17083 6307
rect 18981 6273 19015 6307
rect 20637 6273 20671 6307
rect 1961 6205 1995 6239
rect 3249 6205 3283 6239
rect 7665 6205 7699 6239
rect 8769 6205 8803 6239
rect 10977 6205 11011 6239
rect 14749 6205 14783 6239
rect 18797 6205 18831 6239
rect 20453 6205 20487 6239
rect 5365 6137 5399 6171
rect 9036 6137 9070 6171
rect 11253 6137 11287 6171
rect 12909 6137 12943 6171
rect 18889 6137 18923 6171
rect 10149 6069 10183 6103
rect 12817 6069 12851 6103
rect 14841 6069 14875 6103
rect 16773 6069 16807 6103
rect 16865 6069 16899 6103
rect 20085 6069 20119 6103
rect 20545 6069 20579 6103
rect 1961 5865 1995 5899
rect 3065 5865 3099 5899
rect 4261 5865 4295 5899
rect 5365 5865 5399 5899
rect 6469 5865 6503 5899
rect 9689 5865 9723 5899
rect 9781 5865 9815 5899
rect 12725 5865 12759 5899
rect 13553 5865 13587 5899
rect 14013 5865 14047 5899
rect 14105 5865 14139 5899
rect 15301 5865 15335 5899
rect 17509 5865 17543 5899
rect 17969 5865 18003 5899
rect 19073 5865 19107 5899
rect 19441 5865 19475 5899
rect 11590 5797 11624 5831
rect 19533 5797 19567 5831
rect 1777 5729 1811 5763
rect 2881 5729 2915 5763
rect 4077 5729 4111 5763
rect 5181 5729 5215 5763
rect 6285 5729 6319 5763
rect 7395 5729 7429 5763
rect 8493 5729 8527 5763
rect 9689 5729 9723 5763
rect 10149 5729 10183 5763
rect 15669 5729 15703 5763
rect 15761 5729 15795 5763
rect 17877 5729 17911 5763
rect 10241 5661 10275 5695
rect 10425 5661 10459 5695
rect 11345 5661 11379 5695
rect 14289 5661 14323 5695
rect 15853 5661 15887 5695
rect 18061 5661 18095 5695
rect 19625 5661 19659 5695
rect 7573 5593 7607 5627
rect 13645 5593 13679 5627
rect 8677 5525 8711 5559
rect 1961 5321 1995 5355
rect 3065 5321 3099 5355
rect 4169 5321 4203 5355
rect 5273 5321 5307 5355
rect 7113 5321 7147 5355
rect 8217 5321 8251 5355
rect 9137 5321 9171 5355
rect 10793 5321 10827 5355
rect 12449 5321 12483 5355
rect 14013 5321 14047 5355
rect 16405 5321 16439 5355
rect 18061 5321 18095 5355
rect 19993 5321 20027 5355
rect 9689 5185 9723 5219
rect 11253 5185 11287 5219
rect 11345 5185 11379 5219
rect 13001 5185 13035 5219
rect 14565 5185 14599 5219
rect 17049 5185 17083 5219
rect 18613 5185 18647 5219
rect 20453 5185 20487 5219
rect 20545 5185 20579 5219
rect 1783 5117 1817 5151
rect 2881 5117 2915 5151
rect 3985 5117 4019 5151
rect 5089 5117 5123 5151
rect 6929 5117 6963 5151
rect 8033 5117 8067 5151
rect 9597 5117 9631 5151
rect 12909 5117 12943 5151
rect 14473 5117 14507 5151
rect 16773 5117 16807 5151
rect 20361 5117 20395 5151
rect 9505 5049 9539 5083
rect 18429 5049 18463 5083
rect 11161 4981 11195 5015
rect 12817 4981 12851 5015
rect 14381 4981 14415 5015
rect 16865 4981 16899 5015
rect 18521 4981 18555 5015
rect 1961 4777 1995 4811
rect 4261 4777 4295 4811
rect 6377 4777 6411 4811
rect 7573 4777 7607 4811
rect 8677 4777 8711 4811
rect 10149 4777 10183 4811
rect 11069 4777 11103 4811
rect 11529 4777 11563 4811
rect 12633 4777 12667 4811
rect 13645 4777 13679 4811
rect 14013 4777 14047 4811
rect 15485 4777 15519 4811
rect 16497 4777 16531 4811
rect 18521 4777 18555 4811
rect 19901 4777 19935 4811
rect 14105 4709 14139 4743
rect 16957 4709 16991 4743
rect 1777 4641 1811 4675
rect 2881 4641 2915 4675
rect 4077 4641 4111 4675
rect 5181 4641 5215 4675
rect 7389 4641 7423 4675
rect 8493 4641 8527 4675
rect 9965 4641 9999 4675
rect 11437 4641 11471 4675
rect 15301 4641 15335 4675
rect 16865 4641 16899 4675
rect 18613 4641 18647 4675
rect 19717 4641 19751 4675
rect 11713 4573 11747 4607
rect 14289 4573 14323 4607
rect 17141 4573 17175 4607
rect 18705 4573 18739 4607
rect 3065 4505 3099 4539
rect 5365 4505 5399 4539
rect 18153 4437 18187 4471
rect 10333 4233 10367 4267
rect 5089 4097 5123 4131
rect 6929 4097 6963 4131
rect 13001 4097 13035 4131
rect 13185 4097 13219 4131
rect 14657 4097 14691 4131
rect 16681 4097 16715 4131
rect 18521 4097 18555 4131
rect 18613 4097 18647 4131
rect 20085 4097 20119 4131
rect 20269 4097 20303 4131
rect 1783 4029 1817 4063
rect 2881 4029 2915 4063
rect 3985 4029 4019 4063
rect 7941 4029 7975 4063
rect 9045 4029 9079 4063
rect 10149 4029 10183 4063
rect 11241 4029 11275 4063
rect 14473 4029 14507 4063
rect 17601 4029 17635 4063
rect 18429 4029 18463 4063
rect 18889 4029 18923 4063
rect 16497 3961 16531 3995
rect 19993 3961 20027 3995
rect 1961 3893 1995 3927
rect 3065 3893 3099 3927
rect 4169 3893 4203 3927
rect 8125 3893 8159 3927
rect 9229 3893 9263 3927
rect 11437 3893 11471 3927
rect 12541 3893 12575 3927
rect 12909 3893 12943 3927
rect 14105 3893 14139 3927
rect 14565 3893 14599 3927
rect 16129 3893 16163 3927
rect 16589 3893 16623 3927
rect 18061 3893 18095 3927
rect 19625 3893 19659 3927
rect 2053 3689 2087 3723
rect 2973 3689 3007 3723
rect 10057 3689 10091 3723
rect 11161 3689 11195 3723
rect 12081 3689 12115 3723
rect 12449 3689 12483 3723
rect 13645 3689 13679 3723
rect 14013 3689 14047 3723
rect 16405 3689 16439 3723
rect 18061 3689 18095 3723
rect 19625 3689 19659 3723
rect 8585 3621 8619 3655
rect 12541 3621 12575 3655
rect 14105 3621 14139 3655
rect 19533 3621 19567 3655
rect 1869 3553 1903 3587
rect 4077 3553 4111 3587
rect 6561 3553 6595 3587
rect 9597 3553 9631 3587
rect 9873 3553 9907 3587
rect 10977 3553 11011 3587
rect 17969 3553 18003 3587
rect 7573 3485 7607 3519
rect 9781 3485 9815 3519
rect 12725 3485 12759 3519
rect 14197 3485 14231 3519
rect 16497 3485 16531 3519
rect 16589 3485 16623 3519
rect 18153 3485 18187 3519
rect 19809 3485 19843 3519
rect 4261 3417 4295 3451
rect 16037 3417 16071 3451
rect 17601 3417 17635 3451
rect 19165 3349 19199 3383
rect 1961 3145 1995 3179
rect 5917 3145 5951 3179
rect 10333 3145 10367 3179
rect 11437 3145 11471 3179
rect 16405 3145 16439 3179
rect 8585 3077 8619 3111
rect 18061 3077 18095 3111
rect 13001 3009 13035 3043
rect 14565 3009 14599 3043
rect 14657 3009 14691 3043
rect 17049 3009 17083 3043
rect 18613 3009 18647 3043
rect 1777 2941 1811 2975
rect 2881 2941 2915 2975
rect 7205 2941 7239 2975
rect 10149 2941 10183 2975
rect 11253 2941 11287 2975
rect 12817 2941 12851 2975
rect 14473 2941 14507 2975
rect 16773 2941 16807 2975
rect 18521 2941 18555 2975
rect 19625 2941 19659 2975
rect 7450 2873 7484 2907
rect 16865 2873 16899 2907
rect 18429 2873 18463 2907
rect 3065 2805 3099 2839
rect 14105 2805 14139 2839
rect 19809 2805 19843 2839
rect 8677 2601 8711 2635
rect 10425 2601 10459 2635
rect 11621 2601 11655 2635
rect 13829 2601 13863 2635
rect 14197 2601 14231 2635
rect 16497 2601 16531 2635
rect 16957 2601 16991 2635
rect 19625 2601 19659 2635
rect 15485 2533 15519 2567
rect 1869 2465 1903 2499
rect 11437 2465 11471 2499
rect 12633 2465 12667 2499
rect 12725 2465 12759 2499
rect 16865 2465 16899 2499
rect 18337 2465 18371 2499
rect 19441 2465 19475 2499
rect 7849 2329 7883 2363
rect 14289 2397 14323 2431
rect 14473 2397 14507 2431
rect 17141 2397 17175 2431
rect 18521 2329 18555 2363
rect 2053 2261 2087 2295
rect 12633 2261 12667 2295
rect 12909 2261 12943 2295
rect 13737 2057 13771 2091
rect 13737 1649 13771 1683
<< metal1 >>
rect 3510 21632 3516 21684
rect 3568 21672 3574 21684
rect 5166 21672 5172 21684
rect 3568 21644 5172 21672
rect 3568 21632 3574 21644
rect 5166 21632 5172 21644
rect 5224 21632 5230 21684
rect 15194 21156 15200 21208
rect 15252 21196 15258 21208
rect 17954 21196 17960 21208
rect 15252 21168 17960 21196
rect 15252 21156 15258 21168
rect 17954 21156 17960 21168
rect 18012 21156 18018 21208
rect 17954 20952 17960 21004
rect 18012 20992 18018 21004
rect 18230 20992 18236 21004
rect 18012 20964 18236 20992
rect 18012 20952 18018 20964
rect 18230 20952 18236 20964
rect 18288 20952 18294 21004
rect 4798 20884 4804 20936
rect 4856 20924 4862 20936
rect 5350 20924 5356 20936
rect 4856 20896 5356 20924
rect 4856 20884 4862 20896
rect 5350 20884 5356 20896
rect 5408 20884 5414 20936
rect 3694 20816 3700 20868
rect 3752 20856 3758 20868
rect 6270 20856 6276 20868
rect 3752 20828 6276 20856
rect 3752 20816 3758 20828
rect 6270 20816 6276 20828
rect 6328 20816 6334 20868
rect 3510 20748 3516 20800
rect 3568 20788 3574 20800
rect 4890 20788 4896 20800
rect 3568 20760 4896 20788
rect 3568 20748 3574 20760
rect 4890 20748 4896 20760
rect 4948 20748 4954 20800
rect 8662 20748 8668 20800
rect 8720 20788 8726 20800
rect 18046 20788 18052 20800
rect 8720 20760 18052 20788
rect 8720 20748 8726 20760
rect 18046 20748 18052 20760
rect 18104 20748 18110 20800
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 5258 20544 5264 20596
rect 5316 20584 5322 20596
rect 8754 20584 8760 20596
rect 5316 20556 8760 20584
rect 5316 20544 5322 20556
rect 8754 20544 8760 20556
rect 8812 20544 8818 20596
rect 9306 20544 9312 20596
rect 9364 20584 9370 20596
rect 13906 20584 13912 20596
rect 9364 20556 13912 20584
rect 9364 20544 9370 20556
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 14461 20587 14519 20593
rect 14461 20553 14473 20587
rect 14507 20584 14519 20587
rect 15194 20584 15200 20596
rect 14507 20556 15200 20584
rect 14507 20553 14519 20556
rect 14461 20547 14519 20553
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 15749 20587 15807 20593
rect 15749 20553 15761 20587
rect 15795 20584 15807 20587
rect 17862 20584 17868 20596
rect 15795 20556 17868 20584
rect 15795 20553 15807 20556
rect 15749 20547 15807 20553
rect 17862 20544 17868 20556
rect 17920 20544 17926 20596
rect 7193 20519 7251 20525
rect 1412 20488 7144 20516
rect 1412 20457 1440 20488
rect 1397 20451 1455 20457
rect 1397 20417 1409 20451
rect 1443 20417 1455 20451
rect 1397 20411 1455 20417
rect 2682 20408 2688 20460
rect 2740 20448 2746 20460
rect 2961 20451 3019 20457
rect 2961 20448 2973 20451
rect 2740 20420 2973 20448
rect 2740 20408 2746 20420
rect 2961 20417 2973 20420
rect 3007 20417 3019 20451
rect 2961 20411 3019 20417
rect 3050 20408 3056 20460
rect 3108 20448 3114 20460
rect 5629 20451 5687 20457
rect 5629 20448 5641 20451
rect 3108 20420 5641 20448
rect 3108 20408 3114 20420
rect 5629 20417 5641 20420
rect 5675 20417 5687 20451
rect 5629 20411 5687 20417
rect 2869 20383 2927 20389
rect 2869 20349 2881 20383
rect 2915 20380 2927 20383
rect 6822 20380 6828 20392
rect 2915 20352 6828 20380
rect 2915 20349 2927 20352
rect 2869 20343 2927 20349
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 6917 20383 6975 20389
rect 6917 20349 6929 20383
rect 6963 20380 6975 20383
rect 7015 20383 7073 20389
rect 7015 20380 7027 20383
rect 6963 20352 7027 20380
rect 6963 20349 6975 20352
rect 6917 20343 6975 20349
rect 7015 20349 7027 20352
rect 7061 20349 7073 20383
rect 7116 20380 7144 20488
rect 7193 20485 7205 20519
rect 7239 20516 7251 20519
rect 18690 20516 18696 20528
rect 7239 20488 18696 20516
rect 7239 20485 7251 20488
rect 7193 20479 7251 20485
rect 18690 20476 18696 20488
rect 18748 20476 18754 20528
rect 7282 20408 7288 20460
rect 7340 20448 7346 20460
rect 8665 20451 8723 20457
rect 8665 20448 8677 20451
rect 7340 20420 8677 20448
rect 7340 20408 7346 20420
rect 8665 20417 8677 20420
rect 8711 20417 8723 20451
rect 8665 20411 8723 20417
rect 11054 20408 11060 20460
rect 11112 20448 11118 20460
rect 11241 20451 11299 20457
rect 11241 20448 11253 20451
rect 11112 20420 11253 20448
rect 11112 20408 11118 20420
rect 11241 20417 11253 20420
rect 11287 20417 11299 20451
rect 13262 20448 13268 20460
rect 13223 20420 13268 20448
rect 11241 20411 11299 20417
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 13354 20408 13360 20460
rect 13412 20448 13418 20460
rect 17126 20448 17132 20460
rect 13412 20420 15700 20448
rect 17087 20420 17132 20448
rect 13412 20408 13418 20420
rect 9030 20380 9036 20392
rect 7116 20352 9036 20380
rect 7015 20343 7073 20349
rect 9030 20340 9036 20352
rect 9088 20340 9094 20392
rect 12158 20380 12164 20392
rect 10060 20352 12164 20380
rect 3970 20272 3976 20324
rect 4028 20312 4034 20324
rect 4982 20312 4988 20324
rect 4028 20284 4988 20312
rect 4028 20272 4034 20284
rect 4982 20272 4988 20284
rect 5040 20272 5046 20324
rect 5537 20315 5595 20321
rect 5537 20281 5549 20315
rect 5583 20312 5595 20315
rect 10060 20312 10088 20352
rect 12158 20340 12164 20352
rect 12216 20380 12222 20392
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 12216 20352 13093 20380
rect 12216 20340 12222 20352
rect 13081 20349 13093 20352
rect 13127 20349 13139 20383
rect 13081 20343 13139 20349
rect 14277 20383 14335 20389
rect 14277 20349 14289 20383
rect 14323 20380 14335 20383
rect 14366 20380 14372 20392
rect 14323 20352 14372 20380
rect 14323 20349 14335 20352
rect 14277 20343 14335 20349
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 15194 20340 15200 20392
rect 15252 20380 15258 20392
rect 15565 20383 15623 20389
rect 15565 20380 15577 20383
rect 15252 20352 15577 20380
rect 15252 20340 15258 20352
rect 15565 20349 15577 20352
rect 15611 20349 15623 20383
rect 15672 20380 15700 20420
rect 17126 20408 17132 20420
rect 17184 20408 17190 20460
rect 17310 20448 17316 20460
rect 17271 20420 17316 20448
rect 17310 20408 17316 20420
rect 17368 20408 17374 20460
rect 19613 20451 19671 20457
rect 19613 20417 19625 20451
rect 19659 20448 19671 20451
rect 19886 20448 19892 20460
rect 19659 20420 19892 20448
rect 19659 20417 19671 20420
rect 19613 20411 19671 20417
rect 19886 20408 19892 20420
rect 19944 20408 19950 20460
rect 19429 20383 19487 20389
rect 19429 20380 19441 20383
rect 15672 20352 19441 20380
rect 15565 20343 15623 20349
rect 19429 20349 19441 20352
rect 19475 20349 19487 20383
rect 19429 20343 19487 20349
rect 5583 20284 10088 20312
rect 5583 20281 5595 20284
rect 5537 20275 5595 20281
rect 10410 20272 10416 20324
rect 10468 20312 10474 20324
rect 11149 20315 11207 20321
rect 11149 20312 11161 20315
rect 10468 20284 11161 20312
rect 10468 20272 10474 20284
rect 11149 20281 11161 20284
rect 11195 20281 11207 20315
rect 17034 20312 17040 20324
rect 16995 20284 17040 20312
rect 11149 20275 11207 20281
rect 17034 20272 17040 20284
rect 17092 20272 17098 20324
rect 2222 20204 2228 20256
rect 2280 20244 2286 20256
rect 2409 20247 2467 20253
rect 2409 20244 2421 20247
rect 2280 20216 2421 20244
rect 2280 20204 2286 20216
rect 2409 20213 2421 20216
rect 2455 20213 2467 20247
rect 2409 20207 2467 20213
rect 2774 20204 2780 20256
rect 2832 20244 2838 20256
rect 2832 20216 2877 20244
rect 2832 20204 2838 20216
rect 3878 20204 3884 20256
rect 3936 20244 3942 20256
rect 4065 20247 4123 20253
rect 4065 20244 4077 20247
rect 3936 20216 4077 20244
rect 3936 20204 3942 20216
rect 4065 20213 4077 20216
rect 4111 20213 4123 20247
rect 4065 20207 4123 20213
rect 4706 20204 4712 20256
rect 4764 20244 4770 20256
rect 5077 20247 5135 20253
rect 5077 20244 5089 20247
rect 4764 20216 5089 20244
rect 4764 20204 4770 20216
rect 5077 20213 5089 20216
rect 5123 20213 5135 20247
rect 5077 20207 5135 20213
rect 5258 20204 5264 20256
rect 5316 20244 5322 20256
rect 5445 20247 5503 20253
rect 5445 20244 5457 20247
rect 5316 20216 5457 20244
rect 5316 20204 5322 20216
rect 5445 20213 5457 20216
rect 5491 20213 5503 20247
rect 5445 20207 5503 20213
rect 6917 20247 6975 20253
rect 6917 20213 6929 20247
rect 6963 20244 6975 20247
rect 7650 20244 7656 20256
rect 6963 20216 7656 20244
rect 6963 20213 6975 20216
rect 6917 20207 6975 20213
rect 7650 20204 7656 20216
rect 7708 20204 7714 20256
rect 8113 20247 8171 20253
rect 8113 20213 8125 20247
rect 8159 20244 8171 20247
rect 8202 20244 8208 20256
rect 8159 20216 8208 20244
rect 8159 20213 8171 20216
rect 8113 20207 8171 20213
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 8478 20244 8484 20256
rect 8439 20216 8484 20244
rect 8478 20204 8484 20216
rect 8536 20204 8542 20256
rect 8573 20247 8631 20253
rect 8573 20213 8585 20247
rect 8619 20244 8631 20247
rect 8754 20244 8760 20256
rect 8619 20216 8760 20244
rect 8619 20213 8631 20216
rect 8573 20207 8631 20213
rect 8754 20204 8760 20216
rect 8812 20204 8818 20256
rect 10686 20244 10692 20256
rect 10647 20216 10692 20244
rect 10686 20204 10692 20216
rect 10744 20204 10750 20256
rect 10962 20204 10968 20256
rect 11020 20244 11026 20256
rect 11057 20247 11115 20253
rect 11057 20244 11069 20247
rect 11020 20216 11069 20244
rect 11020 20204 11026 20216
rect 11057 20213 11069 20216
rect 11103 20213 11115 20247
rect 11057 20207 11115 20213
rect 12342 20204 12348 20256
rect 12400 20244 12406 20256
rect 12621 20247 12679 20253
rect 12621 20244 12633 20247
rect 12400 20216 12633 20244
rect 12400 20204 12406 20216
rect 12621 20213 12633 20216
rect 12667 20213 12679 20247
rect 12621 20207 12679 20213
rect 12989 20247 13047 20253
rect 12989 20213 13001 20247
rect 13035 20244 13047 20247
rect 13170 20244 13176 20256
rect 13035 20216 13176 20244
rect 13035 20213 13047 20216
rect 12989 20207 13047 20213
rect 13170 20204 13176 20216
rect 13228 20204 13234 20256
rect 16666 20244 16672 20256
rect 16627 20216 16672 20244
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 18966 20244 18972 20256
rect 18927 20216 18972 20244
rect 18966 20204 18972 20216
rect 19024 20204 19030 20256
rect 19058 20204 19064 20256
rect 19116 20244 19122 20256
rect 19337 20247 19395 20253
rect 19337 20244 19349 20247
rect 19116 20216 19349 20244
rect 19116 20204 19122 20216
rect 19337 20213 19349 20216
rect 19383 20213 19395 20247
rect 19337 20207 19395 20213
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4341 20043 4399 20049
rect 4341 20040 4353 20043
rect 4212 20012 4353 20040
rect 4212 20000 4218 20012
rect 4341 20009 4353 20012
rect 4387 20009 4399 20043
rect 4341 20003 4399 20009
rect 4706 20000 4712 20052
rect 4764 20040 4770 20052
rect 4764 20012 4809 20040
rect 4764 20000 4770 20012
rect 5442 20000 5448 20052
rect 5500 20040 5506 20052
rect 6273 20043 6331 20049
rect 6273 20040 6285 20043
rect 5500 20012 6285 20040
rect 5500 20000 5506 20012
rect 6273 20009 6285 20012
rect 6319 20009 6331 20043
rect 6273 20003 6331 20009
rect 8021 20043 8079 20049
rect 8021 20009 8033 20043
rect 8067 20040 8079 20043
rect 10410 20040 10416 20052
rect 8067 20012 10416 20040
rect 8067 20009 8079 20012
rect 8021 20003 8079 20009
rect 10410 20000 10416 20012
rect 10468 20000 10474 20052
rect 12253 20043 12311 20049
rect 12253 20009 12265 20043
rect 12299 20040 12311 20043
rect 13449 20043 13507 20049
rect 13449 20040 13461 20043
rect 12299 20012 13461 20040
rect 12299 20009 12311 20012
rect 12253 20003 12311 20009
rect 13449 20009 13461 20012
rect 13495 20009 13507 20043
rect 13449 20003 13507 20009
rect 16666 20000 16672 20052
rect 16724 20040 16730 20052
rect 17037 20043 17095 20049
rect 17037 20040 17049 20043
rect 16724 20012 17049 20040
rect 16724 20000 16730 20012
rect 17037 20009 17049 20012
rect 17083 20009 17095 20043
rect 17037 20003 17095 20009
rect 2777 19975 2835 19981
rect 2777 19941 2789 19975
rect 2823 19972 2835 19975
rect 8389 19975 8447 19981
rect 8389 19972 8401 19975
rect 2823 19944 8401 19972
rect 2823 19941 2835 19944
rect 2777 19935 2835 19941
rect 8389 19941 8401 19944
rect 8435 19972 8447 19975
rect 8938 19972 8944 19984
rect 8435 19944 8944 19972
rect 8435 19941 8447 19944
rect 8389 19935 8447 19941
rect 8938 19932 8944 19944
rect 8996 19932 9002 19984
rect 9030 19932 9036 19984
rect 9088 19972 9094 19984
rect 12345 19975 12403 19981
rect 9088 19944 10824 19972
rect 9088 19932 9094 19944
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19904 2927 19907
rect 5718 19904 5724 19916
rect 2915 19876 5724 19904
rect 2915 19873 2927 19876
rect 2869 19867 2927 19873
rect 5718 19864 5724 19876
rect 5776 19904 5782 19916
rect 5776 19876 6500 19904
rect 5776 19864 5782 19876
rect 1397 19839 1455 19845
rect 1397 19805 1409 19839
rect 1443 19836 1455 19839
rect 1854 19836 1860 19848
rect 1443 19808 1860 19836
rect 1443 19805 1455 19808
rect 1397 19799 1455 19805
rect 1854 19796 1860 19808
rect 1912 19796 1918 19848
rect 3050 19836 3056 19848
rect 3011 19808 3056 19836
rect 3050 19796 3056 19808
rect 3108 19796 3114 19848
rect 4801 19839 4859 19845
rect 4801 19805 4813 19839
rect 4847 19805 4859 19839
rect 4801 19799 4859 19805
rect 2409 19771 2467 19777
rect 2409 19737 2421 19771
rect 2455 19768 2467 19771
rect 4816 19768 4844 19799
rect 4890 19796 4896 19848
rect 4948 19836 4954 19848
rect 6362 19836 6368 19848
rect 4948 19808 4993 19836
rect 6323 19808 6368 19836
rect 4948 19796 4954 19808
rect 6362 19796 6368 19808
rect 6420 19796 6426 19848
rect 2455 19740 4844 19768
rect 6472 19768 6500 19876
rect 6822 19864 6828 19916
rect 6880 19904 6886 19916
rect 9944 19907 10002 19913
rect 9944 19904 9956 19907
rect 6880 19876 8616 19904
rect 6880 19864 6886 19876
rect 6549 19839 6607 19845
rect 6549 19805 6561 19839
rect 6595 19836 6607 19839
rect 7282 19836 7288 19848
rect 6595 19808 7288 19836
rect 6595 19805 6607 19808
rect 6549 19799 6607 19805
rect 7282 19796 7288 19808
rect 7340 19796 7346 19848
rect 8481 19839 8539 19845
rect 8481 19805 8493 19839
rect 8527 19805 8539 19839
rect 8481 19799 8539 19805
rect 8496 19768 8524 19799
rect 6472 19740 8524 19768
rect 2455 19737 2467 19740
rect 2409 19731 2467 19737
rect 2866 19660 2872 19712
rect 2924 19700 2930 19712
rect 5442 19700 5448 19712
rect 2924 19672 5448 19700
rect 2924 19660 2930 19672
rect 5442 19660 5448 19672
rect 5500 19660 5506 19712
rect 5905 19703 5963 19709
rect 5905 19669 5917 19703
rect 5951 19700 5963 19703
rect 7282 19700 7288 19712
rect 5951 19672 7288 19700
rect 5951 19669 5963 19672
rect 5905 19663 5963 19669
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 8588 19700 8616 19876
rect 8680 19876 9956 19904
rect 8680 19845 8708 19876
rect 9944 19873 9956 19876
rect 9990 19904 10002 19907
rect 10796 19904 10824 19944
rect 12345 19941 12357 19975
rect 12391 19972 12403 19975
rect 12434 19972 12440 19984
rect 12391 19944 12440 19972
rect 12391 19941 12403 19944
rect 12345 19935 12403 19941
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 13906 19932 13912 19984
rect 13964 19972 13970 19984
rect 15565 19975 15623 19981
rect 15565 19972 15577 19975
rect 13964 19944 15577 19972
rect 13964 19932 13970 19944
rect 15565 19941 15577 19944
rect 15611 19941 15623 19975
rect 15565 19935 15623 19941
rect 13817 19907 13875 19913
rect 13817 19904 13829 19907
rect 9990 19876 10732 19904
rect 10796 19876 13829 19904
rect 9990 19873 10002 19876
rect 9944 19867 10002 19873
rect 8665 19839 8723 19845
rect 8665 19805 8677 19839
rect 8711 19805 8723 19839
rect 8665 19799 8723 19805
rect 9490 19796 9496 19848
rect 9548 19836 9554 19848
rect 9677 19839 9735 19845
rect 9677 19836 9689 19839
rect 9548 19808 9689 19836
rect 9548 19796 9554 19808
rect 9677 19805 9689 19808
rect 9723 19805 9735 19839
rect 9677 19799 9735 19805
rect 10704 19768 10732 19876
rect 13817 19873 13829 19876
rect 13863 19873 13875 19907
rect 14366 19904 14372 19916
rect 13817 19867 13875 19873
rect 13924 19876 14372 19904
rect 11054 19796 11060 19848
rect 11112 19836 11118 19848
rect 13924 19845 13952 19876
rect 14366 19864 14372 19876
rect 14424 19864 14430 19916
rect 15286 19904 15292 19916
rect 15247 19876 15292 19904
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 18233 19907 18291 19913
rect 18233 19873 18245 19907
rect 18279 19904 18291 19907
rect 19613 19907 19671 19913
rect 19613 19904 19625 19907
rect 18279 19876 19625 19904
rect 18279 19873 18291 19876
rect 18233 19867 18291 19873
rect 19613 19873 19625 19876
rect 19659 19873 19671 19907
rect 19613 19867 19671 19873
rect 12437 19839 12495 19845
rect 12437 19836 12449 19839
rect 11112 19808 12449 19836
rect 11112 19796 11118 19808
rect 12437 19805 12449 19808
rect 12483 19805 12495 19839
rect 12437 19799 12495 19805
rect 13909 19839 13967 19845
rect 13909 19805 13921 19839
rect 13955 19805 13967 19839
rect 13909 19799 13967 19805
rect 14001 19839 14059 19845
rect 14001 19805 14013 19839
rect 14047 19805 14059 19839
rect 17126 19836 17132 19848
rect 17087 19808 17132 19836
rect 14001 19799 14059 19805
rect 13262 19768 13268 19780
rect 10704 19740 13268 19768
rect 13262 19728 13268 19740
rect 13320 19768 13326 19780
rect 14016 19768 14044 19799
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 17310 19836 17316 19848
rect 17271 19808 17316 19836
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 19705 19839 19763 19845
rect 19705 19805 19717 19839
rect 19751 19805 19763 19839
rect 19886 19836 19892 19848
rect 19847 19808 19892 19836
rect 19705 19799 19763 19805
rect 13320 19740 14044 19768
rect 13320 19728 13326 19740
rect 14090 19728 14096 19780
rect 14148 19768 14154 19780
rect 19720 19768 19748 19799
rect 19886 19796 19892 19808
rect 19944 19796 19950 19848
rect 14148 19740 19748 19768
rect 14148 19728 14154 19740
rect 10870 19700 10876 19712
rect 8588 19672 10876 19700
rect 10870 19660 10876 19672
rect 10928 19660 10934 19712
rect 11054 19700 11060 19712
rect 11015 19672 11060 19700
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 11882 19700 11888 19712
rect 11843 19672 11888 19700
rect 11882 19660 11888 19672
rect 11940 19660 11946 19712
rect 16669 19703 16727 19709
rect 16669 19669 16681 19703
rect 16715 19700 16727 19703
rect 18046 19700 18052 19712
rect 16715 19672 18052 19700
rect 16715 19669 16727 19672
rect 16669 19663 16727 19669
rect 18046 19660 18052 19672
rect 18104 19660 18110 19712
rect 19242 19700 19248 19712
rect 19203 19672 19248 19700
rect 19242 19660 19248 19672
rect 19300 19660 19306 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 3160 19468 4292 19496
rect 2409 19363 2467 19369
rect 2409 19329 2421 19363
rect 2455 19360 2467 19363
rect 2682 19360 2688 19372
rect 2455 19332 2688 19360
rect 2455 19329 2467 19332
rect 2409 19323 2467 19329
rect 2682 19320 2688 19332
rect 2740 19360 2746 19372
rect 3160 19360 3188 19468
rect 4264 19428 4292 19468
rect 5534 19456 5540 19508
rect 5592 19496 5598 19508
rect 8294 19496 8300 19508
rect 5592 19468 8300 19496
rect 5592 19456 5598 19468
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 16942 19496 16948 19508
rect 16855 19468 16948 19496
rect 16942 19456 16948 19468
rect 17000 19496 17006 19508
rect 17218 19496 17224 19508
rect 17000 19468 17224 19496
rect 17000 19456 17006 19468
rect 17218 19456 17224 19468
rect 17276 19456 17282 19508
rect 4264 19400 7512 19428
rect 3326 19360 3332 19372
rect 2740 19332 3188 19360
rect 3287 19332 3332 19360
rect 2740 19320 2746 19332
rect 3326 19320 3332 19332
rect 3384 19320 3390 19372
rect 7377 19363 7435 19369
rect 7377 19329 7389 19363
rect 7423 19329 7435 19363
rect 7484 19360 7512 19400
rect 7742 19388 7748 19440
rect 7800 19428 7806 19440
rect 8386 19428 8392 19440
rect 7800 19400 8392 19428
rect 7800 19388 7806 19400
rect 8386 19388 8392 19400
rect 8444 19388 8450 19440
rect 8573 19431 8631 19437
rect 8573 19397 8585 19431
rect 8619 19428 8631 19431
rect 8662 19428 8668 19440
rect 8619 19400 8668 19428
rect 8619 19397 8631 19400
rect 8573 19391 8631 19397
rect 8662 19388 8668 19400
rect 8720 19388 8726 19440
rect 17954 19388 17960 19440
rect 18012 19428 18018 19440
rect 18138 19428 18144 19440
rect 18012 19400 18144 19428
rect 18012 19388 18018 19400
rect 18138 19388 18144 19400
rect 18196 19388 18202 19440
rect 7484 19332 9628 19360
rect 7377 19323 7435 19329
rect 5629 19295 5687 19301
rect 5629 19261 5641 19295
rect 5675 19292 5687 19295
rect 6914 19292 6920 19304
rect 5675 19264 6920 19292
rect 5675 19261 5687 19264
rect 5629 19255 5687 19261
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 7282 19292 7288 19304
rect 7243 19264 7288 19292
rect 7282 19252 7288 19264
rect 7340 19252 7346 19304
rect 7392 19292 7420 19323
rect 7650 19292 7656 19304
rect 7392 19264 7656 19292
rect 7650 19252 7656 19264
rect 7708 19252 7714 19304
rect 8202 19252 8208 19304
rect 8260 19252 8266 19304
rect 8389 19295 8447 19301
rect 8389 19261 8401 19295
rect 8435 19292 8447 19295
rect 8570 19292 8576 19304
rect 8435 19264 8576 19292
rect 8435 19261 8447 19264
rect 8389 19255 8447 19261
rect 8570 19252 8576 19264
rect 8628 19252 8634 19304
rect 9490 19292 9496 19304
rect 9451 19264 9496 19292
rect 9490 19252 9496 19264
rect 9548 19252 9554 19304
rect 9600 19292 9628 19332
rect 16666 19320 16672 19372
rect 16724 19360 16730 19372
rect 18690 19360 18696 19372
rect 16724 19332 18696 19360
rect 16724 19320 16730 19332
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 18966 19320 18972 19372
rect 19024 19360 19030 19372
rect 19337 19363 19395 19369
rect 19337 19360 19349 19363
rect 19024 19332 19349 19360
rect 19024 19320 19030 19332
rect 19337 19329 19349 19332
rect 19383 19329 19395 19363
rect 19337 19323 19395 19329
rect 19521 19363 19579 19369
rect 19521 19329 19533 19363
rect 19567 19360 19579 19363
rect 20162 19360 20168 19372
rect 19567 19332 20168 19360
rect 19567 19329 19579 19332
rect 19521 19323 19579 19329
rect 20162 19320 20168 19332
rect 20220 19320 20226 19372
rect 9600 19264 11192 19292
rect 3050 19184 3056 19236
rect 3108 19224 3114 19236
rect 3574 19227 3632 19233
rect 3574 19224 3586 19227
rect 3108 19196 3586 19224
rect 3108 19184 3114 19196
rect 3574 19193 3586 19196
rect 3620 19224 3632 19227
rect 3694 19224 3700 19236
rect 3620 19196 3700 19224
rect 3620 19193 3632 19196
rect 3574 19187 3632 19193
rect 3694 19184 3700 19196
rect 3752 19184 3758 19236
rect 5718 19224 5724 19236
rect 4172 19196 5724 19224
rect 1762 19156 1768 19168
rect 1723 19128 1768 19156
rect 1762 19116 1768 19128
rect 1820 19116 1826 19168
rect 2130 19156 2136 19168
rect 2091 19128 2136 19156
rect 2130 19116 2136 19128
rect 2188 19116 2194 19168
rect 2225 19159 2283 19165
rect 2225 19125 2237 19159
rect 2271 19156 2283 19159
rect 2682 19156 2688 19168
rect 2271 19128 2688 19156
rect 2271 19125 2283 19128
rect 2225 19119 2283 19125
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 3142 19116 3148 19168
rect 3200 19156 3206 19168
rect 4172 19156 4200 19196
rect 5718 19184 5724 19196
rect 5776 19184 5782 19236
rect 8220 19224 8248 19252
rect 8478 19224 8484 19236
rect 8220 19196 8484 19224
rect 8478 19184 8484 19196
rect 8536 19184 8542 19236
rect 9760 19227 9818 19233
rect 9760 19193 9772 19227
rect 9806 19224 9818 19227
rect 11054 19224 11060 19236
rect 9806 19196 11060 19224
rect 9806 19193 9818 19196
rect 9760 19187 9818 19193
rect 11054 19184 11060 19196
rect 11112 19184 11118 19236
rect 11164 19224 11192 19264
rect 11514 19252 11520 19304
rect 11572 19292 11578 19304
rect 13357 19295 13415 19301
rect 13357 19292 13369 19295
rect 11572 19264 13369 19292
rect 11572 19252 11578 19264
rect 13357 19261 13369 19264
rect 13403 19261 13415 19295
rect 13357 19255 13415 19261
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19261 15623 19295
rect 19242 19292 19248 19304
rect 19203 19264 19248 19292
rect 15565 19255 15623 19261
rect 11974 19224 11980 19236
rect 11164 19196 11980 19224
rect 11974 19184 11980 19196
rect 12032 19184 12038 19236
rect 13624 19227 13682 19233
rect 13624 19193 13636 19227
rect 13670 19224 13682 19227
rect 14550 19224 14556 19236
rect 13670 19196 14556 19224
rect 13670 19193 13682 19196
rect 13624 19187 13682 19193
rect 14550 19184 14556 19196
rect 14608 19184 14614 19236
rect 15470 19184 15476 19236
rect 15528 19224 15534 19236
rect 15580 19224 15608 19255
rect 19242 19252 19248 19264
rect 19300 19252 19306 19304
rect 20070 19252 20076 19304
rect 20128 19292 20134 19304
rect 20533 19295 20591 19301
rect 20533 19292 20545 19295
rect 20128 19264 20545 19292
rect 20128 19252 20134 19264
rect 20533 19261 20545 19264
rect 20579 19261 20591 19295
rect 20533 19255 20591 19261
rect 15810 19227 15868 19233
rect 15810 19224 15822 19227
rect 15528 19196 15608 19224
rect 15672 19196 15822 19224
rect 15528 19184 15534 19196
rect 3200 19128 4200 19156
rect 3200 19116 3206 19128
rect 4246 19116 4252 19168
rect 4304 19156 4310 19168
rect 4709 19159 4767 19165
rect 4709 19156 4721 19159
rect 4304 19128 4721 19156
rect 4304 19116 4310 19128
rect 4709 19125 4721 19128
rect 4755 19156 4767 19159
rect 4890 19156 4896 19168
rect 4755 19128 4896 19156
rect 4755 19125 4767 19128
rect 4709 19119 4767 19125
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 5810 19156 5816 19168
rect 5771 19128 5816 19156
rect 5810 19116 5816 19128
rect 5868 19116 5874 19168
rect 6822 19156 6828 19168
rect 6783 19128 6828 19156
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 7190 19156 7196 19168
rect 7151 19128 7196 19156
rect 7190 19116 7196 19128
rect 7248 19116 7254 19168
rect 10778 19116 10784 19168
rect 10836 19156 10842 19168
rect 10873 19159 10931 19165
rect 10873 19156 10885 19159
rect 10836 19128 10885 19156
rect 10836 19116 10842 19128
rect 10873 19125 10885 19128
rect 10919 19125 10931 19159
rect 10873 19119 10931 19125
rect 10962 19116 10968 19168
rect 11020 19156 11026 19168
rect 11698 19156 11704 19168
rect 11020 19128 11704 19156
rect 11020 19116 11026 19128
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 11790 19116 11796 19168
rect 11848 19156 11854 19168
rect 13998 19156 14004 19168
rect 11848 19128 14004 19156
rect 11848 19116 11854 19128
rect 13998 19116 14004 19128
rect 14056 19116 14062 19168
rect 14642 19116 14648 19168
rect 14700 19156 14706 19168
rect 14737 19159 14795 19165
rect 14737 19156 14749 19159
rect 14700 19128 14749 19156
rect 14700 19116 14706 19128
rect 14737 19125 14749 19128
rect 14783 19156 14795 19159
rect 15672 19156 15700 19196
rect 15810 19193 15822 19196
rect 15856 19193 15868 19227
rect 15810 19187 15868 19193
rect 16574 19184 16580 19236
rect 16632 19224 16638 19236
rect 19794 19224 19800 19236
rect 16632 19196 19800 19224
rect 16632 19184 16638 19196
rect 19794 19184 19800 19196
rect 19852 19184 19858 19236
rect 14783 19128 15700 19156
rect 14783 19125 14795 19128
rect 14737 19119 14795 19125
rect 16298 19116 16304 19168
rect 16356 19156 16362 19168
rect 18877 19159 18935 19165
rect 18877 19156 18889 19159
rect 16356 19128 18889 19156
rect 16356 19116 16362 19128
rect 18877 19125 18889 19128
rect 18923 19125 18935 19159
rect 20714 19156 20720 19168
rect 20675 19128 20720 19156
rect 18877 19119 18935 19125
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1394 18952 1400 18964
rect 1355 18924 1400 18952
rect 1394 18912 1400 18924
rect 1452 18912 1458 18964
rect 2777 18955 2835 18961
rect 2777 18921 2789 18955
rect 2823 18952 2835 18955
rect 4062 18952 4068 18964
rect 2823 18924 4068 18952
rect 2823 18921 2835 18924
rect 2777 18915 2835 18921
rect 4062 18912 4068 18924
rect 4120 18912 4126 18964
rect 4154 18912 4160 18964
rect 4212 18952 4218 18964
rect 4525 18955 4583 18961
rect 4525 18952 4537 18955
rect 4212 18924 4537 18952
rect 4212 18912 4218 18924
rect 4525 18921 4537 18924
rect 4571 18921 4583 18955
rect 4525 18915 4583 18921
rect 6733 18955 6791 18961
rect 6733 18921 6745 18955
rect 6779 18952 6791 18955
rect 7837 18955 7895 18961
rect 7837 18952 7849 18955
rect 6779 18924 7849 18952
rect 6779 18921 6791 18924
rect 6733 18915 6791 18921
rect 7837 18921 7849 18924
rect 7883 18921 7895 18955
rect 7837 18915 7895 18921
rect 8202 18912 8208 18964
rect 8260 18952 8266 18964
rect 8297 18955 8355 18961
rect 8297 18952 8309 18955
rect 8260 18924 8309 18952
rect 8260 18912 8266 18924
rect 8297 18921 8309 18924
rect 8343 18921 8355 18955
rect 10410 18952 10416 18964
rect 8297 18915 8355 18921
rect 8404 18924 10416 18952
rect 1578 18844 1584 18896
rect 1636 18884 1642 18896
rect 5810 18884 5816 18896
rect 1636 18856 5816 18884
rect 1636 18844 1642 18856
rect 5810 18844 5816 18856
rect 5868 18844 5874 18896
rect 6641 18887 6699 18893
rect 6641 18853 6653 18887
rect 6687 18884 6699 18887
rect 6822 18884 6828 18896
rect 6687 18856 6828 18884
rect 6687 18853 6699 18856
rect 6641 18847 6699 18853
rect 6822 18844 6828 18856
rect 6880 18844 6886 18896
rect 8404 18884 8432 18924
rect 10410 18912 10416 18924
rect 10468 18912 10474 18964
rect 10686 18952 10692 18964
rect 10647 18924 10692 18952
rect 10686 18912 10692 18924
rect 10744 18912 10750 18964
rect 12526 18912 12532 18964
rect 12584 18952 12590 18964
rect 15194 18952 15200 18964
rect 12584 18924 15200 18952
rect 12584 18912 12590 18924
rect 15194 18912 15200 18924
rect 15252 18912 15258 18964
rect 15289 18955 15347 18961
rect 15289 18921 15301 18955
rect 15335 18952 15347 18955
rect 17034 18952 17040 18964
rect 15335 18924 17040 18952
rect 15335 18921 15347 18924
rect 15289 18915 15347 18921
rect 17034 18912 17040 18924
rect 17092 18912 17098 18964
rect 17310 18912 17316 18964
rect 17368 18952 17374 18964
rect 17681 18955 17739 18961
rect 17681 18952 17693 18955
rect 17368 18924 17693 18952
rect 17368 18912 17374 18924
rect 17681 18921 17693 18924
rect 17727 18921 17739 18955
rect 17681 18915 17739 18921
rect 8128 18856 8432 18884
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18816 2927 18819
rect 2915 18788 4016 18816
rect 2915 18785 2927 18788
rect 2869 18779 2927 18785
rect 3053 18751 3111 18757
rect 3053 18717 3065 18751
rect 3099 18717 3111 18751
rect 3988 18748 4016 18788
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 4212 18788 4445 18816
rect 4212 18776 4218 18788
rect 4433 18785 4445 18788
rect 4479 18785 4491 18819
rect 8128 18816 8156 18856
rect 8754 18844 8760 18896
rect 8812 18884 8818 18896
rect 10597 18887 10655 18893
rect 8812 18856 9812 18884
rect 8812 18844 8818 18856
rect 4433 18779 4491 18785
rect 4632 18788 8156 18816
rect 8205 18819 8263 18825
rect 4632 18748 4660 18788
rect 8205 18785 8217 18819
rect 8251 18816 8263 18819
rect 9674 18816 9680 18828
rect 8251 18788 9680 18816
rect 8251 18785 8263 18788
rect 8205 18779 8263 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 9784 18816 9812 18856
rect 10597 18853 10609 18887
rect 10643 18884 10655 18887
rect 11882 18884 11888 18896
rect 10643 18856 11888 18884
rect 10643 18853 10655 18856
rect 10597 18847 10655 18853
rect 11882 18844 11888 18856
rect 11940 18844 11946 18896
rect 17696 18884 17724 18915
rect 18754 18887 18812 18893
rect 18754 18884 18766 18887
rect 16316 18856 17632 18884
rect 17696 18856 18766 18884
rect 11606 18816 11612 18828
rect 9784 18788 11612 18816
rect 11606 18776 11612 18788
rect 11664 18776 11670 18828
rect 11698 18776 11704 18828
rect 11756 18816 11762 18828
rect 12049 18819 12107 18825
rect 12049 18816 12061 18819
rect 11756 18788 12061 18816
rect 11756 18776 11762 18788
rect 12049 18785 12061 18788
rect 12095 18785 12107 18819
rect 14090 18816 14096 18828
rect 14051 18788 14096 18816
rect 12049 18779 12107 18785
rect 14090 18776 14096 18788
rect 14148 18776 14154 18828
rect 14458 18776 14464 18828
rect 14516 18816 14522 18828
rect 15470 18816 15476 18828
rect 14516 18788 15476 18816
rect 14516 18776 14522 18788
rect 15470 18776 15476 18788
rect 15528 18776 15534 18828
rect 15562 18776 15568 18828
rect 15620 18816 15626 18828
rect 16316 18825 16344 18856
rect 16301 18819 16359 18825
rect 16301 18816 16313 18819
rect 15620 18788 16313 18816
rect 15620 18776 15626 18788
rect 16301 18785 16313 18788
rect 16347 18785 16359 18819
rect 16301 18779 16359 18785
rect 16568 18819 16626 18825
rect 16568 18785 16580 18819
rect 16614 18816 16626 18819
rect 16942 18816 16948 18828
rect 16614 18788 16948 18816
rect 16614 18785 16626 18788
rect 16568 18779 16626 18785
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 17604 18816 17632 18856
rect 18754 18853 18766 18856
rect 18800 18853 18812 18887
rect 18754 18847 18812 18853
rect 17954 18816 17960 18828
rect 17604 18788 17960 18816
rect 17954 18776 17960 18788
rect 18012 18816 18018 18828
rect 18509 18819 18567 18825
rect 18509 18816 18521 18819
rect 18012 18788 18521 18816
rect 18012 18776 18018 18788
rect 18509 18785 18521 18788
rect 18555 18785 18567 18819
rect 18509 18779 18567 18785
rect 3988 18720 4660 18748
rect 4709 18751 4767 18757
rect 3053 18711 3111 18717
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 4798 18748 4804 18760
rect 4755 18720 4804 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 2409 18683 2467 18689
rect 2409 18649 2421 18683
rect 2455 18680 2467 18683
rect 2774 18680 2780 18692
rect 2455 18652 2780 18680
rect 2455 18649 2467 18652
rect 2409 18643 2467 18649
rect 2774 18640 2780 18652
rect 2832 18640 2838 18692
rect 3068 18680 3096 18711
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 4982 18708 4988 18760
rect 5040 18748 5046 18760
rect 5166 18748 5172 18760
rect 5040 18720 5172 18748
rect 5040 18708 5046 18720
rect 5166 18708 5172 18720
rect 5224 18708 5230 18760
rect 6822 18748 6828 18760
rect 6783 18720 6828 18748
rect 6822 18708 6828 18720
rect 6880 18708 6886 18760
rect 7650 18708 7656 18760
rect 7708 18748 7714 18760
rect 8389 18751 8447 18757
rect 8389 18748 8401 18751
rect 7708 18720 8401 18748
rect 7708 18708 7714 18720
rect 8220 18692 8248 18720
rect 8389 18717 8401 18720
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 8662 18708 8668 18760
rect 8720 18748 8726 18760
rect 10594 18748 10600 18760
rect 8720 18720 10600 18748
rect 8720 18708 8726 18720
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 10778 18748 10784 18760
rect 10739 18720 10784 18748
rect 10778 18708 10784 18720
rect 10836 18708 10842 18760
rect 11054 18708 11060 18760
rect 11112 18748 11118 18760
rect 11514 18748 11520 18760
rect 11112 18720 11520 18748
rect 11112 18708 11118 18720
rect 11514 18708 11520 18720
rect 11572 18748 11578 18760
rect 11793 18751 11851 18757
rect 11793 18748 11805 18751
rect 11572 18720 11805 18748
rect 11572 18708 11578 18720
rect 11793 18717 11805 18720
rect 11839 18717 11851 18751
rect 11793 18711 11851 18717
rect 3068 18652 6592 18680
rect 2590 18572 2596 18624
rect 2648 18612 2654 18624
rect 4065 18615 4123 18621
rect 4065 18612 4077 18615
rect 2648 18584 4077 18612
rect 2648 18572 2654 18584
rect 4065 18581 4077 18584
rect 4111 18581 4123 18615
rect 4065 18575 4123 18581
rect 5166 18572 5172 18624
rect 5224 18612 5230 18624
rect 6273 18615 6331 18621
rect 6273 18612 6285 18615
rect 5224 18584 6285 18612
rect 5224 18572 5230 18584
rect 6273 18581 6285 18584
rect 6319 18581 6331 18615
rect 6564 18612 6592 18652
rect 6638 18640 6644 18692
rect 6696 18680 6702 18692
rect 7374 18680 7380 18692
rect 6696 18652 7380 18680
rect 6696 18640 6702 18652
rect 7374 18640 7380 18652
rect 7432 18640 7438 18692
rect 8202 18640 8208 18692
rect 8260 18640 8266 18692
rect 8478 18640 8484 18692
rect 8536 18680 8542 18692
rect 8846 18680 8852 18692
rect 8536 18652 8852 18680
rect 8536 18640 8542 18652
rect 8846 18640 8852 18652
rect 8904 18640 8910 18692
rect 13173 18683 13231 18689
rect 13173 18649 13185 18683
rect 13219 18680 13231 18683
rect 13262 18680 13268 18692
rect 13219 18652 13268 18680
rect 13219 18649 13231 18652
rect 13173 18643 13231 18649
rect 13262 18640 13268 18652
rect 13320 18640 13326 18692
rect 9582 18612 9588 18624
rect 6564 18584 9588 18612
rect 6273 18575 6331 18581
rect 9582 18572 9588 18584
rect 9640 18572 9646 18624
rect 10229 18615 10287 18621
rect 10229 18581 10241 18615
rect 10275 18612 10287 18615
rect 10594 18612 10600 18624
rect 10275 18584 10600 18612
rect 10275 18581 10287 18584
rect 10229 18575 10287 18581
rect 10594 18572 10600 18584
rect 10652 18572 10658 18624
rect 14277 18615 14335 18621
rect 14277 18581 14289 18615
rect 14323 18612 14335 18615
rect 18782 18612 18788 18624
rect 14323 18584 18788 18612
rect 14323 18581 14335 18584
rect 14277 18575 14335 18581
rect 18782 18572 18788 18584
rect 18840 18572 18846 18624
rect 19886 18612 19892 18624
rect 19847 18584 19892 18612
rect 19886 18572 19892 18584
rect 19944 18572 19950 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 4709 18411 4767 18417
rect 2424 18380 4660 18408
rect 2222 18272 2228 18284
rect 2183 18244 2228 18272
rect 2222 18232 2228 18244
rect 2280 18232 2286 18284
rect 2424 18281 2452 18380
rect 4632 18340 4660 18380
rect 4709 18377 4721 18411
rect 4755 18408 4767 18411
rect 4798 18408 4804 18420
rect 4755 18380 4804 18408
rect 4755 18377 4767 18380
rect 4709 18371 4767 18377
rect 4798 18368 4804 18380
rect 4856 18368 4862 18420
rect 11698 18408 11704 18420
rect 6840 18380 11704 18408
rect 6840 18340 6868 18380
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 12434 18368 12440 18420
rect 12492 18408 12498 18420
rect 12492 18380 12537 18408
rect 12492 18368 12498 18380
rect 13538 18368 13544 18420
rect 13596 18408 13602 18420
rect 15654 18408 15660 18420
rect 13596 18380 15660 18408
rect 13596 18368 13602 18380
rect 15654 18368 15660 18380
rect 15712 18368 15718 18420
rect 16393 18411 16451 18417
rect 16393 18377 16405 18411
rect 16439 18408 16451 18411
rect 17126 18408 17132 18420
rect 16439 18380 17132 18408
rect 16439 18377 16451 18380
rect 16393 18371 16451 18377
rect 17126 18368 17132 18380
rect 17184 18368 17190 18420
rect 4632 18312 6868 18340
rect 10410 18300 10416 18352
rect 10468 18340 10474 18352
rect 10962 18340 10968 18352
rect 10468 18312 10968 18340
rect 10468 18300 10474 18312
rect 10962 18300 10968 18312
rect 11020 18300 11026 18352
rect 14001 18343 14059 18349
rect 14001 18309 14013 18343
rect 14047 18309 14059 18343
rect 14001 18303 14059 18309
rect 2409 18275 2467 18281
rect 2409 18241 2421 18275
rect 2455 18241 2467 18275
rect 3326 18272 3332 18284
rect 3287 18244 3332 18272
rect 2409 18235 2467 18241
rect 3326 18232 3332 18244
rect 3384 18232 3390 18284
rect 6546 18232 6552 18284
rect 6604 18272 6610 18284
rect 6825 18275 6883 18281
rect 6825 18272 6837 18275
rect 6604 18244 6837 18272
rect 6604 18232 6610 18244
rect 6825 18241 6837 18244
rect 6871 18241 6883 18275
rect 12894 18272 12900 18284
rect 6825 18235 6883 18241
rect 10888 18244 12900 18272
rect 1762 18164 1768 18216
rect 1820 18204 1826 18216
rect 2133 18207 2191 18213
rect 2133 18204 2145 18207
rect 1820 18176 2145 18204
rect 1820 18164 1826 18176
rect 2133 18173 2145 18176
rect 2179 18173 2191 18207
rect 2133 18167 2191 18173
rect 3970 18164 3976 18216
rect 4028 18204 4034 18216
rect 5537 18207 5595 18213
rect 4028 18176 4384 18204
rect 4028 18164 4034 18176
rect 3050 18096 3056 18148
rect 3108 18136 3114 18148
rect 3574 18139 3632 18145
rect 3574 18136 3586 18139
rect 3108 18108 3586 18136
rect 3108 18096 3114 18108
rect 3574 18105 3586 18108
rect 3620 18136 3632 18139
rect 4246 18136 4252 18148
rect 3620 18108 4252 18136
rect 3620 18105 3632 18108
rect 3574 18099 3632 18105
rect 4246 18096 4252 18108
rect 4304 18096 4310 18148
rect 4356 18136 4384 18176
rect 5537 18173 5549 18207
rect 5583 18204 5595 18207
rect 5626 18204 5632 18216
rect 5583 18176 5632 18204
rect 5583 18173 5595 18176
rect 5537 18167 5595 18173
rect 5626 18164 5632 18176
rect 5684 18164 5690 18216
rect 5718 18164 5724 18216
rect 5776 18204 5782 18216
rect 5776 18176 6776 18204
rect 5776 18164 5782 18176
rect 4356 18108 5764 18136
rect 198 18028 204 18080
rect 256 18068 262 18080
rect 1302 18068 1308 18080
rect 256 18040 1308 18068
rect 256 18028 262 18040
rect 1302 18028 1308 18040
rect 1360 18028 1366 18080
rect 1765 18071 1823 18077
rect 1765 18037 1777 18071
rect 1811 18068 1823 18071
rect 5534 18068 5540 18080
rect 1811 18040 5540 18068
rect 1811 18037 1823 18040
rect 1765 18031 1823 18037
rect 5534 18028 5540 18040
rect 5592 18028 5598 18080
rect 5736 18077 5764 18108
rect 5721 18071 5779 18077
rect 5721 18037 5733 18071
rect 5767 18037 5779 18071
rect 6748 18068 6776 18176
rect 6914 18164 6920 18216
rect 6972 18204 6978 18216
rect 9401 18207 9459 18213
rect 6972 18176 9352 18204
rect 6972 18164 6978 18176
rect 7081 18139 7139 18145
rect 7081 18105 7093 18139
rect 7127 18136 7139 18139
rect 7190 18136 7196 18148
rect 7127 18108 7196 18136
rect 7127 18105 7139 18108
rect 7081 18099 7139 18105
rect 7190 18096 7196 18108
rect 7248 18096 7254 18148
rect 9214 18136 9220 18148
rect 8036 18108 9220 18136
rect 8036 18068 8064 18108
rect 9214 18096 9220 18108
rect 9272 18096 9278 18148
rect 9324 18136 9352 18176
rect 9401 18173 9413 18207
rect 9447 18204 9459 18207
rect 9490 18204 9496 18216
rect 9447 18176 9496 18204
rect 9447 18173 9459 18176
rect 9401 18167 9459 18173
rect 9490 18164 9496 18176
rect 9548 18164 9554 18216
rect 9668 18207 9726 18213
rect 9668 18173 9680 18207
rect 9714 18204 9726 18207
rect 10778 18204 10784 18216
rect 9714 18176 10784 18204
rect 9714 18173 9726 18176
rect 9668 18167 9726 18173
rect 10778 18164 10784 18176
rect 10836 18164 10842 18216
rect 10888 18136 10916 18244
rect 12894 18232 12900 18244
rect 12952 18232 12958 18284
rect 13081 18275 13139 18281
rect 13081 18241 13093 18275
rect 13127 18272 13139 18275
rect 13262 18272 13268 18284
rect 13127 18244 13268 18272
rect 13127 18241 13139 18244
rect 13081 18235 13139 18241
rect 13262 18232 13268 18244
rect 13320 18232 13326 18284
rect 10962 18164 10968 18216
rect 11020 18204 11026 18216
rect 14016 18204 14044 18303
rect 14642 18272 14648 18284
rect 14603 18244 14648 18272
rect 14642 18232 14648 18244
rect 14700 18232 14706 18284
rect 16942 18272 16948 18284
rect 16903 18244 16948 18272
rect 16942 18232 16948 18244
rect 17000 18232 17006 18284
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18785 18275 18843 18281
rect 18785 18272 18797 18275
rect 18012 18244 18797 18272
rect 18012 18232 18018 18244
rect 18785 18241 18797 18244
rect 18831 18241 18843 18275
rect 18785 18235 18843 18241
rect 11020 18176 14044 18204
rect 11020 18164 11026 18176
rect 9324 18108 10916 18136
rect 12805 18139 12863 18145
rect 12805 18105 12817 18139
rect 12851 18136 12863 18139
rect 13538 18136 13544 18148
rect 12851 18108 13544 18136
rect 12851 18105 12863 18108
rect 12805 18099 12863 18105
rect 13538 18096 13544 18108
rect 13596 18096 13602 18148
rect 13630 18096 13636 18148
rect 13688 18136 13694 18148
rect 14461 18139 14519 18145
rect 14461 18136 14473 18139
rect 13688 18108 14473 18136
rect 13688 18096 13694 18108
rect 14461 18105 14473 18108
rect 14507 18105 14519 18139
rect 14461 18099 14519 18105
rect 16761 18139 16819 18145
rect 16761 18105 16773 18139
rect 16807 18136 16819 18139
rect 17770 18136 17776 18148
rect 16807 18108 17776 18136
rect 16807 18105 16819 18108
rect 16761 18099 16819 18105
rect 17770 18096 17776 18108
rect 17828 18096 17834 18148
rect 18800 18136 18828 18235
rect 19052 18207 19110 18213
rect 19052 18173 19064 18207
rect 19098 18204 19110 18207
rect 19886 18204 19892 18216
rect 19098 18176 19892 18204
rect 19098 18173 19110 18176
rect 19052 18167 19110 18173
rect 19886 18164 19892 18176
rect 19944 18164 19950 18216
rect 18966 18136 18972 18148
rect 18800 18108 18972 18136
rect 18966 18096 18972 18108
rect 19024 18096 19030 18148
rect 8202 18068 8208 18080
rect 6748 18040 8064 18068
rect 8163 18040 8208 18068
rect 5721 18031 5779 18037
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 9122 18028 9128 18080
rect 9180 18068 9186 18080
rect 10318 18068 10324 18080
rect 9180 18040 10324 18068
rect 9180 18028 9186 18040
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 10686 18028 10692 18080
rect 10744 18068 10750 18080
rect 10781 18071 10839 18077
rect 10781 18068 10793 18071
rect 10744 18040 10793 18068
rect 10744 18028 10750 18040
rect 10781 18037 10793 18040
rect 10827 18037 10839 18071
rect 10781 18031 10839 18037
rect 12897 18071 12955 18077
rect 12897 18037 12909 18071
rect 12943 18068 12955 18071
rect 13814 18068 13820 18080
rect 12943 18040 13820 18068
rect 12943 18037 12955 18040
rect 12897 18031 12955 18037
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 13906 18028 13912 18080
rect 13964 18068 13970 18080
rect 14369 18071 14427 18077
rect 14369 18068 14381 18071
rect 13964 18040 14381 18068
rect 13964 18028 13970 18040
rect 14369 18037 14381 18040
rect 14415 18037 14427 18071
rect 14369 18031 14427 18037
rect 14550 18028 14556 18080
rect 14608 18068 14614 18080
rect 16853 18071 16911 18077
rect 16853 18068 16865 18071
rect 14608 18040 16865 18068
rect 14608 18028 14614 18040
rect 16853 18037 16865 18040
rect 16899 18068 16911 18071
rect 16942 18068 16948 18080
rect 16899 18040 16948 18068
rect 16899 18037 16911 18040
rect 16853 18031 16911 18037
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 20162 18068 20168 18080
rect 20123 18040 20168 18068
rect 20162 18028 20168 18040
rect 20220 18028 20226 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 2409 17867 2467 17873
rect 2409 17833 2421 17867
rect 2455 17864 2467 17867
rect 4154 17864 4160 17876
rect 2455 17836 4160 17864
rect 2455 17833 2467 17836
rect 2409 17827 2467 17833
rect 4154 17824 4160 17836
rect 4212 17824 4218 17876
rect 5813 17867 5871 17873
rect 5813 17833 5825 17867
rect 5859 17864 5871 17867
rect 7190 17864 7196 17876
rect 5859 17836 7196 17864
rect 5859 17833 5871 17836
rect 5813 17827 5871 17833
rect 7190 17824 7196 17836
rect 7248 17864 7254 17876
rect 9674 17864 9680 17876
rect 7248 17836 8340 17864
rect 9635 17836 9680 17864
rect 7248 17824 7254 17836
rect 3878 17756 3884 17808
rect 3936 17796 3942 17808
rect 4700 17799 4758 17805
rect 3936 17768 4476 17796
rect 3936 17756 3942 17768
rect 2777 17731 2835 17737
rect 2777 17697 2789 17731
rect 2823 17728 2835 17731
rect 4338 17728 4344 17740
rect 2823 17700 4344 17728
rect 2823 17697 2835 17700
rect 2777 17691 2835 17697
rect 4338 17688 4344 17700
rect 4396 17688 4402 17740
rect 4448 17728 4476 17768
rect 4700 17765 4712 17799
rect 4746 17796 4758 17799
rect 4798 17796 4804 17808
rect 4746 17768 4804 17796
rect 4746 17765 4758 17768
rect 4700 17759 4758 17765
rect 4798 17756 4804 17768
rect 4856 17756 4862 17808
rect 5350 17756 5356 17808
rect 5408 17796 5414 17808
rect 6178 17796 6184 17808
rect 5408 17768 6184 17796
rect 5408 17756 5414 17768
rect 6178 17756 6184 17768
rect 6236 17756 6242 17808
rect 6270 17756 6276 17808
rect 6328 17796 6334 17808
rect 6730 17796 6736 17808
rect 6328 17768 6736 17796
rect 6328 17756 6334 17768
rect 6730 17756 6736 17768
rect 6788 17756 6794 17808
rect 6908 17799 6966 17805
rect 6908 17765 6920 17799
rect 6954 17796 6966 17799
rect 8202 17796 8208 17808
rect 6954 17768 8208 17796
rect 6954 17765 6966 17768
rect 6908 17759 6966 17765
rect 8202 17756 8208 17768
rect 8260 17756 8266 17808
rect 8312 17796 8340 17836
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 10137 17867 10195 17873
rect 10137 17833 10149 17867
rect 10183 17864 10195 17867
rect 10226 17864 10232 17876
rect 10183 17836 10232 17864
rect 10183 17833 10195 17836
rect 10137 17827 10195 17833
rect 10226 17824 10232 17836
rect 10284 17824 10290 17876
rect 11698 17824 11704 17876
rect 11756 17864 11762 17876
rect 12989 17867 13047 17873
rect 12989 17864 13001 17867
rect 11756 17836 13001 17864
rect 11756 17824 11762 17836
rect 12989 17833 13001 17836
rect 13035 17833 13047 17867
rect 12989 17827 13047 17833
rect 13262 17824 13268 17876
rect 13320 17864 13326 17876
rect 15657 17867 15715 17873
rect 15657 17864 15669 17867
rect 13320 17836 15669 17864
rect 13320 17824 13326 17836
rect 15657 17833 15669 17836
rect 15703 17833 15715 17867
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 15657 17827 15715 17833
rect 15856 17836 19717 17864
rect 8312 17768 10272 17796
rect 8110 17728 8116 17740
rect 4448 17700 8116 17728
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 9950 17688 9956 17740
rect 10008 17728 10014 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 10008 17700 10057 17728
rect 10008 17688 10014 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17660 1455 17663
rect 2406 17660 2412 17672
rect 1443 17632 2412 17660
rect 1443 17629 1455 17632
rect 1397 17623 1455 17629
rect 2406 17620 2412 17632
rect 2464 17620 2470 17672
rect 2498 17620 2504 17672
rect 2556 17660 2562 17672
rect 2869 17663 2927 17669
rect 2869 17660 2881 17663
rect 2556 17632 2881 17660
rect 2556 17620 2562 17632
rect 2869 17629 2881 17632
rect 2915 17629 2927 17663
rect 3050 17660 3056 17672
rect 3011 17632 3056 17660
rect 2869 17623 2927 17629
rect 3050 17620 3056 17632
rect 3108 17620 3114 17672
rect 3326 17620 3332 17672
rect 3384 17660 3390 17672
rect 4433 17663 4491 17669
rect 4433 17660 4445 17663
rect 3384 17632 4445 17660
rect 3384 17620 3390 17632
rect 4433 17629 4445 17632
rect 4479 17629 4491 17663
rect 4433 17623 4491 17629
rect 4448 17524 4476 17623
rect 6546 17620 6552 17672
rect 6604 17660 6610 17672
rect 6641 17663 6699 17669
rect 6641 17660 6653 17663
rect 6604 17632 6653 17660
rect 6604 17620 6610 17632
rect 6641 17629 6653 17632
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 7650 17620 7656 17672
rect 7708 17660 7714 17672
rect 10134 17660 10140 17672
rect 7708 17632 10140 17660
rect 7708 17620 7714 17632
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 10244 17669 10272 17768
rect 10410 17756 10416 17808
rect 10468 17796 10474 17808
rect 12710 17796 12716 17808
rect 10468 17768 12716 17796
rect 10468 17756 10474 17768
rect 12710 17756 12716 17768
rect 12768 17756 12774 17808
rect 12894 17756 12900 17808
rect 12952 17796 12958 17808
rect 14093 17799 14151 17805
rect 14093 17796 14105 17799
rect 12952 17768 14105 17796
rect 12952 17756 12958 17768
rect 14093 17765 14105 17768
rect 14139 17765 14151 17799
rect 14093 17759 14151 17765
rect 15194 17756 15200 17808
rect 15252 17796 15258 17808
rect 15749 17799 15807 17805
rect 15749 17796 15761 17799
rect 15252 17768 15761 17796
rect 15252 17756 15258 17768
rect 15749 17765 15761 17768
rect 15795 17765 15807 17799
rect 15749 17759 15807 17765
rect 11882 17737 11888 17740
rect 11876 17728 11888 17737
rect 11843 17700 11888 17728
rect 11876 17691 11888 17700
rect 11882 17688 11888 17691
rect 11940 17688 11946 17740
rect 12342 17688 12348 17740
rect 12400 17728 12406 17740
rect 12400 17700 12756 17728
rect 12400 17688 12406 17700
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17629 10287 17663
rect 10229 17623 10287 17629
rect 11054 17620 11060 17672
rect 11112 17660 11118 17672
rect 11609 17663 11667 17669
rect 11609 17660 11621 17663
rect 11112 17632 11621 17660
rect 11112 17620 11118 17632
rect 11609 17629 11621 17632
rect 11655 17629 11667 17663
rect 12728 17660 12756 17700
rect 12802 17688 12808 17740
rect 12860 17728 12866 17740
rect 13817 17731 13875 17737
rect 13817 17728 13829 17731
rect 12860 17700 13829 17728
rect 12860 17688 12866 17700
rect 13817 17697 13829 17700
rect 13863 17697 13875 17731
rect 13817 17691 13875 17697
rect 14366 17688 14372 17740
rect 14424 17728 14430 17740
rect 15856 17728 15884 17836
rect 19705 17833 19717 17836
rect 19751 17833 19763 17867
rect 19705 17827 19763 17833
rect 15930 17756 15936 17808
rect 15988 17756 15994 17808
rect 17586 17756 17592 17808
rect 17644 17796 17650 17808
rect 18141 17799 18199 17805
rect 18141 17796 18153 17799
rect 17644 17768 18153 17796
rect 17644 17756 17650 17768
rect 18141 17765 18153 17768
rect 18187 17765 18199 17799
rect 18141 17759 18199 17765
rect 14424 17700 15884 17728
rect 15948 17728 15976 17756
rect 17954 17728 17960 17740
rect 15948 17700 17960 17728
rect 14424 17688 14430 17700
rect 17954 17688 17960 17700
rect 18012 17728 18018 17740
rect 18049 17731 18107 17737
rect 18049 17728 18061 17731
rect 18012 17700 18061 17728
rect 18012 17688 18018 17700
rect 18049 17697 18061 17700
rect 18095 17697 18107 17731
rect 18049 17691 18107 17697
rect 18598 17688 18604 17740
rect 18656 17728 18662 17740
rect 19613 17731 19671 17737
rect 19613 17728 19625 17731
rect 18656 17700 19625 17728
rect 18656 17688 18662 17700
rect 19613 17697 19625 17700
rect 19659 17697 19671 17731
rect 19613 17691 19671 17697
rect 15010 17660 15016 17672
rect 12728 17632 15016 17660
rect 11609 17623 11667 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15194 17620 15200 17672
rect 15252 17660 15258 17672
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 15252 17632 15853 17660
rect 15252 17620 15258 17632
rect 15841 17629 15853 17632
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 18325 17663 18383 17669
rect 18325 17629 18337 17663
rect 18371 17629 18383 17663
rect 18325 17623 18383 17629
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 6564 17524 6592 17620
rect 8478 17552 8484 17604
rect 8536 17592 8542 17604
rect 11514 17592 11520 17604
rect 8536 17564 11520 17592
rect 8536 17552 8542 17564
rect 11514 17552 11520 17564
rect 11572 17552 11578 17604
rect 12618 17552 12624 17604
rect 12676 17592 12682 17604
rect 15289 17595 15347 17601
rect 15289 17592 15301 17595
rect 12676 17564 15301 17592
rect 12676 17552 12682 17564
rect 15289 17561 15301 17564
rect 15335 17561 15347 17595
rect 18340 17592 18368 17623
rect 18782 17592 18788 17604
rect 18340 17564 18788 17592
rect 15289 17555 15347 17561
rect 18782 17552 18788 17564
rect 18840 17592 18846 17604
rect 19812 17592 19840 17623
rect 20530 17620 20536 17672
rect 20588 17660 20594 17672
rect 20806 17660 20812 17672
rect 20588 17632 20812 17660
rect 20588 17620 20594 17632
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 20438 17592 20444 17604
rect 18840 17564 20444 17592
rect 18840 17552 18846 17564
rect 20438 17552 20444 17564
rect 20496 17552 20502 17604
rect 4448 17496 6592 17524
rect 6822 17484 6828 17536
rect 6880 17524 6886 17536
rect 8021 17527 8079 17533
rect 8021 17524 8033 17527
rect 6880 17496 8033 17524
rect 6880 17484 6886 17496
rect 8021 17493 8033 17496
rect 8067 17493 8079 17527
rect 8021 17487 8079 17493
rect 8110 17484 8116 17536
rect 8168 17524 8174 17536
rect 10226 17524 10232 17536
rect 8168 17496 10232 17524
rect 8168 17484 8174 17496
rect 10226 17484 10232 17496
rect 10284 17484 10290 17536
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 15194 17524 15200 17536
rect 12584 17496 15200 17524
rect 12584 17484 12590 17496
rect 15194 17484 15200 17496
rect 15252 17484 15258 17536
rect 17678 17524 17684 17536
rect 17639 17496 17684 17524
rect 17678 17484 17684 17496
rect 17736 17484 17742 17536
rect 19150 17484 19156 17536
rect 19208 17524 19214 17536
rect 19245 17527 19303 17533
rect 19245 17524 19257 17527
rect 19208 17496 19257 17524
rect 19208 17484 19214 17496
rect 19245 17493 19257 17496
rect 19291 17493 19303 17527
rect 19245 17487 19303 17493
rect 20806 17484 20812 17536
rect 20864 17524 20870 17536
rect 21818 17524 21824 17536
rect 20864 17496 21824 17524
rect 20864 17484 20870 17496
rect 21818 17484 21824 17496
rect 21876 17484 21882 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 3326 17320 3332 17332
rect 2332 17292 3332 17320
rect 2332 17193 2360 17292
rect 3326 17280 3332 17292
rect 3384 17280 3390 17332
rect 3694 17320 3700 17332
rect 3655 17292 3700 17320
rect 3694 17280 3700 17292
rect 3752 17280 3758 17332
rect 4338 17280 4344 17332
rect 4396 17320 4402 17332
rect 4525 17323 4583 17329
rect 4525 17320 4537 17323
rect 4396 17292 4537 17320
rect 4396 17280 4402 17292
rect 4525 17289 4537 17292
rect 4571 17289 4583 17323
rect 4525 17283 4583 17289
rect 5350 17280 5356 17332
rect 5408 17320 5414 17332
rect 7650 17320 7656 17332
rect 5408 17292 7656 17320
rect 5408 17280 5414 17292
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 9306 17320 9312 17332
rect 8220 17292 9312 17320
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17153 2375 17187
rect 3712 17184 3740 17280
rect 3786 17212 3792 17264
rect 3844 17252 3850 17264
rect 8220 17252 8248 17292
rect 9306 17280 9312 17292
rect 9364 17280 9370 17332
rect 9582 17280 9588 17332
rect 9640 17320 9646 17332
rect 12526 17320 12532 17332
rect 9640 17292 12532 17320
rect 9640 17280 9646 17292
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 17954 17280 17960 17332
rect 18012 17280 18018 17332
rect 18966 17280 18972 17332
rect 19024 17280 19030 17332
rect 20438 17320 20444 17332
rect 20399 17292 20444 17320
rect 20438 17280 20444 17292
rect 20496 17280 20502 17332
rect 20898 17280 20904 17332
rect 20956 17320 20962 17332
rect 21174 17320 21180 17332
rect 20956 17292 21180 17320
rect 20956 17280 20962 17292
rect 21174 17280 21180 17292
rect 21232 17280 21238 17332
rect 3844 17224 8248 17252
rect 8297 17255 8355 17261
rect 3844 17212 3850 17224
rect 8297 17221 8309 17255
rect 8343 17252 8355 17255
rect 10134 17252 10140 17264
rect 8343 17224 10140 17252
rect 8343 17221 8355 17224
rect 8297 17215 8355 17221
rect 10134 17212 10140 17224
rect 10192 17212 10198 17264
rect 10226 17212 10232 17264
rect 10284 17252 10290 17264
rect 13814 17252 13820 17264
rect 10284 17224 13820 17252
rect 10284 17212 10290 17224
rect 13814 17212 13820 17224
rect 13872 17212 13878 17264
rect 16209 17255 16267 17261
rect 16209 17221 16221 17255
rect 16255 17252 16267 17255
rect 16255 17224 17816 17252
rect 16255 17221 16267 17224
rect 16209 17215 16267 17221
rect 5077 17187 5135 17193
rect 5077 17184 5089 17187
rect 3712 17156 5089 17184
rect 2317 17147 2375 17153
rect 5077 17153 5089 17156
rect 5123 17153 5135 17187
rect 5077 17147 5135 17153
rect 7374 17144 7380 17196
rect 7432 17184 7438 17196
rect 8757 17187 8815 17193
rect 8757 17184 8769 17187
rect 7432 17156 8769 17184
rect 7432 17144 7438 17156
rect 8757 17153 8769 17156
rect 8803 17153 8815 17187
rect 8757 17147 8815 17153
rect 8941 17187 8999 17193
rect 8941 17153 8953 17187
rect 8987 17184 8999 17187
rect 10686 17184 10692 17196
rect 8987 17156 10692 17184
rect 8987 17153 8999 17156
rect 8941 17147 8999 17153
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 13081 17187 13139 17193
rect 13081 17153 13093 17187
rect 13127 17184 13139 17187
rect 13354 17184 13360 17196
rect 13127 17156 13360 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 13354 17144 13360 17156
rect 13412 17144 13418 17196
rect 15010 17144 15016 17196
rect 15068 17184 15074 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 15068 17156 16681 17184
rect 15068 17144 15074 17156
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 16761 17187 16819 17193
rect 16761 17153 16773 17187
rect 16807 17153 16819 17187
rect 16761 17147 16819 17153
rect 2406 17076 2412 17128
rect 2464 17116 2470 17128
rect 4893 17119 4951 17125
rect 4893 17116 4905 17119
rect 2464 17088 4905 17116
rect 2464 17076 2470 17088
rect 4893 17085 4905 17088
rect 4939 17085 4951 17119
rect 4893 17079 4951 17085
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17116 7067 17119
rect 13722 17116 13728 17128
rect 7055 17088 13728 17116
rect 7055 17085 7067 17088
rect 7009 17079 7067 17085
rect 13722 17076 13728 17088
rect 13780 17076 13786 17128
rect 13998 17116 14004 17128
rect 13959 17088 14004 17116
rect 13998 17076 14004 17088
rect 14056 17076 14062 17128
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 16776 17116 16804 17147
rect 14148 17088 16804 17116
rect 17788 17116 17816 17224
rect 17862 17144 17868 17196
rect 17920 17184 17926 17196
rect 17972 17184 18000 17280
rect 17920 17156 18000 17184
rect 18049 17187 18107 17193
rect 17920 17144 17926 17156
rect 18049 17153 18061 17187
rect 18095 17184 18107 17187
rect 18598 17184 18604 17196
rect 18095 17156 18604 17184
rect 18095 17153 18107 17156
rect 18049 17147 18107 17153
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 18984 17184 19012 17280
rect 19061 17187 19119 17193
rect 19061 17184 19073 17187
rect 18984 17156 19073 17184
rect 19061 17153 19073 17156
rect 19107 17153 19119 17187
rect 19061 17147 19119 17153
rect 20898 17144 20904 17196
rect 20956 17184 20962 17196
rect 22278 17184 22284 17196
rect 20956 17156 22284 17184
rect 20956 17144 20962 17156
rect 22278 17144 22284 17156
rect 22336 17144 22342 17196
rect 18690 17116 18696 17128
rect 17788 17088 18696 17116
rect 14148 17076 14154 17088
rect 18690 17076 18696 17088
rect 18748 17076 18754 17128
rect 19328 17119 19386 17125
rect 19328 17085 19340 17119
rect 19374 17116 19386 17119
rect 20162 17116 20168 17128
rect 19374 17088 20168 17116
rect 19374 17085 19386 17088
rect 19328 17079 19386 17085
rect 20162 17076 20168 17088
rect 20220 17076 20226 17128
rect 2584 17051 2642 17057
rect 2584 17017 2596 17051
rect 2630 17048 2642 17051
rect 3050 17048 3056 17060
rect 2630 17020 3056 17048
rect 2630 17017 2642 17020
rect 2584 17011 2642 17017
rect 3050 17008 3056 17020
rect 3108 17008 3114 17060
rect 7285 17051 7343 17057
rect 7285 17048 7297 17051
rect 7024 17020 7297 17048
rect 7024 16992 7052 17020
rect 7285 17017 7297 17020
rect 7331 17017 7343 17051
rect 7285 17011 7343 17017
rect 8294 17008 8300 17060
rect 8352 17048 8358 17060
rect 8665 17051 8723 17057
rect 8665 17048 8677 17051
rect 8352 17020 8677 17048
rect 8352 17008 8358 17020
rect 8665 17017 8677 17020
rect 8711 17048 8723 17051
rect 9398 17048 9404 17060
rect 8711 17020 9404 17048
rect 8711 17017 8723 17020
rect 8665 17011 8723 17017
rect 9398 17008 9404 17020
rect 9456 17008 9462 17060
rect 10505 17051 10563 17057
rect 10505 17048 10517 17051
rect 9508 17020 10517 17048
rect 4798 16940 4804 16992
rect 4856 16980 4862 16992
rect 4985 16983 5043 16989
rect 4985 16980 4997 16983
rect 4856 16952 4997 16980
rect 4856 16940 4862 16952
rect 4985 16949 4997 16952
rect 5031 16949 5043 16983
rect 4985 16943 5043 16949
rect 7006 16940 7012 16992
rect 7064 16940 7070 16992
rect 7190 16940 7196 16992
rect 7248 16980 7254 16992
rect 9508 16980 9536 17020
rect 10505 17017 10517 17020
rect 10551 17017 10563 17051
rect 10505 17011 10563 17017
rect 11698 17008 11704 17060
rect 11756 17048 11762 17060
rect 11756 17020 12664 17048
rect 11756 17008 11762 17020
rect 7248 16952 9536 16980
rect 10045 16983 10103 16989
rect 7248 16940 7254 16952
rect 10045 16949 10057 16983
rect 10091 16980 10103 16983
rect 10318 16980 10324 16992
rect 10091 16952 10324 16980
rect 10091 16949 10103 16952
rect 10045 16943 10103 16949
rect 10318 16940 10324 16952
rect 10376 16940 10382 16992
rect 10413 16983 10471 16989
rect 10413 16949 10425 16983
rect 10459 16980 10471 16983
rect 10870 16980 10876 16992
rect 10459 16952 10876 16980
rect 10459 16949 10471 16952
rect 10413 16943 10471 16949
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 12437 16983 12495 16989
rect 12437 16949 12449 16983
rect 12483 16980 12495 16983
rect 12526 16980 12532 16992
rect 12483 16952 12532 16980
rect 12483 16949 12495 16952
rect 12437 16943 12495 16949
rect 12526 16940 12532 16952
rect 12584 16940 12590 16992
rect 12636 16980 12664 17020
rect 12710 17008 12716 17060
rect 12768 17048 12774 17060
rect 12897 17051 12955 17057
rect 12897 17048 12909 17051
rect 12768 17020 12909 17048
rect 12768 17008 12774 17020
rect 12897 17017 12909 17020
rect 12943 17017 12955 17051
rect 12897 17011 12955 17017
rect 14182 17008 14188 17060
rect 14240 17057 14246 17060
rect 14240 17051 14304 17057
rect 14240 17017 14258 17051
rect 14292 17017 14304 17051
rect 14240 17011 14304 17017
rect 14240 17008 14246 17011
rect 12805 16983 12863 16989
rect 12805 16980 12817 16983
rect 12636 16952 12817 16980
rect 12805 16949 12817 16952
rect 12851 16949 12863 16983
rect 12805 16943 12863 16949
rect 14642 16940 14648 16992
rect 14700 16980 14706 16992
rect 15381 16983 15439 16989
rect 15381 16980 15393 16983
rect 14700 16952 15393 16980
rect 14700 16940 14706 16952
rect 15381 16949 15393 16952
rect 15427 16949 15439 16983
rect 15381 16943 15439 16949
rect 15930 16940 15936 16992
rect 15988 16980 15994 16992
rect 16206 16980 16212 16992
rect 15988 16952 16212 16980
rect 15988 16940 15994 16952
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 16298 16940 16304 16992
rect 16356 16980 16362 16992
rect 16577 16983 16635 16989
rect 16577 16980 16589 16983
rect 16356 16952 16589 16980
rect 16356 16940 16362 16952
rect 16577 16949 16589 16952
rect 16623 16949 16635 16983
rect 16577 16943 16635 16949
rect 17954 16940 17960 16992
rect 18012 16980 18018 16992
rect 18598 16980 18604 16992
rect 18012 16952 18604 16980
rect 18012 16940 18018 16952
rect 18598 16940 18604 16952
rect 18656 16940 18662 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 2409 16779 2467 16785
rect 2409 16745 2421 16779
rect 2455 16776 2467 16779
rect 2498 16776 2504 16788
rect 2455 16748 2504 16776
rect 2455 16745 2467 16748
rect 2409 16739 2467 16745
rect 2498 16736 2504 16748
rect 2556 16736 2562 16788
rect 4154 16736 4160 16788
rect 4212 16776 4218 16788
rect 8665 16779 8723 16785
rect 8665 16776 8677 16779
rect 4212 16748 8677 16776
rect 4212 16736 4218 16748
rect 8665 16745 8677 16748
rect 8711 16745 8723 16779
rect 8665 16739 8723 16745
rect 10505 16779 10563 16785
rect 10505 16745 10517 16779
rect 10551 16776 10563 16779
rect 10962 16776 10968 16788
rect 10551 16748 10968 16776
rect 10551 16745 10563 16748
rect 10505 16739 10563 16745
rect 10962 16736 10968 16748
rect 11020 16736 11026 16788
rect 11974 16776 11980 16788
rect 11935 16748 11980 16776
rect 11974 16736 11980 16748
rect 12032 16736 12038 16788
rect 12802 16776 12808 16788
rect 12763 16748 12808 16776
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 13265 16779 13323 16785
rect 13265 16745 13277 16779
rect 13311 16776 13323 16779
rect 13311 16748 13400 16776
rect 13311 16745 13323 16748
rect 13265 16739 13323 16745
rect 2777 16711 2835 16717
rect 2777 16677 2789 16711
rect 2823 16708 2835 16711
rect 2866 16708 2872 16720
rect 2823 16680 2872 16708
rect 2823 16677 2835 16680
rect 2777 16671 2835 16677
rect 2866 16668 2872 16680
rect 2924 16668 2930 16720
rect 5350 16708 5356 16720
rect 3896 16680 5356 16708
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 1486 16640 1492 16652
rect 1443 16612 1492 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 1486 16600 1492 16612
rect 1544 16640 1550 16652
rect 1673 16643 1731 16649
rect 1673 16640 1685 16643
rect 1544 16612 1685 16640
rect 1544 16600 1550 16612
rect 1673 16609 1685 16612
rect 1719 16609 1731 16643
rect 3896 16640 3924 16680
rect 5350 16668 5356 16680
rect 5408 16668 5414 16720
rect 5721 16711 5779 16717
rect 5721 16677 5733 16711
rect 5767 16708 5779 16711
rect 6270 16708 6276 16720
rect 5767 16680 6276 16708
rect 5767 16677 5779 16680
rect 5721 16671 5779 16677
rect 6270 16668 6276 16680
rect 6328 16668 6334 16720
rect 13372 16708 13400 16748
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 18785 16779 18843 16785
rect 18785 16776 18797 16779
rect 13780 16748 18797 16776
rect 13780 16736 13786 16748
rect 18785 16745 18797 16748
rect 18831 16745 18843 16779
rect 19150 16776 19156 16788
rect 19111 16748 19156 16776
rect 18785 16739 18843 16745
rect 19150 16736 19156 16748
rect 19208 16736 19214 16788
rect 13538 16708 13544 16720
rect 7208 16680 11652 16708
rect 13372 16680 13544 16708
rect 4062 16640 4068 16652
rect 1673 16603 1731 16609
rect 2884 16612 3924 16640
rect 4023 16612 4068 16640
rect 2884 16581 2912 16612
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 4341 16643 4399 16649
rect 4341 16609 4353 16643
rect 4387 16640 4399 16643
rect 7208 16640 7236 16680
rect 4387 16612 5764 16640
rect 4387 16609 4399 16612
rect 4341 16603 4399 16609
rect 5736 16584 5764 16612
rect 5828 16612 7236 16640
rect 7285 16643 7343 16649
rect 2869 16575 2927 16581
rect 2869 16541 2881 16575
rect 2915 16541 2927 16575
rect 2869 16535 2927 16541
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16572 3111 16575
rect 3694 16572 3700 16584
rect 3099 16544 3700 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 3694 16532 3700 16544
rect 3752 16532 3758 16584
rect 5718 16532 5724 16584
rect 5776 16532 5782 16584
rect 5828 16581 5856 16612
rect 7285 16609 7297 16643
rect 7331 16640 7343 16643
rect 8294 16640 8300 16652
rect 7331 16612 8300 16640
rect 7331 16609 7343 16612
rect 7285 16603 7343 16609
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16640 8539 16643
rect 9214 16640 9220 16652
rect 8527 16612 9220 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 9582 16600 9588 16652
rect 9640 16640 9646 16652
rect 10853 16643 10911 16649
rect 10853 16640 10865 16643
rect 9640 16612 10865 16640
rect 9640 16600 9646 16612
rect 10853 16609 10865 16612
rect 10899 16609 10911 16643
rect 10853 16603 10911 16609
rect 5813 16575 5871 16581
rect 5813 16541 5825 16575
rect 5859 16541 5871 16575
rect 5813 16535 5871 16541
rect 5997 16575 6055 16581
rect 5997 16541 6009 16575
rect 6043 16541 6055 16575
rect 7374 16572 7380 16584
rect 7335 16544 7380 16572
rect 5997 16535 6055 16541
rect 1854 16464 1860 16516
rect 1912 16504 1918 16516
rect 3786 16504 3792 16516
rect 1912 16476 3792 16504
rect 1912 16464 1918 16476
rect 3786 16464 3792 16476
rect 3844 16464 3850 16516
rect 5442 16464 5448 16516
rect 5500 16504 5506 16516
rect 6012 16504 6040 16535
rect 7374 16532 7380 16544
rect 7432 16532 7438 16584
rect 7469 16575 7527 16581
rect 7469 16541 7481 16575
rect 7515 16541 7527 16575
rect 7469 16535 7527 16541
rect 10505 16575 10563 16581
rect 10505 16541 10517 16575
rect 10551 16572 10563 16575
rect 10597 16575 10655 16581
rect 10597 16572 10609 16575
rect 10551 16544 10609 16572
rect 10551 16541 10563 16544
rect 10505 16535 10563 16541
rect 10597 16541 10609 16544
rect 10643 16541 10655 16575
rect 10597 16535 10655 16541
rect 7484 16504 7512 16535
rect 5500 16476 7512 16504
rect 5500 16464 5506 16476
rect 5350 16436 5356 16448
rect 5311 16408 5356 16436
rect 5350 16396 5356 16408
rect 5408 16396 5414 16448
rect 5534 16396 5540 16448
rect 5592 16436 5598 16448
rect 6917 16439 6975 16445
rect 6917 16436 6929 16439
rect 5592 16408 6929 16436
rect 5592 16396 5598 16408
rect 6917 16405 6929 16408
rect 6963 16405 6975 16439
rect 6917 16399 6975 16405
rect 8110 16396 8116 16448
rect 8168 16436 8174 16448
rect 11238 16436 11244 16448
rect 8168 16408 11244 16436
rect 8168 16396 8174 16408
rect 11238 16396 11244 16408
rect 11296 16396 11302 16448
rect 11624 16436 11652 16680
rect 13538 16668 13544 16680
rect 13596 16668 13602 16720
rect 14182 16668 14188 16720
rect 14240 16708 14246 16720
rect 16482 16708 16488 16720
rect 14240 16680 16488 16708
rect 14240 16668 14246 16680
rect 16482 16668 16488 16680
rect 16540 16708 16546 16720
rect 16540 16680 17448 16708
rect 16540 16668 16546 16680
rect 11974 16600 11980 16652
rect 12032 16640 12038 16652
rect 13173 16643 13231 16649
rect 13173 16640 13185 16643
rect 12032 16612 13185 16640
rect 12032 16600 12038 16612
rect 13173 16609 13185 16612
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 13280 16612 13492 16640
rect 12066 16532 12072 16584
rect 12124 16572 12130 16584
rect 13280 16572 13308 16612
rect 12124 16544 13308 16572
rect 13357 16575 13415 16581
rect 12124 16532 12130 16544
rect 13357 16541 13369 16575
rect 13403 16541 13415 16575
rect 13464 16572 13492 16612
rect 13814 16600 13820 16652
rect 13872 16640 13878 16652
rect 14734 16640 14740 16652
rect 13872 16612 14740 16640
rect 13872 16600 13878 16612
rect 14734 16600 14740 16612
rect 14792 16600 14798 16652
rect 15562 16600 15568 16652
rect 15620 16640 15626 16652
rect 16025 16643 16083 16649
rect 16025 16640 16037 16643
rect 15620 16612 16037 16640
rect 15620 16600 15626 16612
rect 16025 16609 16037 16612
rect 16071 16609 16083 16643
rect 16025 16603 16083 16609
rect 16292 16643 16350 16649
rect 16292 16609 16304 16643
rect 16338 16640 16350 16643
rect 17126 16640 17132 16652
rect 16338 16612 17132 16640
rect 16338 16609 16350 16612
rect 16292 16603 16350 16609
rect 17126 16600 17132 16612
rect 17184 16600 17190 16652
rect 15286 16572 15292 16584
rect 13464 16544 15292 16572
rect 13357 16535 13415 16541
rect 12250 16464 12256 16516
rect 12308 16504 12314 16516
rect 13372 16504 13400 16535
rect 15286 16532 15292 16544
rect 15344 16532 15350 16584
rect 12308 16476 13400 16504
rect 12308 16464 12314 16476
rect 14826 16464 14832 16516
rect 14884 16504 14890 16516
rect 15838 16504 15844 16516
rect 14884 16476 15844 16504
rect 14884 16464 14890 16476
rect 15838 16464 15844 16476
rect 15896 16464 15902 16516
rect 17420 16513 17448 16680
rect 17678 16668 17684 16720
rect 17736 16708 17742 16720
rect 19245 16711 19303 16717
rect 19245 16708 19257 16711
rect 17736 16680 19257 16708
rect 17736 16668 17742 16680
rect 19245 16677 19257 16680
rect 19291 16677 19303 16711
rect 19245 16671 19303 16677
rect 19150 16532 19156 16584
rect 19208 16572 19214 16584
rect 19337 16575 19395 16581
rect 19337 16572 19349 16575
rect 19208 16544 19349 16572
rect 19208 16532 19214 16544
rect 19337 16541 19349 16544
rect 19383 16541 19395 16575
rect 19337 16535 19395 16541
rect 17405 16507 17463 16513
rect 17405 16473 17417 16507
rect 17451 16473 17463 16507
rect 17405 16467 17463 16473
rect 12434 16436 12440 16448
rect 11624 16408 12440 16436
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 3050 16232 3056 16244
rect 3011 16204 3056 16232
rect 3050 16192 3056 16204
rect 3108 16192 3114 16244
rect 7558 16192 7564 16244
rect 7616 16232 7622 16244
rect 8570 16232 8576 16244
rect 7616 16204 8576 16232
rect 7616 16192 7622 16204
rect 8570 16192 8576 16204
rect 8628 16192 8634 16244
rect 10413 16235 10471 16241
rect 10413 16201 10425 16235
rect 10459 16232 10471 16235
rect 11882 16232 11888 16244
rect 10459 16204 11888 16232
rect 10459 16201 10471 16204
rect 10413 16195 10471 16201
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 9582 16164 9588 16176
rect 9495 16136 9588 16164
rect 9582 16124 9588 16136
rect 9640 16164 9646 16176
rect 10226 16164 10232 16176
rect 9640 16136 10232 16164
rect 9640 16124 9646 16136
rect 10226 16124 10232 16136
rect 10284 16164 10290 16176
rect 10284 16136 11008 16164
rect 10284 16124 10290 16136
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 3896 16068 5181 16096
rect 1673 16031 1731 16037
rect 1673 15997 1685 16031
rect 1719 16028 1731 16031
rect 3326 16028 3332 16040
rect 1719 16000 3332 16028
rect 1719 15997 1731 16000
rect 1673 15991 1731 15997
rect 3326 15988 3332 16000
rect 3384 15988 3390 16040
rect 3896 15972 3924 16068
rect 5169 16065 5181 16068
rect 5215 16065 5227 16099
rect 5169 16059 5227 16065
rect 10318 16056 10324 16108
rect 10376 16096 10382 16108
rect 10980 16105 11008 16136
rect 10873 16099 10931 16105
rect 10873 16096 10885 16099
rect 10376 16068 10885 16096
rect 10376 16056 10382 16068
rect 10873 16065 10885 16068
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 10965 16099 11023 16105
rect 10965 16065 10977 16099
rect 11011 16065 11023 16099
rect 10965 16059 11023 16065
rect 15562 16056 15568 16108
rect 15620 16096 15626 16108
rect 15746 16096 15752 16108
rect 15620 16068 15752 16096
rect 15620 16056 15626 16068
rect 15746 16056 15752 16068
rect 15804 16056 15810 16108
rect 19518 16056 19524 16108
rect 19576 16096 19582 16108
rect 20530 16096 20536 16108
rect 19576 16068 20536 16096
rect 19576 16056 19582 16068
rect 20530 16056 20536 16068
rect 20588 16056 20594 16108
rect 4985 16031 5043 16037
rect 4985 15997 4997 16031
rect 5031 16028 5043 16031
rect 5350 16028 5356 16040
rect 5031 16000 5356 16028
rect 5031 15997 5043 16000
rect 4985 15991 5043 15997
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 16028 6975 16031
rect 8110 16028 8116 16040
rect 6963 16000 8116 16028
rect 6963 15997 6975 16000
rect 6917 15991 6975 15997
rect 8110 15988 8116 16000
rect 8168 15988 8174 16040
rect 8205 16031 8263 16037
rect 8205 15997 8217 16031
rect 8251 16028 8263 16031
rect 8294 16028 8300 16040
rect 8251 16000 8300 16028
rect 8251 15997 8263 16000
rect 8205 15991 8263 15997
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 8472 16031 8530 16037
rect 8472 15997 8484 16031
rect 8518 16028 8530 16031
rect 10686 16028 10692 16040
rect 8518 16000 10692 16028
rect 8518 15997 8530 16000
rect 8472 15991 8530 15997
rect 10686 15988 10692 16000
rect 10744 15988 10750 16040
rect 12618 15988 12624 16040
rect 12676 16028 12682 16040
rect 13357 16031 13415 16037
rect 13357 16028 13369 16031
rect 12676 16000 13369 16028
rect 12676 15988 12682 16000
rect 13357 15997 13369 16000
rect 13403 15997 13415 16031
rect 13357 15991 13415 15997
rect 13624 16031 13682 16037
rect 13624 15997 13636 16031
rect 13670 16028 13682 16031
rect 14090 16028 14096 16040
rect 13670 16000 14096 16028
rect 13670 15997 13682 16000
rect 13624 15991 13682 15997
rect 1940 15963 1998 15969
rect 1940 15929 1952 15963
rect 1986 15960 1998 15963
rect 3878 15960 3884 15972
rect 1986 15932 3884 15960
rect 1986 15929 1998 15932
rect 1940 15923 1998 15929
rect 3878 15920 3884 15932
rect 3936 15920 3942 15972
rect 4062 15920 4068 15972
rect 4120 15960 4126 15972
rect 5077 15963 5135 15969
rect 4120 15932 5028 15960
rect 4120 15920 4126 15932
rect 1578 15852 1584 15904
rect 1636 15892 1642 15904
rect 2314 15892 2320 15904
rect 1636 15864 2320 15892
rect 1636 15852 1642 15864
rect 2314 15852 2320 15864
rect 2372 15852 2378 15904
rect 4614 15892 4620 15904
rect 4575 15864 4620 15892
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 5000 15892 5028 15932
rect 5077 15929 5089 15963
rect 5123 15960 5135 15963
rect 5534 15960 5540 15972
rect 5123 15932 5540 15960
rect 5123 15929 5135 15932
rect 5077 15923 5135 15929
rect 5534 15920 5540 15932
rect 5592 15920 5598 15972
rect 7193 15963 7251 15969
rect 7193 15929 7205 15963
rect 7239 15960 7251 15963
rect 7558 15960 7564 15972
rect 7239 15932 7564 15960
rect 7239 15929 7251 15932
rect 7193 15923 7251 15929
rect 7558 15920 7564 15932
rect 7616 15920 7622 15972
rect 10410 15920 10416 15972
rect 10468 15960 10474 15972
rect 10781 15963 10839 15969
rect 10781 15960 10793 15963
rect 10468 15932 10793 15960
rect 10468 15920 10474 15932
rect 10781 15929 10793 15932
rect 10827 15929 10839 15963
rect 10781 15923 10839 15929
rect 10870 15920 10876 15972
rect 10928 15960 10934 15972
rect 12066 15960 12072 15972
rect 10928 15932 12072 15960
rect 10928 15920 10934 15932
rect 12066 15920 12072 15932
rect 12124 15920 12130 15972
rect 13372 15960 13400 15991
rect 14090 15988 14096 16000
rect 14148 15988 14154 16040
rect 15764 16028 15792 16056
rect 18782 16037 18788 16040
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 15764 16000 18521 16028
rect 18509 15997 18521 16000
rect 18555 15997 18567 16031
rect 18776 16028 18788 16037
rect 18743 16000 18788 16028
rect 18509 15991 18567 15997
rect 18776 15991 18788 16000
rect 18782 15988 18788 15991
rect 18840 15988 18846 16040
rect 13998 15960 14004 15972
rect 13372 15932 14004 15960
rect 13998 15920 14004 15932
rect 14056 15920 14062 15972
rect 16016 15963 16074 15969
rect 14476 15932 15976 15960
rect 14476 15892 14504 15932
rect 15948 15904 15976 15932
rect 16016 15929 16028 15963
rect 16062 15960 16074 15963
rect 16390 15960 16396 15972
rect 16062 15932 16396 15960
rect 16062 15929 16074 15932
rect 16016 15923 16074 15929
rect 16390 15920 16396 15932
rect 16448 15920 16454 15972
rect 19334 15960 19340 15972
rect 19076 15932 19340 15960
rect 5000 15864 14504 15892
rect 14550 15852 14556 15904
rect 14608 15892 14614 15904
rect 14737 15895 14795 15901
rect 14737 15892 14749 15895
rect 14608 15864 14749 15892
rect 14608 15852 14614 15864
rect 14737 15861 14749 15864
rect 14783 15892 14795 15895
rect 15194 15892 15200 15904
rect 14783 15864 15200 15892
rect 14783 15861 14795 15864
rect 14737 15855 14795 15861
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 15930 15852 15936 15904
rect 15988 15852 15994 15904
rect 17126 15892 17132 15904
rect 17087 15864 17132 15892
rect 17126 15852 17132 15864
rect 17184 15852 17190 15904
rect 18782 15852 18788 15904
rect 18840 15892 18846 15904
rect 19076 15892 19104 15932
rect 19334 15920 19340 15932
rect 19392 15920 19398 15972
rect 18840 15864 19104 15892
rect 18840 15852 18846 15864
rect 19150 15852 19156 15904
rect 19208 15892 19214 15904
rect 19889 15895 19947 15901
rect 19889 15892 19901 15895
rect 19208 15864 19901 15892
rect 19208 15852 19214 15864
rect 19889 15861 19901 15864
rect 19935 15861 19947 15895
rect 19889 15855 19947 15861
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 2869 15691 2927 15697
rect 2869 15657 2881 15691
rect 2915 15688 2927 15691
rect 4614 15688 4620 15700
rect 2915 15660 4620 15688
rect 2915 15657 2927 15660
rect 2869 15651 2927 15657
rect 4614 15648 4620 15660
rect 4672 15648 4678 15700
rect 8294 15688 8300 15700
rect 6472 15660 8300 15688
rect 1397 15623 1455 15629
rect 1397 15589 1409 15623
rect 1443 15620 1455 15623
rect 1765 15623 1823 15629
rect 1765 15620 1777 15623
rect 1443 15592 1777 15620
rect 1443 15589 1455 15592
rect 1397 15583 1455 15589
rect 1765 15589 1777 15592
rect 1811 15620 1823 15623
rect 1811 15592 6408 15620
rect 1811 15589 1823 15592
rect 1765 15583 1823 15589
rect 2774 15512 2780 15564
rect 2832 15552 2838 15564
rect 2832 15524 2877 15552
rect 2832 15512 2838 15524
rect 3326 15512 3332 15564
rect 3384 15552 3390 15564
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 3384 15524 4077 15552
rect 3384 15512 3390 15524
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 4332 15555 4390 15561
rect 4332 15521 4344 15555
rect 4378 15552 4390 15555
rect 5442 15552 5448 15564
rect 4378 15524 5448 15552
rect 4378 15521 4390 15524
rect 4332 15515 4390 15521
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 3050 15484 3056 15496
rect 3011 15456 3056 15484
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 6380 15484 6408 15592
rect 6472 15561 6500 15660
rect 8294 15648 8300 15660
rect 8352 15688 8358 15700
rect 8665 15691 8723 15697
rect 8665 15688 8677 15691
rect 8352 15660 8677 15688
rect 8352 15648 8358 15660
rect 8665 15657 8677 15660
rect 8711 15688 8723 15691
rect 8846 15688 8852 15700
rect 8711 15660 8852 15688
rect 8711 15657 8723 15660
rect 8665 15651 8723 15657
rect 8846 15648 8852 15660
rect 8904 15688 8910 15700
rect 9490 15688 9496 15700
rect 8904 15660 9496 15688
rect 8904 15648 8910 15660
rect 9490 15648 9496 15660
rect 9548 15648 9554 15700
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 10045 15691 10103 15697
rect 9732 15660 9777 15688
rect 9732 15648 9738 15660
rect 10045 15657 10057 15691
rect 10091 15688 10103 15691
rect 11241 15691 11299 15697
rect 11241 15688 11253 15691
rect 10091 15660 11253 15688
rect 10091 15657 10103 15660
rect 10045 15651 10103 15657
rect 11241 15657 11253 15660
rect 11287 15657 11299 15691
rect 11241 15651 11299 15657
rect 11701 15691 11759 15697
rect 11701 15657 11713 15691
rect 11747 15688 11759 15691
rect 12434 15688 12440 15700
rect 11747 15660 12440 15688
rect 11747 15657 11759 15660
rect 11701 15651 11759 15657
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 13998 15648 14004 15700
rect 14056 15688 14062 15700
rect 14366 15688 14372 15700
rect 14056 15660 14372 15688
rect 14056 15648 14062 15660
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 15286 15648 15292 15700
rect 15344 15688 15350 15700
rect 19705 15691 19763 15697
rect 19705 15688 19717 15691
rect 15344 15660 19717 15688
rect 15344 15648 15350 15660
rect 19705 15657 19717 15660
rect 19751 15657 19763 15691
rect 19705 15651 19763 15657
rect 6724 15623 6782 15629
rect 6724 15589 6736 15623
rect 6770 15620 6782 15623
rect 6822 15620 6828 15632
rect 6770 15592 6828 15620
rect 6770 15589 6782 15592
rect 6724 15583 6782 15589
rect 6822 15580 6828 15592
rect 6880 15580 6886 15632
rect 10778 15620 10784 15632
rect 6932 15592 10784 15620
rect 6457 15555 6515 15561
rect 6457 15521 6469 15555
rect 6503 15521 6515 15555
rect 6932 15552 6960 15592
rect 10778 15580 10784 15592
rect 10836 15580 10842 15632
rect 11146 15580 11152 15632
rect 11204 15620 11210 15632
rect 11882 15620 11888 15632
rect 11204 15592 11888 15620
rect 11204 15580 11210 15592
rect 11882 15580 11888 15592
rect 11940 15620 11946 15632
rect 13265 15623 13323 15629
rect 13265 15620 13277 15623
rect 11940 15592 13277 15620
rect 11940 15580 11946 15592
rect 13265 15589 13277 15592
rect 13311 15589 13323 15623
rect 18046 15620 18052 15632
rect 13265 15583 13323 15589
rect 13372 15592 18052 15620
rect 6457 15515 6515 15521
rect 6564 15524 6960 15552
rect 6564 15484 6592 15524
rect 7098 15512 7104 15564
rect 7156 15552 7162 15564
rect 8849 15555 8907 15561
rect 8849 15552 8861 15555
rect 7156 15524 8861 15552
rect 7156 15512 7162 15524
rect 8849 15521 8861 15524
rect 8895 15521 8907 15555
rect 8849 15515 8907 15521
rect 8938 15512 8944 15564
rect 8996 15552 9002 15564
rect 11514 15552 11520 15564
rect 8996 15524 11520 15552
rect 8996 15512 9002 15524
rect 11514 15512 11520 15524
rect 11572 15512 11578 15564
rect 11609 15555 11667 15561
rect 11609 15521 11621 15555
rect 11655 15552 11667 15555
rect 12066 15552 12072 15564
rect 11655 15524 12072 15552
rect 11655 15521 11667 15524
rect 11609 15515 11667 15521
rect 12066 15512 12072 15524
rect 12124 15512 12130 15564
rect 13078 15512 13084 15564
rect 13136 15552 13142 15564
rect 13173 15555 13231 15561
rect 13173 15552 13185 15555
rect 13136 15524 13185 15552
rect 13136 15512 13142 15524
rect 13173 15521 13185 15524
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 10134 15484 10140 15496
rect 6380 15456 6592 15484
rect 10095 15456 10140 15484
rect 10134 15444 10140 15456
rect 10192 15444 10198 15496
rect 10318 15484 10324 15496
rect 10279 15456 10324 15484
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 10686 15444 10692 15496
rect 10744 15484 10750 15496
rect 11793 15487 11851 15493
rect 11793 15484 11805 15487
rect 10744 15456 11805 15484
rect 10744 15444 10750 15456
rect 11793 15453 11805 15456
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 13372 15484 13400 15592
rect 18046 15580 18052 15592
rect 18104 15580 18110 15632
rect 14553 15555 14611 15561
rect 14553 15521 14565 15555
rect 14599 15552 14611 15555
rect 15562 15552 15568 15564
rect 14599 15524 15568 15552
rect 14599 15521 14611 15524
rect 14553 15515 14611 15521
rect 15562 15512 15568 15524
rect 15620 15512 15626 15564
rect 16476 15555 16534 15561
rect 16476 15521 16488 15555
rect 16522 15552 16534 15555
rect 17678 15552 17684 15564
rect 16522 15524 17684 15552
rect 16522 15521 16534 15524
rect 16476 15515 16534 15521
rect 17678 15512 17684 15524
rect 17736 15512 17742 15564
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 19613 15555 19671 15561
rect 19613 15552 19625 15555
rect 19392 15524 19625 15552
rect 19392 15512 19398 15524
rect 19613 15521 19625 15524
rect 19659 15521 19671 15555
rect 19613 15515 19671 15521
rect 12216 15456 13400 15484
rect 13449 15487 13507 15493
rect 12216 15444 12222 15456
rect 13449 15453 13461 15487
rect 13495 15484 13507 15487
rect 13538 15484 13544 15496
rect 13495 15456 13544 15484
rect 13495 15453 13507 15456
rect 13449 15447 13507 15453
rect 7466 15376 7472 15428
rect 7524 15416 7530 15428
rect 7837 15419 7895 15425
rect 7837 15416 7849 15419
rect 7524 15388 7849 15416
rect 7524 15376 7530 15388
rect 7837 15385 7849 15388
rect 7883 15416 7895 15419
rect 13464 15416 13492 15447
rect 13538 15444 13544 15456
rect 13596 15444 13602 15496
rect 14366 15444 14372 15496
rect 14424 15484 14430 15496
rect 16209 15487 16267 15493
rect 16209 15484 16221 15487
rect 14424 15456 16221 15484
rect 14424 15444 14430 15456
rect 16209 15453 16221 15456
rect 16255 15453 16267 15487
rect 16209 15447 16267 15453
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15484 19947 15487
rect 20254 15484 20260 15496
rect 19935 15456 20260 15484
rect 19935 15453 19947 15456
rect 19889 15447 19947 15453
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 7883 15388 13492 15416
rect 7883 15385 7895 15388
rect 7837 15379 7895 15385
rect 1946 15308 1952 15360
rect 2004 15348 2010 15360
rect 2409 15351 2467 15357
rect 2409 15348 2421 15351
rect 2004 15320 2421 15348
rect 2004 15308 2010 15320
rect 2409 15317 2421 15320
rect 2455 15317 2467 15351
rect 2409 15311 2467 15317
rect 3878 15308 3884 15360
rect 3936 15348 3942 15360
rect 5445 15351 5503 15357
rect 5445 15348 5457 15351
rect 3936 15320 5457 15348
rect 3936 15308 3942 15320
rect 5445 15317 5457 15320
rect 5491 15317 5503 15351
rect 5445 15311 5503 15317
rect 6178 15308 6184 15360
rect 6236 15348 6242 15360
rect 9306 15348 9312 15360
rect 6236 15320 9312 15348
rect 6236 15308 6242 15320
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 12805 15351 12863 15357
rect 12805 15348 12817 15351
rect 11112 15320 12817 15348
rect 11112 15308 11118 15320
rect 12805 15317 12817 15320
rect 12851 15317 12863 15351
rect 12805 15311 12863 15317
rect 16390 15308 16396 15360
rect 16448 15348 16454 15360
rect 17589 15351 17647 15357
rect 17589 15348 17601 15351
rect 16448 15320 17601 15348
rect 16448 15308 16454 15320
rect 17589 15317 17601 15320
rect 17635 15317 17647 15351
rect 17589 15311 17647 15317
rect 19245 15351 19303 15357
rect 19245 15317 19257 15351
rect 19291 15348 19303 15351
rect 19610 15348 19616 15360
rect 19291 15320 19616 15348
rect 19291 15317 19303 15320
rect 19245 15311 19303 15317
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 2774 15104 2780 15156
rect 2832 15144 2838 15156
rect 3329 15147 3387 15153
rect 3329 15144 3341 15147
rect 2832 15116 3341 15144
rect 2832 15104 2838 15116
rect 3329 15113 3341 15116
rect 3375 15113 3387 15147
rect 3329 15107 3387 15113
rect 6086 15104 6092 15156
rect 6144 15144 6150 15156
rect 6457 15147 6515 15153
rect 6457 15144 6469 15147
rect 6144 15116 6469 15144
rect 6144 15104 6150 15116
rect 6457 15113 6469 15116
rect 6503 15144 6515 15147
rect 6546 15144 6552 15156
rect 6503 15116 6552 15144
rect 6503 15113 6515 15116
rect 6457 15107 6515 15113
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 14737 15147 14795 15153
rect 14737 15144 14749 15147
rect 8772 15116 14749 15144
rect 7742 15076 7748 15088
rect 2424 15048 7748 15076
rect 2424 15017 2452 15048
rect 7742 15036 7748 15048
rect 7800 15036 7806 15088
rect 2409 15011 2467 15017
rect 2409 14977 2421 15011
rect 2455 14977 2467 15011
rect 3878 15008 3884 15020
rect 3839 14980 3884 15008
rect 2409 14971 2467 14977
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 5442 15008 5448 15020
rect 5403 14980 5448 15008
rect 5442 14968 5448 14980
rect 5500 14968 5506 15020
rect 7374 15008 7380 15020
rect 7335 14980 7380 15008
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 2133 14943 2191 14949
rect 2133 14909 2145 14943
rect 2179 14940 2191 14943
rect 6546 14940 6552 14952
rect 2179 14912 6552 14940
rect 2179 14909 2191 14912
rect 2133 14903 2191 14909
rect 6546 14900 6552 14912
rect 6604 14900 6610 14952
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14940 6699 14943
rect 7098 14940 7104 14952
rect 6687 14912 7104 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 7098 14900 7104 14912
rect 7156 14900 7162 14952
rect 7285 14943 7343 14949
rect 7285 14909 7297 14943
rect 7331 14940 7343 14943
rect 8772 14940 8800 15116
rect 14737 15113 14749 15116
rect 14783 15113 14795 15147
rect 16298 15144 16304 15156
rect 16259 15116 16304 15144
rect 14737 15107 14795 15113
rect 16298 15104 16304 15116
rect 16356 15104 16362 15156
rect 10321 15079 10379 15085
rect 10321 15045 10333 15079
rect 10367 15076 10379 15079
rect 11146 15076 11152 15088
rect 10367 15048 11152 15076
rect 10367 15045 10379 15048
rect 10321 15039 10379 15045
rect 11146 15036 11152 15048
rect 11204 15076 11210 15088
rect 12250 15076 12256 15088
rect 11204 15048 12256 15076
rect 11204 15036 11210 15048
rect 12250 15036 12256 15048
rect 12308 15036 12314 15088
rect 13909 15079 13967 15085
rect 13909 15045 13921 15079
rect 13955 15076 13967 15079
rect 14090 15076 14096 15088
rect 13955 15048 14096 15076
rect 13955 15045 13967 15048
rect 13909 15039 13967 15045
rect 14090 15036 14096 15048
rect 14148 15036 14154 15088
rect 14366 15036 14372 15088
rect 14424 15076 14430 15088
rect 18782 15076 18788 15088
rect 14424 15048 18788 15076
rect 14424 15036 14430 15048
rect 18782 15036 18788 15048
rect 18840 15036 18846 15088
rect 8846 14968 8852 15020
rect 8904 15008 8910 15020
rect 8941 15011 8999 15017
rect 8941 15008 8953 15011
rect 8904 14980 8953 15008
rect 8904 14968 8910 14980
rect 8941 14977 8953 14980
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 10686 14968 10692 15020
rect 10744 15008 10750 15020
rect 10744 14980 11376 15008
rect 10744 14968 10750 14980
rect 7331 14912 8800 14940
rect 9208 14943 9266 14949
rect 7331 14909 7343 14912
rect 7285 14903 7343 14909
rect 9208 14909 9220 14943
rect 9254 14940 9266 14943
rect 9582 14940 9588 14952
rect 9254 14912 9588 14940
rect 9254 14909 9266 14912
rect 9208 14903 9266 14909
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 11238 14940 11244 14952
rect 11199 14912 11244 14940
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 11348 14940 11376 14980
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 12529 15011 12587 15017
rect 12529 15008 12541 15011
rect 12492 14980 12541 15008
rect 12492 14968 12498 14980
rect 12529 14977 12541 14980
rect 12575 14977 12587 15011
rect 12529 14971 12587 14977
rect 13538 14968 13544 15020
rect 13596 15008 13602 15020
rect 15289 15011 15347 15017
rect 15289 15008 15301 15011
rect 13596 14980 15301 15008
rect 13596 14968 13602 14980
rect 15289 14977 15301 14980
rect 15335 14977 15347 15011
rect 15289 14971 15347 14977
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 15197 14943 15255 14949
rect 15197 14940 15209 14943
rect 11348 14912 15209 14940
rect 15197 14909 15209 14912
rect 15243 14909 15255 14943
rect 16868 14940 16896 14971
rect 15197 14903 15255 14909
rect 15304 14912 16896 14940
rect 2225 14875 2283 14881
rect 2225 14841 2237 14875
rect 2271 14872 2283 14875
rect 7193 14875 7251 14881
rect 2271 14844 6868 14872
rect 2271 14841 2283 14844
rect 2225 14835 2283 14841
rect 1765 14807 1823 14813
rect 1765 14773 1777 14807
rect 1811 14804 1823 14807
rect 2314 14804 2320 14816
rect 1811 14776 2320 14804
rect 1811 14773 1823 14776
rect 1765 14767 1823 14773
rect 2314 14764 2320 14776
rect 2372 14764 2378 14816
rect 3694 14804 3700 14816
rect 3655 14776 3700 14804
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 3789 14807 3847 14813
rect 3789 14773 3801 14807
rect 3835 14804 3847 14807
rect 4893 14807 4951 14813
rect 4893 14804 4905 14807
rect 3835 14776 4905 14804
rect 3835 14773 3847 14776
rect 3789 14767 3847 14773
rect 4893 14773 4905 14776
rect 4939 14773 4951 14807
rect 4893 14767 4951 14773
rect 4982 14764 4988 14816
rect 5040 14804 5046 14816
rect 5261 14807 5319 14813
rect 5261 14804 5273 14807
rect 5040 14776 5273 14804
rect 5040 14764 5046 14776
rect 5261 14773 5273 14776
rect 5307 14773 5319 14807
rect 5261 14767 5319 14773
rect 5353 14807 5411 14813
rect 5353 14773 5365 14807
rect 5399 14804 5411 14807
rect 5534 14804 5540 14816
rect 5399 14776 5540 14804
rect 5399 14773 5411 14776
rect 5353 14767 5411 14773
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 6840 14813 6868 14844
rect 7193 14841 7205 14875
rect 7239 14872 7251 14875
rect 11054 14872 11060 14884
rect 7239 14844 11060 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 11054 14832 11060 14844
rect 11112 14832 11118 14884
rect 12796 14875 12854 14881
rect 12796 14841 12808 14875
rect 12842 14872 12854 14875
rect 12842 14844 12940 14872
rect 12842 14841 12854 14844
rect 12796 14835 12854 14841
rect 6825 14807 6883 14813
rect 6825 14773 6837 14807
rect 6871 14773 6883 14807
rect 6825 14767 6883 14773
rect 8386 14764 8392 14816
rect 8444 14804 8450 14816
rect 11330 14804 11336 14816
rect 8444 14776 11336 14804
rect 8444 14764 8450 14776
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 11425 14807 11483 14813
rect 11425 14773 11437 14807
rect 11471 14804 11483 14807
rect 12434 14804 12440 14816
rect 11471 14776 12440 14804
rect 11471 14773 11483 14776
rect 11425 14767 11483 14773
rect 12434 14764 12440 14776
rect 12492 14764 12498 14816
rect 12912 14804 12940 14844
rect 13170 14832 13176 14884
rect 13228 14872 13234 14884
rect 15105 14875 15163 14881
rect 15105 14872 15117 14875
rect 13228 14844 15117 14872
rect 13228 14832 13234 14844
rect 15105 14841 15117 14844
rect 15151 14841 15163 14875
rect 15105 14835 15163 14841
rect 13446 14804 13452 14816
rect 12912 14776 13452 14804
rect 13446 14764 13452 14776
rect 13504 14804 13510 14816
rect 15304 14804 15332 14912
rect 18782 14900 18788 14952
rect 18840 14940 18846 14952
rect 19150 14949 19156 14952
rect 18877 14943 18935 14949
rect 18877 14940 18889 14943
rect 18840 14912 18889 14940
rect 18840 14900 18846 14912
rect 18877 14909 18889 14912
rect 18923 14909 18935 14943
rect 18877 14903 18935 14909
rect 19144 14903 19156 14949
rect 19208 14940 19214 14952
rect 19208 14912 19244 14940
rect 19150 14900 19156 14903
rect 19208 14900 19214 14912
rect 16669 14875 16727 14881
rect 16669 14841 16681 14875
rect 16715 14872 16727 14875
rect 16942 14872 16948 14884
rect 16715 14844 16948 14872
rect 16715 14841 16727 14844
rect 16669 14835 16727 14841
rect 16942 14832 16948 14844
rect 17000 14832 17006 14884
rect 13504 14776 15332 14804
rect 16761 14807 16819 14813
rect 13504 14764 13510 14776
rect 16761 14773 16773 14807
rect 16807 14804 16819 14807
rect 17310 14804 17316 14816
rect 16807 14776 17316 14804
rect 16807 14773 16819 14776
rect 16761 14767 16819 14773
rect 17310 14764 17316 14776
rect 17368 14764 17374 14816
rect 20254 14804 20260 14816
rect 20215 14776 20260 14804
rect 20254 14764 20260 14776
rect 20312 14764 20318 14816
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 2866 14600 2872 14612
rect 2827 14572 2872 14600
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 3694 14560 3700 14612
rect 3752 14600 3758 14612
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 3752 14572 4077 14600
rect 3752 14560 3758 14572
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 4065 14563 4123 14569
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 13998 14600 14004 14612
rect 6604 14572 14004 14600
rect 6604 14560 6610 14572
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 14277 14603 14335 14609
rect 14277 14569 14289 14603
rect 14323 14600 14335 14603
rect 14366 14600 14372 14612
rect 14323 14572 14372 14600
rect 14323 14569 14335 14572
rect 14277 14563 14335 14569
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 15289 14603 15347 14609
rect 15289 14569 15301 14603
rect 15335 14600 15347 14603
rect 19334 14600 19340 14612
rect 15335 14572 19340 14600
rect 15335 14569 15347 14572
rect 15289 14563 15347 14569
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 19610 14600 19616 14612
rect 19571 14572 19616 14600
rect 19610 14560 19616 14572
rect 19668 14560 19674 14612
rect 6356 14535 6414 14541
rect 6356 14501 6368 14535
rect 6402 14532 6414 14535
rect 7466 14532 7472 14544
rect 6402 14504 7472 14532
rect 6402 14501 6414 14504
rect 6356 14495 6414 14501
rect 7466 14492 7472 14504
rect 7524 14492 7530 14544
rect 9030 14492 9036 14544
rect 9088 14532 9094 14544
rect 12710 14532 12716 14544
rect 9088 14504 12716 14532
rect 9088 14492 9094 14504
rect 12710 14492 12716 14504
rect 12768 14492 12774 14544
rect 15562 14492 15568 14544
rect 15620 14532 15626 14544
rect 15620 14504 18736 14532
rect 15620 14492 15626 14504
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 2832 14436 2877 14464
rect 2832 14424 2838 14436
rect 3786 14424 3792 14476
rect 3844 14464 3850 14476
rect 4433 14467 4491 14473
rect 4433 14464 4445 14467
rect 3844 14436 4445 14464
rect 3844 14424 3850 14436
rect 4433 14433 4445 14436
rect 4479 14433 4491 14467
rect 4433 14427 4491 14433
rect 4525 14467 4583 14473
rect 4525 14433 4537 14467
rect 4571 14464 4583 14467
rect 5442 14464 5448 14476
rect 4571 14436 5448 14464
rect 4571 14433 4583 14436
rect 4525 14427 4583 14433
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 6086 14464 6092 14476
rect 6047 14436 6092 14464
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 8297 14467 8355 14473
rect 8297 14433 8309 14467
rect 8343 14433 8355 14467
rect 8297 14427 8355 14433
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14396 1455 14399
rect 2682 14396 2688 14408
rect 1443 14368 2688 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14396 3111 14399
rect 3418 14396 3424 14408
rect 3099 14368 3424 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 3418 14356 3424 14368
rect 3476 14356 3482 14408
rect 4709 14399 4767 14405
rect 4709 14365 4721 14399
rect 4755 14396 4767 14399
rect 4890 14396 4896 14408
rect 4755 14368 4896 14396
rect 4755 14365 4767 14368
rect 4709 14359 4767 14365
rect 4890 14356 4896 14368
rect 4948 14396 4954 14408
rect 5350 14396 5356 14408
rect 4948 14368 5356 14396
rect 4948 14356 4954 14368
rect 5350 14356 5356 14368
rect 5408 14356 5414 14408
rect 2498 14288 2504 14340
rect 2556 14328 2562 14340
rect 3694 14328 3700 14340
rect 2556 14300 3700 14328
rect 2556 14288 2562 14300
rect 3694 14288 3700 14300
rect 3752 14328 3758 14340
rect 4982 14328 4988 14340
rect 3752 14300 4988 14328
rect 3752 14288 3758 14300
rect 4982 14288 4988 14300
rect 5040 14288 5046 14340
rect 8312 14328 8340 14427
rect 9490 14424 9496 14476
rect 9548 14464 9554 14476
rect 9674 14464 9680 14476
rect 9548 14436 9680 14464
rect 9548 14424 9554 14436
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 9944 14467 10002 14473
rect 9944 14433 9956 14467
rect 9990 14464 10002 14467
rect 11146 14464 11152 14476
rect 9990 14436 11152 14464
rect 9990 14433 10002 14436
rect 9944 14427 10002 14433
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 12152 14467 12210 14473
rect 12152 14433 12164 14467
rect 12198 14464 12210 14467
rect 12434 14464 12440 14476
rect 12198 14436 12440 14464
rect 12198 14433 12210 14436
rect 12152 14427 12210 14433
rect 12434 14424 12440 14436
rect 12492 14464 12498 14476
rect 13354 14464 13360 14476
rect 12492 14436 13360 14464
rect 12492 14424 12498 14436
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 14090 14464 14096 14476
rect 14051 14436 14096 14464
rect 14090 14424 14096 14436
rect 14148 14424 14154 14476
rect 15746 14424 15752 14476
rect 15804 14464 15810 14476
rect 16301 14467 16359 14473
rect 16301 14464 16313 14467
rect 15804 14436 16313 14464
rect 15804 14424 15810 14436
rect 16301 14433 16313 14436
rect 16347 14433 16359 14467
rect 16301 14427 16359 14433
rect 16568 14467 16626 14473
rect 16568 14433 16580 14467
rect 16614 14464 16626 14467
rect 17034 14464 17040 14476
rect 16614 14436 17040 14464
rect 16614 14433 16626 14436
rect 16568 14427 16626 14433
rect 17034 14424 17040 14436
rect 17092 14424 17098 14476
rect 18708 14473 18736 14504
rect 18693 14467 18751 14473
rect 18693 14433 18705 14467
rect 18739 14433 18751 14467
rect 18693 14427 18751 14433
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14396 8631 14399
rect 8846 14396 8852 14408
rect 8619 14368 8852 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 8846 14356 8852 14368
rect 8904 14356 8910 14408
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 11606 14396 11612 14408
rect 11112 14368 11612 14396
rect 11112 14356 11118 14368
rect 11606 14356 11612 14368
rect 11664 14396 11670 14408
rect 11885 14399 11943 14405
rect 11885 14396 11897 14399
rect 11664 14368 11897 14396
rect 11664 14356 11670 14368
rect 11885 14365 11897 14368
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 14550 14396 14556 14408
rect 14424 14368 14556 14396
rect 14424 14356 14430 14368
rect 14550 14356 14556 14368
rect 14608 14356 14614 14408
rect 19702 14396 19708 14408
rect 19663 14368 19708 14396
rect 19702 14356 19708 14368
rect 19760 14356 19766 14408
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14396 19947 14399
rect 20162 14396 20168 14408
rect 19935 14368 20168 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 20162 14356 20168 14368
rect 20220 14356 20226 14408
rect 9490 14328 9496 14340
rect 8312 14300 9496 14328
rect 9490 14288 9496 14300
rect 9548 14288 9554 14340
rect 13265 14331 13323 14337
rect 10612 14300 11376 14328
rect 2409 14263 2467 14269
rect 2409 14229 2421 14263
rect 2455 14260 2467 14263
rect 5994 14260 6000 14272
rect 2455 14232 6000 14260
rect 2455 14229 2467 14232
rect 2409 14223 2467 14229
rect 5994 14220 6000 14232
rect 6052 14220 6058 14272
rect 7374 14220 7380 14272
rect 7432 14260 7438 14272
rect 7469 14263 7527 14269
rect 7469 14260 7481 14263
rect 7432 14232 7481 14260
rect 7432 14220 7438 14232
rect 7469 14229 7481 14232
rect 7515 14260 7527 14263
rect 10612 14260 10640 14300
rect 7515 14232 10640 14260
rect 11057 14263 11115 14269
rect 7515 14229 7527 14232
rect 7469 14223 7527 14229
rect 11057 14229 11069 14263
rect 11103 14260 11115 14263
rect 11238 14260 11244 14272
rect 11103 14232 11244 14260
rect 11103 14229 11115 14232
rect 11057 14223 11115 14229
rect 11238 14220 11244 14232
rect 11296 14220 11302 14272
rect 11348 14260 11376 14300
rect 13265 14297 13277 14331
rect 13311 14328 13323 14331
rect 13446 14328 13452 14340
rect 13311 14300 13452 14328
rect 13311 14297 13323 14300
rect 13265 14291 13323 14297
rect 13446 14288 13452 14300
rect 13504 14328 13510 14340
rect 13722 14328 13728 14340
rect 13504 14300 13728 14328
rect 13504 14288 13510 14300
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 17678 14328 17684 14340
rect 17639 14300 17684 14328
rect 17678 14288 17684 14300
rect 17736 14288 17742 14340
rect 13170 14260 13176 14272
rect 11348 14232 13176 14260
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 13354 14220 13360 14272
rect 13412 14260 13418 14272
rect 16114 14260 16120 14272
rect 13412 14232 16120 14260
rect 13412 14220 13418 14232
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 18138 14220 18144 14272
rect 18196 14260 18202 14272
rect 18509 14263 18567 14269
rect 18509 14260 18521 14263
rect 18196 14232 18521 14260
rect 18196 14220 18202 14232
rect 18509 14229 18521 14232
rect 18555 14260 18567 14263
rect 18782 14260 18788 14272
rect 18555 14232 18788 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 19242 14260 19248 14272
rect 19203 14232 19248 14260
rect 19242 14220 19248 14232
rect 19300 14220 19306 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 1765 14059 1823 14065
rect 1765 14025 1777 14059
rect 1811 14056 1823 14059
rect 6086 14056 6092 14068
rect 1811 14028 6092 14056
rect 1811 14025 1823 14028
rect 1765 14019 1823 14025
rect 6086 14016 6092 14028
rect 6144 14016 6150 14068
rect 6546 14016 6552 14068
rect 6604 14056 6610 14068
rect 6604 14028 7788 14056
rect 6604 14016 6610 14028
rect 4709 13991 4767 13997
rect 4709 13957 4721 13991
rect 4755 13988 4767 13991
rect 4890 13988 4896 14000
rect 4755 13960 4896 13988
rect 4755 13957 4767 13960
rect 4709 13951 4767 13957
rect 4890 13948 4896 13960
rect 4948 13948 4954 14000
rect 5074 13948 5080 14000
rect 5132 13988 5138 14000
rect 5534 13988 5540 14000
rect 5132 13960 5540 13988
rect 5132 13948 5138 13960
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 5721 13991 5779 13997
rect 5721 13957 5733 13991
rect 5767 13957 5779 13991
rect 7760 13988 7788 14028
rect 7834 14016 7840 14068
rect 7892 14056 7898 14068
rect 8205 14059 8263 14065
rect 8205 14056 8217 14059
rect 7892 14028 8217 14056
rect 7892 14016 7898 14028
rect 8205 14025 8217 14028
rect 8251 14025 8263 14059
rect 9030 14056 9036 14068
rect 8991 14028 9036 14056
rect 8205 14019 8263 14025
rect 9030 14016 9036 14028
rect 9088 14016 9094 14068
rect 13998 14056 14004 14068
rect 9140 14028 13124 14056
rect 13959 14028 14004 14056
rect 9140 13988 9168 14028
rect 7760 13960 9168 13988
rect 5721 13951 5779 13957
rect 2409 13923 2467 13929
rect 2409 13889 2421 13923
rect 2455 13920 2467 13923
rect 5736 13920 5764 13951
rect 9306 13948 9312 14000
rect 9364 13988 9370 14000
rect 10686 13988 10692 14000
rect 9364 13960 10692 13988
rect 9364 13948 9370 13960
rect 2455 13892 3464 13920
rect 2455 13889 2467 13892
rect 2409 13883 2467 13889
rect 3436 13864 3464 13892
rect 4356 13892 5764 13920
rect 2222 13852 2228 13864
rect 2183 13824 2228 13852
rect 2222 13812 2228 13824
rect 2280 13812 2286 13864
rect 3326 13852 3332 13864
rect 3287 13824 3332 13852
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 3418 13812 3424 13864
rect 3476 13812 3482 13864
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 4356 13852 4384 13892
rect 6178 13880 6184 13932
rect 6236 13920 6242 13932
rect 9508 13929 9536 13960
rect 10686 13948 10692 13960
rect 10744 13948 10750 14000
rect 10781 13991 10839 13997
rect 10781 13957 10793 13991
rect 10827 13988 10839 13991
rect 11698 13988 11704 14000
rect 10827 13960 11704 13988
rect 10827 13957 10839 13960
rect 10781 13951 10839 13957
rect 11698 13948 11704 13960
rect 11756 13948 11762 14000
rect 12158 13948 12164 14000
rect 12216 13988 12222 14000
rect 12437 13991 12495 13997
rect 12437 13988 12449 13991
rect 12216 13960 12449 13988
rect 12216 13948 12222 13960
rect 12437 13957 12449 13960
rect 12483 13957 12495 13991
rect 12437 13951 12495 13957
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6236 13892 6837 13920
rect 6236 13880 6242 13892
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13920 9551 13923
rect 9677 13923 9735 13929
rect 9539 13892 9573 13920
rect 9539 13889 9551 13892
rect 9493 13883 9551 13889
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 11330 13920 11336 13932
rect 9723 13892 11336 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 11330 13880 11336 13892
rect 11388 13880 11394 13932
rect 12710 13920 12716 13932
rect 12544 13892 12716 13920
rect 4120 13824 4384 13852
rect 5537 13855 5595 13861
rect 4120 13812 4126 13824
rect 5537 13821 5549 13855
rect 5583 13852 5595 13855
rect 5902 13852 5908 13864
rect 5583 13824 5908 13852
rect 5583 13821 5595 13824
rect 5537 13815 5595 13821
rect 5902 13812 5908 13824
rect 5960 13812 5966 13864
rect 7092 13855 7150 13861
rect 7092 13821 7104 13855
rect 7138 13852 7150 13855
rect 7374 13852 7380 13864
rect 7138 13824 7380 13852
rect 7138 13821 7150 13824
rect 7092 13815 7150 13821
rect 7374 13812 7380 13824
rect 7432 13812 7438 13864
rect 12544 13852 12572 13892
rect 12710 13880 12716 13892
rect 12768 13880 12774 13932
rect 13096 13929 13124 14028
rect 13998 14016 14004 14028
rect 14056 14016 14062 14068
rect 15562 14056 15568 14068
rect 15523 14028 15568 14056
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 16114 14016 16120 14068
rect 16172 14056 16178 14068
rect 17954 14056 17960 14068
rect 16172 14028 17960 14056
rect 16172 14016 16178 14028
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 13446 13948 13452 14000
rect 13504 13988 13510 14000
rect 18782 13988 18788 14000
rect 13504 13960 18788 13988
rect 13504 13948 13510 13960
rect 18782 13948 18788 13960
rect 18840 13948 18846 14000
rect 13081 13923 13139 13929
rect 13081 13889 13093 13923
rect 13127 13889 13139 13923
rect 13081 13883 13139 13889
rect 13170 13880 13176 13932
rect 13228 13920 13234 13932
rect 14553 13923 14611 13929
rect 14553 13920 14565 13923
rect 13228 13892 14565 13920
rect 13228 13880 13234 13892
rect 14553 13889 14565 13892
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 15562 13880 15568 13932
rect 15620 13920 15626 13932
rect 16022 13920 16028 13932
rect 15620 13892 16028 13920
rect 15620 13880 15626 13892
rect 16022 13880 16028 13892
rect 16080 13880 16086 13932
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 17494 13920 17500 13932
rect 17083 13892 17500 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 12894 13852 12900 13864
rect 7484 13824 12572 13852
rect 12855 13824 12900 13852
rect 2133 13787 2191 13793
rect 2133 13753 2145 13787
rect 2179 13784 2191 13787
rect 2498 13784 2504 13796
rect 2179 13756 2504 13784
rect 2179 13753 2191 13756
rect 2133 13747 2191 13753
rect 2498 13744 2504 13756
rect 2556 13744 2562 13796
rect 2866 13744 2872 13796
rect 2924 13784 2930 13796
rect 3574 13787 3632 13793
rect 3574 13784 3586 13787
rect 2924 13756 3586 13784
rect 2924 13744 2930 13756
rect 3574 13753 3586 13756
rect 3620 13753 3632 13787
rect 3574 13747 3632 13753
rect 5534 13676 5540 13728
rect 5592 13716 5598 13728
rect 7484 13716 7512 13824
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 13814 13812 13820 13864
rect 13872 13852 13878 13864
rect 15749 13855 15807 13861
rect 15749 13852 15761 13855
rect 13872 13824 15761 13852
rect 13872 13812 13878 13824
rect 15749 13821 15761 13824
rect 15795 13821 15807 13855
rect 16850 13852 16856 13864
rect 16811 13824 16856 13852
rect 15749 13815 15807 13821
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 18138 13812 18144 13864
rect 18196 13852 18202 13864
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 18196 13824 18797 13852
rect 18196 13812 18202 13824
rect 18785 13821 18797 13824
rect 18831 13821 18843 13855
rect 18785 13815 18843 13821
rect 19052 13855 19110 13861
rect 19052 13821 19064 13855
rect 19098 13852 19110 13855
rect 20254 13852 20260 13864
rect 19098 13824 20260 13852
rect 19098 13821 19110 13824
rect 19052 13815 19110 13821
rect 8294 13744 8300 13796
rect 8352 13784 8358 13796
rect 9401 13787 9459 13793
rect 9401 13784 9413 13787
rect 8352 13756 9413 13784
rect 8352 13744 8358 13756
rect 9401 13753 9413 13756
rect 9447 13753 9459 13787
rect 9401 13747 9459 13753
rect 10502 13744 10508 13796
rect 10560 13784 10566 13796
rect 11146 13784 11152 13796
rect 10560 13756 11152 13784
rect 10560 13744 10566 13756
rect 11146 13744 11152 13756
rect 11204 13744 11210 13796
rect 11241 13787 11299 13793
rect 11241 13753 11253 13787
rect 11287 13784 11299 13787
rect 11882 13784 11888 13796
rect 11287 13756 11888 13784
rect 11287 13753 11299 13756
rect 11241 13747 11299 13753
rect 11882 13744 11888 13756
rect 11940 13744 11946 13796
rect 12710 13744 12716 13796
rect 12768 13784 12774 13796
rect 14461 13787 14519 13793
rect 14461 13784 14473 13787
rect 12768 13756 14473 13784
rect 12768 13744 12774 13756
rect 14461 13753 14473 13756
rect 14507 13753 14519 13787
rect 18800 13784 18828 13815
rect 20254 13812 20260 13824
rect 20312 13812 20318 13864
rect 19518 13784 19524 13796
rect 18800 13756 19524 13784
rect 14461 13747 14519 13753
rect 19518 13744 19524 13756
rect 19576 13744 19582 13796
rect 5592 13688 7512 13716
rect 5592 13676 5598 13688
rect 8754 13676 8760 13728
rect 8812 13716 8818 13728
rect 9030 13716 9036 13728
rect 8812 13688 9036 13716
rect 8812 13676 8818 13688
rect 9030 13676 9036 13688
rect 9088 13716 9094 13728
rect 9582 13716 9588 13728
rect 9088 13688 9588 13716
rect 9088 13676 9094 13688
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 9858 13676 9864 13728
rect 9916 13716 9922 13728
rect 12805 13719 12863 13725
rect 12805 13716 12817 13719
rect 9916 13688 12817 13716
rect 9916 13676 9922 13688
rect 12805 13685 12817 13688
rect 12851 13685 12863 13719
rect 12805 13679 12863 13685
rect 12986 13676 12992 13728
rect 13044 13716 13050 13728
rect 14369 13719 14427 13725
rect 14369 13716 14381 13719
rect 13044 13688 14381 13716
rect 13044 13676 13050 13688
rect 14369 13685 14381 13688
rect 14415 13685 14427 13719
rect 16390 13716 16396 13728
rect 16351 13688 16396 13716
rect 14369 13679 14427 13685
rect 16390 13676 16396 13688
rect 16448 13676 16454 13728
rect 16758 13716 16764 13728
rect 16719 13688 16764 13716
rect 16758 13676 16764 13688
rect 16816 13676 16822 13728
rect 20162 13716 20168 13728
rect 20123 13688 20168 13716
rect 20162 13676 20168 13688
rect 20220 13676 20226 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 4433 13515 4491 13521
rect 4433 13481 4445 13515
rect 4479 13512 4491 13515
rect 5629 13515 5687 13521
rect 5629 13512 5641 13515
rect 4479 13484 5641 13512
rect 4479 13481 4491 13484
rect 4433 13475 4491 13481
rect 5629 13481 5641 13484
rect 5675 13481 5687 13515
rect 6086 13512 6092 13524
rect 6047 13484 6092 13512
rect 5629 13475 5687 13481
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7469 13515 7527 13521
rect 7469 13512 7481 13515
rect 7156 13484 7481 13512
rect 7156 13472 7162 13484
rect 7469 13481 7481 13484
rect 7515 13481 7527 13515
rect 7469 13475 7527 13481
rect 8021 13515 8079 13521
rect 8021 13481 8033 13515
rect 8067 13512 8079 13515
rect 10137 13515 10195 13521
rect 10137 13512 10149 13515
rect 8067 13484 10149 13512
rect 8067 13481 8079 13484
rect 8021 13475 8079 13481
rect 10137 13481 10149 13484
rect 10183 13481 10195 13515
rect 10137 13475 10195 13481
rect 10686 13472 10692 13524
rect 10744 13472 10750 13524
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 11020 13484 16344 13512
rect 11020 13472 11026 13484
rect 2590 13444 2596 13456
rect 1780 13416 2596 13444
rect 1780 13385 1808 13416
rect 2590 13404 2596 13416
rect 2648 13444 2654 13456
rect 3326 13444 3332 13456
rect 2648 13416 3332 13444
rect 2648 13404 2654 13416
rect 3326 13404 3332 13416
rect 3384 13404 3390 13456
rect 5994 13444 6000 13456
rect 5955 13416 6000 13444
rect 5994 13404 6000 13416
rect 6052 13404 6058 13456
rect 10704 13444 10732 13472
rect 6104 13416 10732 13444
rect 1765 13379 1823 13385
rect 1765 13345 1777 13379
rect 1811 13345 1823 13379
rect 1765 13339 1823 13345
rect 2032 13379 2090 13385
rect 2032 13345 2044 13379
rect 2078 13376 2090 13379
rect 3050 13376 3056 13388
rect 2078 13348 3056 13376
rect 2078 13345 2090 13348
rect 2032 13339 2090 13345
rect 3050 13336 3056 13348
rect 3108 13336 3114 13388
rect 3142 13336 3148 13388
rect 3200 13376 3206 13388
rect 4338 13376 4344 13388
rect 3200 13348 4344 13376
rect 3200 13336 3206 13348
rect 4338 13336 4344 13348
rect 4396 13336 4402 13388
rect 4525 13379 4583 13385
rect 4525 13345 4537 13379
rect 4571 13376 4583 13379
rect 5718 13376 5724 13388
rect 4571 13348 5724 13376
rect 4571 13345 4583 13348
rect 4525 13339 4583 13345
rect 5718 13336 5724 13348
rect 5776 13336 5782 13388
rect 3068 13308 3096 13336
rect 4617 13311 4675 13317
rect 4617 13308 4629 13311
rect 3068 13280 4629 13308
rect 4617 13277 4629 13280
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 5994 13268 6000 13320
rect 6052 13308 6058 13320
rect 6104 13308 6132 13416
rect 11330 13404 11336 13456
rect 11388 13444 11394 13456
rect 11514 13453 11520 13456
rect 11508 13444 11520 13453
rect 11388 13416 11520 13444
rect 11388 13404 11394 13416
rect 11508 13407 11520 13416
rect 11514 13404 11520 13407
rect 11572 13404 11578 13456
rect 13817 13447 13875 13453
rect 13817 13444 13829 13447
rect 11716 13416 13829 13444
rect 7653 13379 7711 13385
rect 7653 13345 7665 13379
rect 7699 13345 7711 13379
rect 7653 13339 7711 13345
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13376 8447 13379
rect 9858 13376 9864 13388
rect 8435 13348 9864 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 6270 13308 6276 13320
rect 6052 13280 6132 13308
rect 6231 13280 6276 13308
rect 6052 13268 6058 13280
rect 6270 13268 6276 13280
rect 6328 13268 6334 13320
rect 7668 13252 7696 13339
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 10045 13379 10103 13385
rect 10045 13345 10057 13379
rect 10091 13376 10103 13379
rect 10686 13376 10692 13388
rect 10091 13348 10692 13376
rect 10091 13345 10103 13348
rect 10045 13339 10103 13345
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 11716 13376 11744 13416
rect 13817 13413 13829 13416
rect 13863 13413 13875 13447
rect 16316 13444 16344 13484
rect 16390 13472 16396 13524
rect 16448 13512 16454 13524
rect 16577 13515 16635 13521
rect 16577 13512 16589 13515
rect 16448 13484 16589 13512
rect 16448 13472 16454 13484
rect 16577 13481 16589 13484
rect 16623 13481 16635 13515
rect 16577 13475 16635 13481
rect 18046 13444 18052 13456
rect 16316 13416 18052 13444
rect 13817 13407 13875 13413
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 10980 13348 11744 13376
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13277 8539 13311
rect 8481 13271 8539 13277
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 8754 13308 8760 13320
rect 8711 13280 8760 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 7650 13200 7656 13252
rect 7708 13200 7714 13252
rect 8496 13240 8524 13271
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 10226 13308 10232 13320
rect 10187 13280 10232 13308
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 9030 13240 9036 13252
rect 8496 13212 9036 13240
rect 9030 13200 9036 13212
rect 9088 13200 9094 13252
rect 9306 13200 9312 13252
rect 9364 13240 9370 13252
rect 10980 13240 11008 13348
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 13538 13376 13544 13388
rect 12676 13348 13544 13376
rect 12676 13336 12682 13348
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 13909 13379 13967 13385
rect 13909 13376 13921 13379
rect 13648 13348 13921 13376
rect 11054 13268 11060 13320
rect 11112 13308 11118 13320
rect 11241 13311 11299 13317
rect 11241 13308 11253 13311
rect 11112 13280 11253 13308
rect 11112 13268 11118 13280
rect 11241 13277 11253 13280
rect 11287 13277 11299 13311
rect 13648 13308 13676 13348
rect 13909 13345 13921 13348
rect 13955 13345 13967 13379
rect 13909 13339 13967 13345
rect 16485 13379 16543 13385
rect 16485 13345 16497 13379
rect 16531 13376 16543 13379
rect 17402 13376 17408 13388
rect 16531 13348 17408 13376
rect 16531 13345 16543 13348
rect 16485 13339 16543 13345
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 17678 13376 17684 13388
rect 17639 13348 17684 13376
rect 17678 13336 17684 13348
rect 17736 13336 17742 13388
rect 17954 13385 17960 13388
rect 17948 13376 17960 13385
rect 17867 13348 17960 13376
rect 17948 13339 17960 13348
rect 18012 13376 18018 13388
rect 18782 13376 18788 13388
rect 18012 13348 18788 13376
rect 17954 13336 17960 13339
rect 18012 13336 18018 13348
rect 18782 13336 18788 13348
rect 18840 13336 18846 13388
rect 13998 13308 14004 13320
rect 11241 13271 11299 13277
rect 12268 13280 13676 13308
rect 13959 13280 14004 13308
rect 9364 13212 11008 13240
rect 9364 13200 9370 13212
rect 2866 13132 2872 13184
rect 2924 13172 2930 13184
rect 3145 13175 3203 13181
rect 3145 13172 3157 13175
rect 2924 13144 3157 13172
rect 2924 13132 2930 13144
rect 3145 13141 3157 13144
rect 3191 13141 3203 13175
rect 4062 13172 4068 13184
rect 4023 13144 4068 13172
rect 3145 13135 3203 13141
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 5810 13132 5816 13184
rect 5868 13172 5874 13184
rect 8294 13172 8300 13184
rect 5868 13144 8300 13172
rect 5868 13132 5874 13144
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 9677 13175 9735 13181
rect 9677 13141 9689 13175
rect 9723 13172 9735 13175
rect 12268 13172 12296 13280
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 16761 13311 16819 13317
rect 16761 13277 16773 13311
rect 16807 13277 16819 13311
rect 16761 13271 16819 13277
rect 9723 13144 12296 13172
rect 9723 13141 9735 13144
rect 9677 13135 9735 13141
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 12621 13175 12679 13181
rect 12621 13172 12633 13175
rect 12492 13144 12633 13172
rect 12492 13132 12498 13144
rect 12621 13141 12633 13144
rect 12667 13172 12679 13175
rect 13170 13172 13176 13184
rect 12667 13144 13176 13172
rect 12667 13141 12679 13144
rect 12621 13135 12679 13141
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 13446 13172 13452 13184
rect 13407 13144 13452 13172
rect 13446 13132 13452 13144
rect 13504 13132 13510 13184
rect 15194 13132 15200 13184
rect 15252 13172 15258 13184
rect 16117 13175 16175 13181
rect 16117 13172 16129 13175
rect 15252 13144 16129 13172
rect 15252 13132 15258 13144
rect 16117 13141 16129 13144
rect 16163 13141 16175 13175
rect 16776 13172 16804 13271
rect 17954 13172 17960 13184
rect 16776 13144 17960 13172
rect 16117 13135 16175 13141
rect 17954 13132 17960 13144
rect 18012 13132 18018 13184
rect 19061 13175 19119 13181
rect 19061 13141 19073 13175
rect 19107 13172 19119 13175
rect 19334 13172 19340 13184
rect 19107 13144 19340 13172
rect 19107 13141 19119 13144
rect 19061 13135 19119 13141
rect 19334 13132 19340 13144
rect 19392 13172 19398 13184
rect 19610 13172 19616 13184
rect 19392 13144 19616 13172
rect 19392 13132 19398 13144
rect 19610 13132 19616 13144
rect 19668 13132 19674 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 5776 12940 6837 12968
rect 5776 12928 5782 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 9861 12971 9919 12977
rect 6825 12931 6883 12937
rect 7300 12940 9444 12968
rect 2590 12792 2596 12844
rect 2648 12832 2654 12844
rect 2869 12835 2927 12841
rect 2869 12832 2881 12835
rect 2648 12804 2881 12832
rect 2648 12792 2654 12804
rect 2869 12801 2881 12804
rect 2915 12801 2927 12835
rect 5629 12835 5687 12841
rect 5629 12832 5641 12835
rect 2869 12795 2927 12801
rect 4264 12804 5641 12832
rect 4264 12776 4292 12804
rect 5629 12801 5641 12804
rect 5675 12832 5687 12835
rect 6270 12832 6276 12844
rect 5675 12804 6276 12832
rect 5675 12801 5687 12804
rect 5629 12795 5687 12801
rect 6270 12792 6276 12804
rect 6328 12792 6334 12844
rect 7300 12841 7328 12940
rect 9416 12900 9444 12940
rect 9861 12937 9873 12971
rect 9907 12968 9919 12971
rect 10226 12968 10232 12980
rect 9907 12940 10232 12968
rect 9907 12937 9919 12940
rect 9861 12931 9919 12937
rect 10226 12928 10232 12940
rect 10284 12928 10290 12980
rect 10686 12968 10692 12980
rect 10647 12940 10692 12968
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 12066 12968 12072 12980
rect 11848 12940 12072 12968
rect 11848 12928 11854 12940
rect 12066 12928 12072 12940
rect 12124 12968 12130 12980
rect 14090 12968 14096 12980
rect 12124 12940 14096 12968
rect 12124 12928 12130 12940
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 17129 12971 17187 12977
rect 17129 12968 17141 12971
rect 17092 12940 17141 12968
rect 17092 12928 17098 12940
rect 17129 12937 17141 12940
rect 17175 12968 17187 12971
rect 17175 12940 18368 12968
rect 17175 12937 17187 12940
rect 17129 12931 17187 12937
rect 18340 12912 18368 12940
rect 18782 12928 18788 12980
rect 18840 12968 18846 12980
rect 20717 12971 20775 12977
rect 20717 12968 20729 12971
rect 18840 12940 20729 12968
rect 18840 12928 18846 12940
rect 20717 12937 20729 12940
rect 20763 12937 20775 12971
rect 20717 12931 20775 12937
rect 10410 12900 10416 12912
rect 9416 12872 10416 12900
rect 10410 12860 10416 12872
rect 10468 12860 10474 12912
rect 11882 12860 11888 12912
rect 11940 12900 11946 12912
rect 14458 12900 14464 12912
rect 11940 12872 14464 12900
rect 11940 12860 11946 12872
rect 14458 12860 14464 12872
rect 14516 12860 14522 12912
rect 18322 12860 18328 12912
rect 18380 12860 18386 12912
rect 19334 12860 19340 12912
rect 19392 12860 19398 12912
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 11238 12832 11244 12844
rect 7377 12795 7435 12801
rect 9876 12804 11244 12832
rect 1581 12767 1639 12773
rect 1581 12733 1593 12767
rect 1627 12764 1639 12767
rect 2406 12764 2412 12776
rect 1627 12736 2412 12764
rect 1627 12733 1639 12736
rect 1581 12727 1639 12733
rect 2406 12724 2412 12736
rect 2464 12724 2470 12776
rect 3136 12767 3194 12773
rect 3136 12733 3148 12767
rect 3182 12764 3194 12767
rect 4246 12764 4252 12776
rect 3182 12736 4252 12764
rect 3182 12733 3194 12736
rect 3136 12727 3194 12733
rect 4246 12724 4252 12736
rect 4304 12724 4310 12776
rect 5074 12764 5080 12776
rect 4724 12736 5080 12764
rect 4724 12708 4752 12736
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 5442 12764 5448 12776
rect 5403 12736 5448 12764
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5534 12724 5540 12776
rect 5592 12764 5598 12776
rect 6288 12764 6316 12792
rect 7392 12764 7420 12795
rect 8754 12773 8760 12776
rect 5592 12736 5637 12764
rect 6288 12736 7420 12764
rect 8481 12767 8539 12773
rect 5592 12724 5598 12736
rect 8481 12733 8493 12767
rect 8527 12733 8539 12767
rect 8748 12764 8760 12773
rect 8667 12736 8760 12764
rect 8481 12727 8539 12733
rect 8748 12727 8760 12736
rect 8812 12764 8818 12776
rect 9876 12764 9904 12804
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 12253 12835 12311 12841
rect 12253 12801 12265 12835
rect 12299 12832 12311 12835
rect 12618 12832 12624 12844
rect 12299 12804 12624 12832
rect 12299 12801 12311 12804
rect 12253 12795 12311 12801
rect 12618 12792 12624 12804
rect 12676 12792 12682 12844
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12768 12804 13001 12832
rect 12768 12792 12774 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 14550 12832 14556 12844
rect 14511 12804 14556 12832
rect 12989 12795 13047 12801
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 15746 12832 15752 12844
rect 15707 12804 15752 12832
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 19352 12832 19380 12860
rect 17972 12804 19380 12832
rect 11054 12764 11060 12776
rect 8812 12736 9904 12764
rect 11015 12736 11060 12764
rect 1854 12696 1860 12708
rect 1815 12668 1860 12696
rect 1854 12656 1860 12668
rect 1912 12656 1918 12708
rect 2516 12668 4375 12696
rect 2516 12640 2544 12668
rect 2498 12588 2504 12640
rect 2556 12588 2562 12640
rect 3050 12588 3056 12640
rect 3108 12628 3114 12640
rect 4249 12631 4307 12637
rect 4249 12628 4261 12631
rect 3108 12600 4261 12628
rect 3108 12588 3114 12600
rect 4249 12597 4261 12600
rect 4295 12597 4307 12631
rect 4347 12628 4375 12668
rect 4706 12656 4712 12708
rect 4764 12656 4770 12708
rect 5092 12696 5120 12724
rect 5092 12668 5948 12696
rect 5077 12631 5135 12637
rect 5077 12628 5089 12631
rect 4347 12600 5089 12628
rect 4249 12591 4307 12597
rect 5077 12597 5089 12600
rect 5123 12597 5135 12631
rect 5920 12628 5948 12668
rect 6730 12656 6736 12708
rect 6788 12696 6794 12708
rect 7193 12699 7251 12705
rect 7193 12696 7205 12699
rect 6788 12668 7205 12696
rect 6788 12656 6794 12668
rect 7193 12665 7205 12668
rect 7239 12665 7251 12699
rect 8496 12696 8524 12727
rect 8754 12724 8760 12727
rect 8812 12724 8818 12736
rect 11054 12724 11060 12736
rect 11112 12724 11118 12776
rect 13446 12764 13452 12776
rect 11164 12736 13452 12764
rect 9674 12696 9680 12708
rect 8496 12668 9680 12696
rect 7193 12659 7251 12665
rect 9674 12656 9680 12668
rect 9732 12656 9738 12708
rect 9766 12656 9772 12708
rect 9824 12696 9830 12708
rect 11164 12696 11192 12736
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 16016 12767 16074 12773
rect 16016 12733 16028 12767
rect 16062 12764 16074 12767
rect 17972 12764 18000 12804
rect 16062 12736 18000 12764
rect 18049 12767 18107 12773
rect 16062 12733 16074 12736
rect 16016 12727 16074 12733
rect 18049 12733 18061 12767
rect 18095 12764 18107 12767
rect 18690 12764 18696 12776
rect 18095 12736 18696 12764
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 18874 12724 18880 12776
rect 18932 12764 18938 12776
rect 19150 12764 19156 12776
rect 18932 12736 19156 12764
rect 18932 12724 18938 12736
rect 19150 12724 19156 12736
rect 19208 12724 19214 12776
rect 19337 12767 19395 12773
rect 19337 12733 19349 12767
rect 19383 12764 19395 12767
rect 19383 12736 19564 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 9824 12668 11192 12696
rect 9824 12656 9830 12668
rect 11422 12656 11428 12708
rect 11480 12696 11486 12708
rect 12897 12699 12955 12705
rect 12897 12696 12909 12699
rect 11480 12668 12909 12696
rect 11480 12656 11486 12668
rect 12897 12665 12909 12668
rect 12943 12665 12955 12699
rect 12897 12659 12955 12665
rect 13262 12656 13268 12708
rect 13320 12696 13326 12708
rect 14461 12699 14519 12705
rect 14461 12696 14473 12699
rect 13320 12668 14473 12696
rect 13320 12656 13326 12668
rect 14461 12665 14473 12668
rect 14507 12665 14519 12699
rect 14461 12659 14519 12665
rect 15286 12656 15292 12708
rect 15344 12696 15350 12708
rect 18230 12696 18236 12708
rect 15344 12668 18236 12696
rect 15344 12656 15350 12668
rect 18230 12656 18236 12668
rect 18288 12656 18294 12708
rect 18325 12699 18383 12705
rect 18325 12665 18337 12699
rect 18371 12696 18383 12699
rect 18598 12696 18604 12708
rect 18371 12668 18604 12696
rect 18371 12665 18383 12668
rect 18325 12659 18383 12665
rect 18598 12656 18604 12668
rect 18656 12656 18662 12708
rect 19536 12640 19564 12736
rect 19604 12699 19662 12705
rect 19604 12665 19616 12699
rect 19650 12696 19662 12699
rect 19978 12696 19984 12708
rect 19650 12668 19984 12696
rect 19650 12665 19662 12668
rect 19604 12659 19662 12665
rect 19978 12656 19984 12668
rect 20036 12656 20042 12708
rect 10502 12628 10508 12640
rect 5920 12600 10508 12628
rect 5077 12591 5135 12597
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 11149 12631 11207 12637
rect 11149 12628 11161 12631
rect 10744 12600 11161 12628
rect 10744 12588 10750 12600
rect 11149 12597 11161 12600
rect 11195 12628 11207 12631
rect 12253 12631 12311 12637
rect 12253 12628 12265 12631
rect 11195 12600 12265 12628
rect 11195 12597 11207 12600
rect 11149 12591 11207 12597
rect 12253 12597 12265 12600
rect 12299 12597 12311 12631
rect 12253 12591 12311 12597
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12802 12628 12808 12640
rect 12492 12600 12537 12628
rect 12763 12600 12808 12628
rect 12492 12588 12498 12600
rect 12802 12588 12808 12600
rect 12860 12588 12866 12640
rect 12986 12588 12992 12640
rect 13044 12628 13050 12640
rect 14001 12631 14059 12637
rect 14001 12628 14013 12631
rect 13044 12600 14013 12628
rect 13044 12588 13050 12600
rect 14001 12597 14013 12600
rect 14047 12597 14059 12631
rect 14001 12591 14059 12597
rect 14090 12588 14096 12640
rect 14148 12628 14154 12640
rect 14369 12631 14427 12637
rect 14369 12628 14381 12631
rect 14148 12600 14381 12628
rect 14148 12588 14154 12600
rect 14369 12597 14381 12600
rect 14415 12597 14427 12631
rect 14369 12591 14427 12597
rect 18506 12588 18512 12640
rect 18564 12628 18570 12640
rect 19518 12628 19524 12640
rect 18564 12600 19524 12628
rect 18564 12588 18570 12600
rect 19518 12588 19524 12600
rect 19576 12588 19582 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 2685 12427 2743 12433
rect 2685 12393 2697 12427
rect 2731 12424 2743 12427
rect 4062 12424 4068 12436
rect 2731 12396 4068 12424
rect 2731 12393 2743 12396
rect 2685 12387 2743 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 6270 12424 6276 12436
rect 6231 12396 6276 12424
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 7190 12384 7196 12436
rect 7248 12424 7254 12436
rect 7466 12424 7472 12436
rect 7248 12396 7472 12424
rect 7248 12384 7254 12396
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 8021 12427 8079 12433
rect 8021 12393 8033 12427
rect 8067 12424 8079 12427
rect 11054 12424 11060 12436
rect 8067 12396 11060 12424
rect 8067 12393 8079 12396
rect 8021 12387 8079 12393
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 11330 12384 11336 12436
rect 11388 12424 11394 12436
rect 12066 12424 12072 12436
rect 11388 12396 12072 12424
rect 11388 12384 11394 12396
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 12253 12427 12311 12433
rect 12253 12393 12265 12427
rect 12299 12424 12311 12427
rect 13998 12424 14004 12436
rect 12299 12396 14004 12424
rect 12299 12393 12311 12396
rect 12253 12387 12311 12393
rect 13998 12384 14004 12396
rect 14056 12384 14062 12436
rect 16132 12396 17612 12424
rect 3418 12316 3424 12368
rect 3476 12356 3482 12368
rect 5160 12359 5218 12365
rect 5160 12356 5172 12359
rect 3476 12328 5172 12356
rect 3476 12316 3482 12328
rect 5160 12325 5172 12328
rect 5206 12356 5218 12359
rect 6546 12356 6552 12368
rect 5206 12328 6552 12356
rect 5206 12325 5218 12328
rect 5160 12319 5218 12325
rect 6546 12316 6552 12328
rect 6604 12316 6610 12368
rect 8386 12356 8392 12368
rect 8299 12328 8392 12356
rect 8386 12316 8392 12328
rect 8444 12356 8450 12368
rect 8662 12356 8668 12368
rect 8444 12328 8668 12356
rect 8444 12316 8450 12328
rect 8662 12316 8668 12328
rect 8720 12316 8726 12368
rect 9490 12316 9496 12368
rect 9548 12356 9554 12368
rect 9944 12359 10002 12365
rect 9548 12328 9812 12356
rect 9548 12316 9554 12328
rect 2222 12248 2228 12300
rect 2280 12288 2286 12300
rect 2593 12291 2651 12297
rect 2593 12288 2605 12291
rect 2280 12260 2605 12288
rect 2280 12248 2286 12260
rect 2593 12257 2605 12260
rect 2639 12257 2651 12291
rect 2593 12251 2651 12257
rect 3326 12248 3332 12300
rect 3384 12288 3390 12300
rect 4893 12291 4951 12297
rect 4893 12288 4905 12291
rect 3384 12260 4905 12288
rect 3384 12248 3390 12260
rect 4893 12257 4905 12260
rect 4939 12257 4951 12291
rect 4893 12251 4951 12257
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 7742 12288 7748 12300
rect 7248 12260 7748 12288
rect 7248 12248 7254 12260
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8202 12288 8208 12300
rect 7975 12260 8208 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 9674 12288 9680 12300
rect 9635 12260 9680 12288
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 9784 12288 9812 12328
rect 9944 12325 9956 12359
rect 9990 12356 10002 12359
rect 10042 12356 10048 12368
rect 9990 12328 10048 12356
rect 9990 12325 10002 12328
rect 9944 12319 10002 12325
rect 10042 12316 10048 12328
rect 10100 12356 10106 12368
rect 10226 12356 10232 12368
rect 10100 12328 10232 12356
rect 10100 12316 10106 12328
rect 10226 12316 10232 12328
rect 10284 12316 10290 12368
rect 10778 12316 10784 12368
rect 10836 12356 10842 12368
rect 11698 12356 11704 12368
rect 10836 12328 11704 12356
rect 10836 12316 10842 12328
rect 11698 12316 11704 12328
rect 11756 12316 11762 12368
rect 15749 12359 15807 12365
rect 15749 12356 15761 12359
rect 12544 12328 15761 12356
rect 12544 12288 12572 12328
rect 15749 12325 15761 12328
rect 15795 12325 15807 12359
rect 15749 12319 15807 12325
rect 9784 12260 12572 12288
rect 12621 12291 12679 12297
rect 12621 12257 12633 12291
rect 12667 12257 12679 12291
rect 12621 12251 12679 12257
rect 13072 12291 13130 12297
rect 13072 12257 13084 12291
rect 13118 12288 13130 12291
rect 13814 12288 13820 12300
rect 13118 12260 13820 12288
rect 13118 12257 13130 12260
rect 13072 12251 13130 12257
rect 2866 12220 2872 12232
rect 2827 12192 2872 12220
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 8478 12220 8484 12232
rect 8439 12192 8484 12220
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12220 8631 12223
rect 9122 12220 9128 12232
rect 8619 12192 9128 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 12250 12180 12256 12232
rect 12308 12220 12314 12232
rect 12636 12220 12664 12251
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 14826 12248 14832 12300
rect 14884 12288 14890 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 14884 12260 15669 12288
rect 14884 12248 14890 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15764 12288 15792 12319
rect 15838 12316 15844 12368
rect 15896 12356 15902 12368
rect 16132 12356 16160 12396
rect 15896 12328 16160 12356
rect 15896 12316 15902 12328
rect 17218 12316 17224 12368
rect 17276 12356 17282 12368
rect 17497 12359 17555 12365
rect 17497 12356 17509 12359
rect 17276 12328 17509 12356
rect 17276 12316 17282 12328
rect 17497 12325 17509 12328
rect 17543 12325 17555 12359
rect 17584 12356 17612 12396
rect 19058 12384 19064 12436
rect 19116 12424 19122 12436
rect 20070 12424 20076 12436
rect 19116 12396 20076 12424
rect 19116 12384 19122 12396
rect 20070 12384 20076 12396
rect 20128 12384 20134 12436
rect 19334 12356 19340 12368
rect 17584 12328 19340 12356
rect 17497 12319 17555 12325
rect 19334 12316 19340 12328
rect 19392 12316 19398 12368
rect 16114 12288 16120 12300
rect 15764 12260 16120 12288
rect 15657 12251 15715 12257
rect 16114 12248 16120 12260
rect 16172 12248 16178 12300
rect 17405 12291 17463 12297
rect 17405 12288 17417 12291
rect 16684 12260 17417 12288
rect 12308 12192 12664 12220
rect 12805 12223 12863 12229
rect 12308 12180 12314 12192
rect 12805 12189 12817 12223
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 2225 12155 2283 12161
rect 2225 12121 2237 12155
rect 2271 12152 2283 12155
rect 3418 12152 3424 12164
rect 2271 12124 3424 12152
rect 2271 12121 2283 12124
rect 2225 12115 2283 12121
rect 3418 12112 3424 12124
rect 3476 12112 3482 12164
rect 3694 12112 3700 12164
rect 3752 12152 3758 12164
rect 4614 12152 4620 12164
rect 3752 12124 4620 12152
rect 3752 12112 3758 12124
rect 4614 12112 4620 12124
rect 4672 12112 4678 12164
rect 7650 12112 7656 12164
rect 7708 12152 7714 12164
rect 7745 12155 7803 12161
rect 7745 12152 7757 12155
rect 7708 12124 7757 12152
rect 7708 12112 7714 12124
rect 7745 12121 7757 12124
rect 7791 12152 7803 12155
rect 8662 12152 8668 12164
rect 7791 12124 8668 12152
rect 7791 12121 7803 12124
rect 7745 12115 7803 12121
rect 8662 12112 8668 12124
rect 8720 12112 8726 12164
rect 11146 12112 11152 12164
rect 11204 12152 11210 12164
rect 11330 12152 11336 12164
rect 11204 12124 11336 12152
rect 11204 12112 11210 12124
rect 11330 12112 11336 12124
rect 11388 12112 11394 12164
rect 12437 12155 12495 12161
rect 12437 12121 12449 12155
rect 12483 12152 12495 12155
rect 12618 12152 12624 12164
rect 12483 12124 12624 12152
rect 12483 12121 12495 12124
rect 12437 12115 12495 12121
rect 12618 12112 12624 12124
rect 12676 12112 12682 12164
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 6914 12084 6920 12096
rect 4120 12056 6920 12084
rect 4120 12044 4126 12056
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 10042 12044 10048 12096
rect 10100 12084 10106 12096
rect 11057 12087 11115 12093
rect 11057 12084 11069 12087
rect 10100 12056 11069 12084
rect 10100 12044 10106 12056
rect 11057 12053 11069 12056
rect 11103 12084 11115 12087
rect 12253 12087 12311 12093
rect 12253 12084 12265 12087
rect 11103 12056 12265 12084
rect 11103 12053 11115 12056
rect 11057 12047 11115 12053
rect 12253 12053 12265 12056
rect 12299 12053 12311 12087
rect 12820 12084 12848 12183
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 15841 12223 15899 12229
rect 15841 12220 15853 12223
rect 15804 12192 15853 12220
rect 15804 12180 15810 12192
rect 15841 12189 15853 12192
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 13078 12084 13084 12096
rect 12820 12056 13084 12084
rect 12253 12047 12311 12053
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 13722 12084 13728 12096
rect 13228 12056 13728 12084
rect 13228 12044 13234 12056
rect 13722 12044 13728 12056
rect 13780 12044 13786 12096
rect 14090 12044 14096 12096
rect 14148 12084 14154 12096
rect 14185 12087 14243 12093
rect 14185 12084 14197 12087
rect 14148 12056 14197 12084
rect 14148 12044 14154 12056
rect 14185 12053 14197 12056
rect 14231 12084 14243 12087
rect 14550 12084 14556 12096
rect 14231 12056 14556 12084
rect 14231 12053 14243 12056
rect 14185 12047 14243 12053
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 14826 12084 14832 12096
rect 14787 12056 14832 12084
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 15289 12087 15347 12093
rect 15289 12053 15301 12087
rect 15335 12084 15347 12087
rect 15838 12084 15844 12096
rect 15335 12056 15844 12084
rect 15335 12053 15347 12056
rect 15289 12047 15347 12053
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 16114 12044 16120 12096
rect 16172 12084 16178 12096
rect 16684 12084 16712 12260
rect 17405 12257 17417 12260
rect 17451 12257 17463 12291
rect 17405 12251 17463 12257
rect 18506 12248 18512 12300
rect 18564 12288 18570 12300
rect 18601 12291 18659 12297
rect 18601 12288 18613 12291
rect 18564 12260 18613 12288
rect 18564 12248 18570 12260
rect 18601 12257 18613 12260
rect 18647 12257 18659 12291
rect 18857 12291 18915 12297
rect 18857 12288 18869 12291
rect 18601 12251 18659 12257
rect 18708 12260 18869 12288
rect 17681 12223 17739 12229
rect 17681 12189 17693 12223
rect 17727 12220 17739 12223
rect 18708 12220 18736 12260
rect 18857 12257 18869 12260
rect 18903 12288 18915 12291
rect 20622 12288 20628 12300
rect 18903 12260 20628 12288
rect 18903 12257 18915 12260
rect 18857 12251 18915 12257
rect 20622 12248 20628 12260
rect 20680 12248 20686 12300
rect 17727 12192 18736 12220
rect 17727 12189 17739 12192
rect 17681 12183 17739 12189
rect 17034 12084 17040 12096
rect 16172 12056 16712 12084
rect 16995 12056 17040 12084
rect 16172 12044 16178 12056
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 19978 12084 19984 12096
rect 19939 12056 19984 12084
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 2222 11880 2228 11892
rect 2183 11852 2228 11880
rect 2222 11840 2228 11852
rect 2280 11840 2286 11892
rect 3789 11883 3847 11889
rect 3789 11849 3801 11883
rect 3835 11849 3847 11883
rect 3789 11843 3847 11849
rect 2498 11704 2504 11756
rect 2556 11744 2562 11756
rect 2685 11747 2743 11753
rect 2685 11744 2697 11747
rect 2556 11716 2697 11744
rect 2556 11704 2562 11716
rect 2685 11713 2697 11716
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 3142 11744 3148 11756
rect 2915 11716 3148 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 3142 11704 3148 11716
rect 3200 11704 3206 11756
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11676 2651 11679
rect 3804 11676 3832 11843
rect 8202 11840 8208 11892
rect 8260 11840 8266 11892
rect 9306 11880 9312 11892
rect 9267 11852 9312 11880
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 11054 11840 11060 11892
rect 11112 11880 11118 11892
rect 13814 11880 13820 11892
rect 11112 11852 13676 11880
rect 13775 11852 13820 11880
rect 11112 11840 11118 11852
rect 8220 11812 8248 11840
rect 11517 11815 11575 11821
rect 8220 11784 9812 11812
rect 9784 11756 9812 11784
rect 11517 11781 11529 11815
rect 11563 11781 11575 11815
rect 13648 11812 13676 11852
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 16393 11883 16451 11889
rect 16393 11849 16405 11883
rect 16439 11880 16451 11883
rect 16758 11880 16764 11892
rect 16439 11852 16764 11880
rect 16439 11849 16451 11852
rect 16393 11843 16451 11849
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 18690 11880 18696 11892
rect 18012 11852 18696 11880
rect 18012 11840 18018 11852
rect 18690 11840 18696 11852
rect 18748 11840 18754 11892
rect 19613 11883 19671 11889
rect 19613 11849 19625 11883
rect 19659 11880 19671 11883
rect 19702 11880 19708 11892
rect 19659 11852 19708 11880
rect 19659 11849 19671 11852
rect 19613 11843 19671 11849
rect 19702 11840 19708 11852
rect 19760 11840 19766 11892
rect 13648 11784 15792 11812
rect 11517 11775 11575 11781
rect 4246 11704 4252 11756
rect 4304 11744 4310 11756
rect 4341 11747 4399 11753
rect 4341 11744 4353 11747
rect 4304 11716 4353 11744
rect 4304 11704 4310 11716
rect 4341 11713 4353 11716
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11744 5779 11747
rect 6638 11744 6644 11756
rect 5767 11716 6644 11744
rect 5767 11713 5779 11716
rect 5721 11707 5779 11713
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 9766 11704 9772 11756
rect 9824 11704 9830 11756
rect 9950 11744 9956 11756
rect 9911 11716 9956 11744
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 10042 11704 10048 11756
rect 10100 11704 10106 11756
rect 11532 11744 11560 11775
rect 15197 11747 15255 11753
rect 15197 11744 15209 11747
rect 11532 11716 12020 11744
rect 2639 11648 3832 11676
rect 5445 11679 5503 11685
rect 2639 11645 2651 11648
rect 2593 11639 2651 11645
rect 5445 11645 5457 11679
rect 5491 11676 5503 11679
rect 6914 11676 6920 11688
rect 5491 11648 6920 11676
rect 5491 11645 5503 11648
rect 5445 11639 5503 11645
rect 6914 11636 6920 11648
rect 6972 11636 6978 11688
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11645 7067 11679
rect 7009 11639 7067 11645
rect 7276 11679 7334 11685
rect 7276 11645 7288 11679
rect 7322 11676 7334 11679
rect 10060 11676 10088 11704
rect 7322 11648 10088 11676
rect 10137 11679 10195 11685
rect 7322 11645 7334 11648
rect 7276 11639 7334 11645
rect 10137 11645 10149 11679
rect 10183 11676 10195 11679
rect 10226 11676 10232 11688
rect 10183 11648 10232 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 2958 11568 2964 11620
rect 3016 11608 3022 11620
rect 3970 11608 3976 11620
rect 3016 11580 3976 11608
rect 3016 11568 3022 11580
rect 3970 11568 3976 11580
rect 4028 11568 4034 11620
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 5258 11608 5264 11620
rect 4203 11580 5264 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 5258 11568 5264 11580
rect 5316 11568 5322 11620
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 6638 11608 6644 11620
rect 5592 11580 6644 11608
rect 5592 11568 5598 11580
rect 6638 11568 6644 11580
rect 6696 11608 6702 11620
rect 7024 11608 7052 11639
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 10410 11685 10416 11688
rect 10404 11676 10416 11685
rect 10371 11648 10416 11676
rect 10404 11639 10416 11648
rect 10410 11636 10416 11639
rect 10468 11636 10474 11688
rect 9677 11611 9735 11617
rect 9677 11608 9689 11611
rect 6696 11580 7052 11608
rect 9416 11580 9689 11608
rect 6696 11568 6702 11580
rect 3694 11500 3700 11552
rect 3752 11540 3758 11552
rect 4249 11543 4307 11549
rect 4249 11540 4261 11543
rect 3752 11512 4261 11540
rect 3752 11500 3758 11512
rect 4249 11509 4261 11512
rect 4295 11509 4307 11543
rect 4249 11503 4307 11509
rect 7742 11500 7748 11552
rect 7800 11540 7806 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 7800 11512 8401 11540
rect 7800 11500 7806 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 8389 11503 8447 11509
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 9416 11540 9444 11580
rect 9677 11577 9689 11580
rect 9723 11577 9735 11611
rect 11992 11608 12020 11716
rect 13832 11716 15209 11744
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11676 12495 11679
rect 13078 11676 13084 11688
rect 12483 11648 13084 11676
rect 12483 11645 12495 11648
rect 12437 11639 12495 11645
rect 13078 11636 13084 11648
rect 13136 11676 13142 11688
rect 13446 11676 13452 11688
rect 13136 11648 13452 11676
rect 13136 11636 13142 11648
rect 13446 11636 13452 11648
rect 13504 11636 13510 11688
rect 12710 11617 12716 11620
rect 12704 11608 12716 11617
rect 11992 11580 12716 11608
rect 9677 11571 9735 11577
rect 12704 11571 12716 11580
rect 12768 11608 12774 11620
rect 13722 11608 13728 11620
rect 12768 11580 13728 11608
rect 12710 11568 12716 11571
rect 12768 11568 12774 11580
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 9272 11512 9444 11540
rect 9769 11543 9827 11549
rect 9272 11500 9278 11512
rect 9769 11509 9781 11543
rect 9815 11540 9827 11543
rect 9858 11540 9864 11552
rect 9815 11512 9864 11540
rect 9815 11509 9827 11512
rect 9769 11503 9827 11509
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 11606 11540 11612 11552
rect 11567 11512 11612 11540
rect 11606 11500 11612 11512
rect 11664 11500 11670 11552
rect 13078 11500 13084 11552
rect 13136 11540 13142 11552
rect 13832 11540 13860 11716
rect 15197 11713 15209 11716
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 15010 11676 15016 11688
rect 14971 11648 15016 11676
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 15764 11676 15792 11784
rect 16500 11784 18644 11812
rect 16500 11676 16528 11784
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 15764 11648 16528 11676
rect 16574 11636 16580 11688
rect 16632 11676 16638 11688
rect 16960 11676 16988 11707
rect 16632 11648 16988 11676
rect 16632 11636 16638 11648
rect 17034 11636 17040 11688
rect 17092 11676 17098 11688
rect 18417 11679 18475 11685
rect 18417 11676 18429 11679
rect 17092 11648 18429 11676
rect 17092 11636 17098 11648
rect 18417 11645 18429 11648
rect 18463 11645 18475 11679
rect 18417 11639 18475 11645
rect 14274 11568 14280 11620
rect 14332 11608 14338 11620
rect 14550 11608 14556 11620
rect 14332 11580 14556 11608
rect 14332 11568 14338 11580
rect 14550 11568 14556 11580
rect 14608 11608 14614 11620
rect 15105 11611 15163 11617
rect 15105 11608 15117 11611
rect 14608 11580 15117 11608
rect 14608 11568 14614 11580
rect 15105 11577 15117 11580
rect 15151 11577 15163 11611
rect 15105 11571 15163 11577
rect 16482 11568 16488 11620
rect 16540 11608 16546 11620
rect 16761 11611 16819 11617
rect 16761 11608 16773 11611
rect 16540 11580 16773 11608
rect 16540 11568 16546 11580
rect 16761 11577 16773 11580
rect 16807 11577 16819 11611
rect 18616 11608 18644 11784
rect 18693 11747 18751 11753
rect 18693 11713 18705 11747
rect 18739 11744 18751 11747
rect 19978 11744 19984 11756
rect 18739 11716 19984 11744
rect 18739 11713 18751 11716
rect 18693 11707 18751 11713
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 20254 11744 20260 11756
rect 20215 11716 20260 11744
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 19981 11611 20039 11617
rect 19981 11608 19993 11611
rect 18616 11580 19993 11608
rect 16761 11571 16819 11577
rect 19981 11577 19993 11580
rect 20027 11608 20039 11611
rect 20346 11608 20352 11620
rect 20027 11580 20352 11608
rect 20027 11577 20039 11580
rect 19981 11571 20039 11577
rect 20346 11568 20352 11580
rect 20404 11568 20410 11620
rect 13136 11512 13860 11540
rect 13136 11500 13142 11512
rect 14458 11500 14464 11552
rect 14516 11540 14522 11552
rect 14645 11543 14703 11549
rect 14645 11540 14657 11543
rect 14516 11512 14657 11540
rect 14516 11500 14522 11512
rect 14645 11509 14657 11512
rect 14691 11509 14703 11543
rect 14645 11503 14703 11509
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 16853 11543 16911 11549
rect 16853 11540 16865 11543
rect 16724 11512 16865 11540
rect 16724 11500 16730 11512
rect 16853 11509 16865 11512
rect 16899 11540 16911 11543
rect 17034 11540 17040 11552
rect 16899 11512 17040 11540
rect 16899 11509 16911 11512
rect 16853 11503 16911 11509
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 18046 11540 18052 11552
rect 18007 11512 18052 11540
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 18509 11543 18567 11549
rect 18509 11509 18521 11543
rect 18555 11540 18567 11543
rect 19150 11540 19156 11552
rect 18555 11512 19156 11540
rect 18555 11509 18567 11512
rect 18509 11503 18567 11509
rect 19150 11500 19156 11512
rect 19208 11500 19214 11552
rect 19521 11543 19579 11549
rect 19521 11509 19533 11543
rect 19567 11540 19579 11543
rect 20070 11540 20076 11552
rect 19567 11512 20076 11540
rect 19567 11509 19579 11512
rect 19521 11503 19579 11509
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 6604 11308 6745 11336
rect 6604 11296 6610 11308
rect 6733 11305 6745 11308
rect 6779 11336 6791 11339
rect 6822 11336 6828 11348
rect 6779 11308 6828 11336
rect 6779 11305 6791 11308
rect 6733 11299 6791 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 7929 11339 7987 11345
rect 7929 11336 7941 11339
rect 7156 11308 7941 11336
rect 7156 11296 7162 11308
rect 7929 11305 7941 11308
rect 7975 11336 7987 11339
rect 8570 11336 8576 11348
rect 7975 11308 8576 11336
rect 7975 11305 7987 11308
rect 7929 11299 7987 11305
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 9766 11296 9772 11348
rect 9824 11336 9830 11348
rect 11793 11339 11851 11345
rect 11793 11336 11805 11339
rect 9824 11308 11805 11336
rect 9824 11296 9830 11308
rect 11793 11305 11805 11308
rect 11839 11336 11851 11339
rect 12250 11336 12256 11348
rect 11839 11308 12256 11336
rect 11839 11305 11851 11308
rect 11793 11299 11851 11305
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 15657 11339 15715 11345
rect 15657 11305 15669 11339
rect 15703 11336 15715 11339
rect 16482 11336 16488 11348
rect 15703 11308 16488 11336
rect 15703 11305 15715 11308
rect 15657 11299 15715 11305
rect 16482 11296 16488 11308
rect 16540 11296 16546 11348
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 19702 11336 19708 11348
rect 19484 11308 19708 11336
rect 19484 11296 19490 11308
rect 19702 11296 19708 11308
rect 19760 11296 19766 11348
rect 4522 11228 4528 11280
rect 4580 11268 4586 11280
rect 10226 11268 10232 11280
rect 4580 11240 10232 11268
rect 4580 11228 4586 11240
rect 10226 11228 10232 11240
rect 10284 11228 10290 11280
rect 12713 11271 12771 11277
rect 12713 11237 12725 11271
rect 12759 11268 12771 11271
rect 13998 11268 14004 11280
rect 12759 11240 14004 11268
rect 12759 11237 12771 11240
rect 12713 11231 12771 11237
rect 13998 11228 14004 11240
rect 14056 11228 14062 11280
rect 14185 11271 14243 11277
rect 14185 11237 14197 11271
rect 14231 11268 14243 11271
rect 15749 11271 15807 11277
rect 14231 11240 15424 11268
rect 14231 11237 14243 11240
rect 14185 11231 14243 11237
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 2777 11203 2835 11209
rect 2777 11200 2789 11203
rect 1443 11172 2789 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 2777 11169 2789 11172
rect 2823 11169 2835 11203
rect 4062 11200 4068 11212
rect 4023 11172 4068 11200
rect 2777 11163 2835 11169
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11200 4399 11203
rect 4706 11200 4712 11212
rect 4387 11172 4712 11200
rect 4387 11169 4399 11172
rect 4341 11163 4399 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5620 11203 5678 11209
rect 5620 11169 5632 11203
rect 5666 11200 5678 11203
rect 6178 11200 6184 11212
rect 5666 11172 6184 11200
rect 5666 11169 5678 11172
rect 5620 11163 5678 11169
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 6972 11172 8616 11200
rect 6972 11160 6978 11172
rect 1854 11092 1860 11144
rect 1912 11132 1918 11144
rect 2406 11132 2412 11144
rect 1912 11104 2412 11132
rect 1912 11092 1918 11104
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3142 11132 3148 11144
rect 3099 11104 3148 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 2884 11064 2912 11095
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11101 5411 11135
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 5353 11095 5411 11101
rect 6371 11104 8033 11132
rect 4706 11064 4712 11076
rect 2884 11036 4712 11064
rect 4706 11024 4712 11036
rect 4764 11024 4770 11076
rect 2406 10996 2412 11008
rect 2367 10968 2412 10996
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 5368 10996 5396 11095
rect 5534 10996 5540 11008
rect 5368 10968 5540 10996
rect 5534 10956 5540 10968
rect 5592 10956 5598 11008
rect 5718 10956 5724 11008
rect 5776 10996 5782 11008
rect 6371 10996 6399 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11101 8171 11135
rect 8588 11132 8616 11172
rect 8662 11160 8668 11212
rect 8720 11200 8726 11212
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 8720 11172 9321 11200
rect 8720 11160 8726 11172
rect 9309 11169 9321 11172
rect 9355 11169 9367 11203
rect 9309 11163 9367 11169
rect 9950 11160 9956 11212
rect 10008 11200 10014 11212
rect 10505 11203 10563 11209
rect 10505 11200 10517 11203
rect 10008 11172 10517 11200
rect 10008 11160 10014 11172
rect 10505 11169 10517 11172
rect 10551 11169 10563 11203
rect 10505 11163 10563 11169
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 12805 11203 12863 11209
rect 12805 11200 12817 11203
rect 12492 11172 12817 11200
rect 12492 11160 12498 11172
rect 12805 11169 12817 11172
rect 12851 11169 12863 11203
rect 12805 11163 12863 11169
rect 13909 11203 13967 11209
rect 13909 11169 13921 11203
rect 13955 11200 13967 11203
rect 15194 11200 15200 11212
rect 13955 11172 15200 11200
rect 13955 11169 13967 11172
rect 13909 11163 13967 11169
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 15396 11200 15424 11240
rect 15749 11237 15761 11271
rect 15795 11268 15807 11271
rect 16666 11268 16672 11280
rect 15795 11240 16672 11268
rect 15795 11237 15807 11240
rect 15749 11231 15807 11237
rect 16666 11228 16672 11240
rect 16724 11228 16730 11280
rect 17494 11228 17500 11280
rect 17552 11277 17558 11280
rect 17552 11271 17616 11277
rect 17552 11237 17570 11271
rect 17604 11237 17616 11271
rect 17552 11231 17616 11237
rect 17552 11228 17558 11231
rect 17862 11228 17868 11280
rect 17920 11268 17926 11280
rect 19978 11268 19984 11280
rect 17920 11240 19984 11268
rect 17920 11228 17926 11240
rect 19978 11228 19984 11240
rect 20036 11228 20042 11280
rect 15396 11172 18368 11200
rect 9490 11132 9496 11144
rect 8588 11104 9496 11132
rect 8113 11095 8171 11101
rect 7742 11024 7748 11076
rect 7800 11064 7806 11076
rect 8128 11064 8156 11095
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 11146 11092 11152 11144
rect 11204 11132 11210 11144
rect 12989 11135 13047 11141
rect 11204 11104 12388 11132
rect 11204 11092 11210 11104
rect 7800 11036 8156 11064
rect 7800 11024 7806 11036
rect 8754 11024 8760 11076
rect 8812 11064 8818 11076
rect 12250 11064 12256 11076
rect 8812 11036 12256 11064
rect 8812 11024 8818 11036
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 12360 11073 12388 11104
rect 12989 11101 13001 11135
rect 13035 11132 13047 11135
rect 13814 11132 13820 11144
rect 13035 11104 13820 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 15838 11132 15844 11144
rect 15799 11104 15844 11132
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 17313 11135 17371 11141
rect 17313 11101 17325 11135
rect 17359 11101 17371 11135
rect 18340 11132 18368 11172
rect 19242 11160 19248 11212
rect 19300 11200 19306 11212
rect 19521 11203 19579 11209
rect 19521 11200 19533 11203
rect 19300 11172 19533 11200
rect 19300 11160 19306 11172
rect 19521 11169 19533 11172
rect 19567 11169 19579 11203
rect 19521 11163 19579 11169
rect 19426 11132 19432 11144
rect 18340 11104 19432 11132
rect 17313 11095 17371 11101
rect 12345 11067 12403 11073
rect 12345 11033 12357 11067
rect 12391 11033 12403 11067
rect 15286 11064 15292 11076
rect 15247 11036 15292 11064
rect 12345 11027 12403 11033
rect 15286 11024 15292 11036
rect 15344 11024 15350 11076
rect 17126 11024 17132 11076
rect 17184 11064 17190 11076
rect 17328 11064 17356 11095
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 19797 11135 19855 11141
rect 19797 11101 19809 11135
rect 19843 11132 19855 11135
rect 20254 11132 20260 11144
rect 19843 11104 20260 11132
rect 19843 11101 19855 11104
rect 19797 11095 19855 11101
rect 20254 11092 20260 11104
rect 20312 11092 20318 11144
rect 17184 11036 17356 11064
rect 17184 11024 17190 11036
rect 7558 10996 7564 11008
rect 5776 10968 6399 10996
rect 7519 10968 7564 10996
rect 5776 10956 5782 10968
rect 7558 10956 7564 10968
rect 7616 10956 7622 11008
rect 8570 10956 8576 11008
rect 8628 10996 8634 11008
rect 9125 10999 9183 11005
rect 9125 10996 9137 10999
rect 8628 10968 9137 10996
rect 8628 10956 8634 10968
rect 9125 10965 9137 10968
rect 9171 10965 9183 10999
rect 9125 10959 9183 10965
rect 9306 10956 9312 11008
rect 9364 10996 9370 11008
rect 15378 10996 15384 11008
rect 9364 10968 15384 10996
rect 9364 10956 9370 10968
rect 15378 10956 15384 10968
rect 15436 10956 15442 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 1118 10752 1124 10804
rect 1176 10792 1182 10804
rect 1486 10792 1492 10804
rect 1176 10764 1492 10792
rect 1176 10752 1182 10764
rect 1486 10752 1492 10764
rect 1544 10752 1550 10804
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 8478 10792 8484 10804
rect 5215 10764 8484 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 9122 10752 9128 10804
rect 9180 10792 9186 10804
rect 9490 10792 9496 10804
rect 9180 10764 9496 10792
rect 9180 10752 9186 10764
rect 9490 10752 9496 10764
rect 9548 10752 9554 10804
rect 10229 10795 10287 10801
rect 10229 10761 10241 10795
rect 10275 10792 10287 10795
rect 10410 10792 10416 10804
rect 10275 10764 10416 10792
rect 10275 10761 10287 10764
rect 10229 10755 10287 10761
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 12437 10795 12495 10801
rect 12437 10761 12449 10795
rect 12483 10792 12495 10795
rect 12802 10792 12808 10804
rect 12483 10764 12808 10792
rect 12483 10761 12495 10764
rect 12437 10755 12495 10761
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 17678 10792 17684 10804
rect 13004 10764 17684 10792
rect 2682 10684 2688 10736
rect 2740 10724 2746 10736
rect 4062 10724 4068 10736
rect 2740 10696 4068 10724
rect 2740 10684 2746 10696
rect 4062 10684 4068 10696
rect 4120 10684 4126 10736
rect 8570 10724 8576 10736
rect 5092 10696 8576 10724
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2498 10656 2504 10668
rect 2363 10628 2504 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 3881 10659 3939 10665
rect 3881 10656 3893 10659
rect 3200 10628 3893 10656
rect 3200 10616 3206 10628
rect 3881 10625 3893 10628
rect 3927 10656 3939 10659
rect 3970 10656 3976 10668
rect 3927 10628 3976 10656
rect 3927 10625 3939 10628
rect 3881 10619 3939 10625
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10588 2099 10591
rect 2406 10588 2412 10600
rect 2087 10560 2412 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 3326 10588 3332 10600
rect 2700 10560 3332 10588
rect 2133 10523 2191 10529
rect 2133 10489 2145 10523
rect 2179 10520 2191 10523
rect 2700 10520 2728 10560
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 3605 10591 3663 10597
rect 3605 10557 3617 10591
rect 3651 10588 3663 10591
rect 3694 10588 3700 10600
rect 3651 10560 3700 10588
rect 3651 10557 3663 10560
rect 3605 10551 3663 10557
rect 3694 10548 3700 10560
rect 3752 10548 3758 10600
rect 5092 10597 5120 10696
rect 8570 10684 8576 10696
rect 8628 10684 8634 10736
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 5718 10656 5724 10668
rect 5675 10628 5724 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 5077 10591 5135 10597
rect 5077 10557 5089 10591
rect 5123 10557 5135 10591
rect 5077 10551 5135 10557
rect 5534 10548 5540 10600
rect 5592 10548 5598 10600
rect 5552 10520 5580 10548
rect 2179 10492 2728 10520
rect 4908 10492 5580 10520
rect 5828 10520 5856 10619
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7616 10628 7757 10656
rect 7616 10616 7622 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10656 7987 10659
rect 8478 10656 8484 10668
rect 7975 10628 8484 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 10428 10656 10456 10752
rect 12710 10684 12716 10736
rect 12768 10724 12774 10736
rect 13004 10724 13032 10764
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 20070 10752 20076 10804
rect 20128 10792 20134 10804
rect 20622 10792 20628 10804
rect 20128 10764 20628 10792
rect 20128 10752 20134 10764
rect 20622 10752 20628 10764
rect 20680 10792 20686 10804
rect 20809 10795 20867 10801
rect 20809 10792 20821 10795
rect 20680 10764 20821 10792
rect 20680 10752 20686 10764
rect 20809 10761 20821 10764
rect 20855 10761 20867 10795
rect 20809 10755 20867 10761
rect 15565 10727 15623 10733
rect 12768 10696 13032 10724
rect 13096 10696 14964 10724
rect 12768 10684 12774 10696
rect 13096 10668 13124 10696
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 10428 10628 13001 10656
rect 12989 10625 13001 10628
rect 13035 10656 13047 10659
rect 13078 10656 13084 10668
rect 13035 10628 13084 10656
rect 13035 10625 13047 10628
rect 12989 10619 13047 10625
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 14274 10656 14280 10668
rect 14200 10628 14280 10656
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10588 7711 10591
rect 8386 10588 8392 10600
rect 7699 10560 8392 10588
rect 7699 10557 7711 10560
rect 7653 10551 7711 10557
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 8849 10591 8907 10597
rect 8849 10588 8861 10591
rect 8812 10560 8861 10588
rect 8812 10548 8818 10560
rect 8849 10557 8861 10560
rect 8895 10588 8907 10591
rect 10134 10588 10140 10600
rect 8895 10560 10140 10588
rect 8895 10557 8907 10560
rect 8849 10551 8907 10557
rect 10134 10548 10140 10560
rect 10192 10548 10198 10600
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10588 11115 10591
rect 14200 10588 14228 10628
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 14458 10656 14464 10668
rect 14419 10628 14464 10656
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 14645 10659 14703 10665
rect 14645 10625 14657 10659
rect 14691 10656 14703 10659
rect 14826 10656 14832 10668
rect 14691 10628 14832 10656
rect 14691 10625 14703 10628
rect 14645 10619 14703 10625
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 14936 10656 14964 10696
rect 15565 10693 15577 10727
rect 15611 10724 15623 10727
rect 15746 10724 15752 10736
rect 15611 10696 15752 10724
rect 15611 10693 15623 10696
rect 15565 10687 15623 10693
rect 15746 10684 15752 10696
rect 15804 10684 15810 10736
rect 17696 10724 17724 10752
rect 18230 10724 18236 10736
rect 17696 10696 18236 10724
rect 18230 10684 18236 10696
rect 18288 10684 18294 10736
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 14936 10628 16129 10656
rect 16117 10625 16129 10628
rect 16163 10625 16175 10659
rect 16117 10619 16175 10625
rect 17313 10591 17371 10597
rect 17313 10588 17325 10591
rect 11103 10560 14228 10588
rect 14261 10560 17325 10588
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 9122 10529 9128 10532
rect 9094 10523 9128 10529
rect 9094 10520 9106 10523
rect 5828 10492 9106 10520
rect 2179 10489 2191 10492
rect 2133 10483 2191 10489
rect 1670 10452 1676 10464
rect 1631 10424 1676 10452
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 3234 10452 3240 10464
rect 3195 10424 3240 10452
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 3694 10412 3700 10464
rect 3752 10452 3758 10464
rect 4908 10461 4936 10492
rect 9094 10489 9106 10492
rect 9180 10520 9186 10532
rect 9180 10492 9242 10520
rect 9094 10483 9128 10489
rect 9122 10480 9128 10483
rect 9180 10480 9186 10492
rect 9674 10480 9680 10532
rect 9732 10520 9738 10532
rect 11333 10523 11391 10529
rect 11333 10520 11345 10523
rect 9732 10492 11345 10520
rect 9732 10480 9738 10492
rect 11333 10489 11345 10492
rect 11379 10489 11391 10523
rect 11333 10483 11391 10489
rect 12342 10480 12348 10532
rect 12400 10520 12406 10532
rect 14261 10520 14289 10560
rect 17313 10557 17325 10560
rect 17359 10557 17371 10591
rect 18046 10588 18052 10600
rect 18007 10560 18052 10588
rect 17313 10551 17371 10557
rect 18046 10548 18052 10560
rect 18104 10548 18110 10600
rect 19242 10548 19248 10600
rect 19300 10588 19306 10600
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 19300 10560 19441 10588
rect 19300 10548 19306 10560
rect 19429 10557 19441 10560
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 12400 10492 14289 10520
rect 14369 10523 14427 10529
rect 12400 10480 12406 10492
rect 14369 10489 14381 10523
rect 14415 10520 14427 10523
rect 14458 10520 14464 10532
rect 14415 10492 14464 10520
rect 14415 10489 14427 10492
rect 14369 10483 14427 10489
rect 14458 10480 14464 10492
rect 14516 10480 14522 10532
rect 15562 10480 15568 10532
rect 15620 10520 15626 10532
rect 16025 10523 16083 10529
rect 16025 10520 16037 10523
rect 15620 10492 16037 10520
rect 15620 10480 15626 10492
rect 16025 10489 16037 10492
rect 16071 10489 16083 10523
rect 16025 10483 16083 10489
rect 16482 10480 16488 10532
rect 16540 10520 16546 10532
rect 18325 10523 18383 10529
rect 18325 10520 18337 10523
rect 16540 10492 18337 10520
rect 16540 10480 16546 10492
rect 18325 10489 18337 10492
rect 18371 10489 18383 10523
rect 18325 10483 18383 10489
rect 19696 10523 19754 10529
rect 19696 10489 19708 10523
rect 19742 10520 19754 10523
rect 19886 10520 19892 10532
rect 19742 10492 19892 10520
rect 19742 10489 19754 10492
rect 19696 10483 19754 10489
rect 19886 10480 19892 10492
rect 19944 10480 19950 10532
rect 21082 10480 21088 10532
rect 21140 10520 21146 10532
rect 22738 10520 22744 10532
rect 21140 10492 22744 10520
rect 21140 10480 21146 10492
rect 22738 10480 22744 10492
rect 22796 10480 22802 10532
rect 4893 10455 4951 10461
rect 3752 10424 3797 10452
rect 3752 10412 3758 10424
rect 4893 10421 4905 10455
rect 4939 10421 4951 10455
rect 4893 10415 4951 10421
rect 5537 10455 5595 10461
rect 5537 10421 5549 10455
rect 5583 10452 5595 10455
rect 7098 10452 7104 10464
rect 5583 10424 7104 10452
rect 5583 10421 5595 10424
rect 5537 10415 5595 10421
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 7282 10452 7288 10464
rect 7243 10424 7288 10452
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 9306 10452 9312 10464
rect 7524 10424 9312 10452
rect 7524 10412 7530 10424
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12805 10455 12863 10461
rect 12805 10452 12817 10455
rect 12492 10424 12817 10452
rect 12492 10412 12498 10424
rect 12805 10421 12817 10424
rect 12851 10421 12863 10455
rect 12805 10415 12863 10421
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13078 10452 13084 10464
rect 12943 10424 13084 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13078 10412 13084 10424
rect 13136 10452 13142 10464
rect 13262 10452 13268 10464
rect 13136 10424 13268 10452
rect 13136 10412 13142 10424
rect 13262 10412 13268 10424
rect 13320 10412 13326 10464
rect 13998 10452 14004 10464
rect 13959 10424 14004 10452
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 15746 10412 15752 10464
rect 15804 10452 15810 10464
rect 15933 10455 15991 10461
rect 15933 10452 15945 10455
rect 15804 10424 15945 10452
rect 15804 10412 15810 10424
rect 15933 10421 15945 10424
rect 15979 10421 15991 10455
rect 17126 10452 17132 10464
rect 17087 10424 17132 10452
rect 15933 10415 15991 10421
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 1670 10208 1676 10260
rect 1728 10248 1734 10260
rect 2593 10251 2651 10257
rect 2593 10248 2605 10251
rect 1728 10220 2605 10248
rect 1728 10208 1734 10220
rect 2593 10217 2605 10220
rect 2639 10217 2651 10251
rect 2593 10211 2651 10217
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 8478 10248 8484 10260
rect 4028 10220 8484 10248
rect 4028 10208 4034 10220
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 8662 10208 8668 10260
rect 8720 10248 8726 10260
rect 12342 10248 12348 10260
rect 8720 10220 11008 10248
rect 12303 10220 12348 10248
rect 8720 10208 8726 10220
rect 2774 10140 2780 10192
rect 2832 10180 2838 10192
rect 3418 10180 3424 10192
rect 2832 10152 3424 10180
rect 2832 10140 2838 10152
rect 3418 10140 3424 10152
rect 3476 10140 3482 10192
rect 5534 10180 5540 10192
rect 4816 10152 5540 10180
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 3694 10112 3700 10124
rect 2731 10084 3700 10112
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 3694 10072 3700 10084
rect 3752 10072 3758 10124
rect 4816 10121 4844 10152
rect 5534 10140 5540 10152
rect 5592 10180 5598 10192
rect 5718 10180 5724 10192
rect 5592 10152 5724 10180
rect 5592 10140 5598 10152
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 7368 10183 7426 10189
rect 7368 10149 7380 10183
rect 7414 10180 7426 10183
rect 7742 10180 7748 10192
rect 7414 10152 7748 10180
rect 7414 10149 7426 10152
rect 7368 10143 7426 10149
rect 7742 10140 7748 10152
rect 7800 10140 7806 10192
rect 10870 10140 10876 10192
rect 10928 10140 10934 10192
rect 10980 10180 11008 10220
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 13814 10248 13820 10260
rect 12492 10220 13820 10248
rect 12492 10208 12498 10220
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 14185 10251 14243 10257
rect 14185 10217 14197 10251
rect 14231 10248 14243 10251
rect 16114 10248 16120 10260
rect 14231 10220 16120 10248
rect 14231 10217 14243 10220
rect 14185 10211 14243 10217
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 17494 10248 17500 10260
rect 17455 10220 17500 10248
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 12894 10180 12900 10192
rect 10980 10152 12900 10180
rect 12894 10140 12900 10152
rect 12952 10140 12958 10192
rect 12989 10183 13047 10189
rect 12989 10149 13001 10183
rect 13035 10180 13047 10183
rect 13262 10180 13268 10192
rect 13035 10152 13268 10180
rect 13035 10149 13047 10152
rect 12989 10143 13047 10149
rect 13262 10140 13268 10152
rect 13320 10140 13326 10192
rect 15562 10140 15568 10192
rect 15620 10180 15626 10192
rect 15746 10180 15752 10192
rect 15620 10152 15752 10180
rect 15620 10140 15626 10152
rect 15746 10140 15752 10152
rect 15804 10140 15810 10192
rect 16384 10183 16442 10189
rect 16384 10149 16396 10183
rect 16430 10180 16442 10183
rect 16574 10180 16580 10192
rect 16430 10152 16580 10180
rect 16430 10149 16442 10152
rect 16384 10143 16442 10149
rect 16574 10140 16580 10152
rect 16632 10140 16638 10192
rect 18690 10140 18696 10192
rect 18748 10180 18754 10192
rect 18846 10183 18904 10189
rect 18846 10180 18858 10183
rect 18748 10152 18858 10180
rect 18748 10140 18754 10152
rect 18846 10149 18858 10152
rect 18892 10149 18904 10183
rect 18846 10143 18904 10149
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 5068 10115 5126 10121
rect 5068 10081 5080 10115
rect 5114 10112 5126 10115
rect 6546 10112 6552 10124
rect 5114 10084 6552 10112
rect 5114 10081 5126 10084
rect 5068 10075 5126 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 6638 10072 6644 10124
rect 6696 10112 6702 10124
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 6696 10084 7113 10112
rect 6696 10072 6702 10084
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 10778 10112 10784 10124
rect 10739 10084 10784 10112
rect 7101 10075 7159 10081
rect 10778 10072 10784 10084
rect 10836 10072 10842 10124
rect 10888 10112 10916 10140
rect 12529 10115 12587 10121
rect 10888 10084 11008 10112
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 10980 10053 11008 10084
rect 12529 10081 12541 10115
rect 12575 10112 12587 10115
rect 12618 10112 12624 10124
rect 12575 10084 12624 10112
rect 12575 10081 12587 10084
rect 12529 10075 12587 10081
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10112 13139 10115
rect 13998 10112 14004 10124
rect 13127 10084 14004 10112
rect 13127 10081 13139 10084
rect 13081 10075 13139 10081
rect 13998 10072 14004 10084
rect 14056 10072 14062 10124
rect 17126 10112 17132 10124
rect 16132 10084 17132 10112
rect 10873 10047 10931 10053
rect 10873 10044 10885 10047
rect 8352 10016 10885 10044
rect 8352 10004 8358 10016
rect 10873 10013 10885 10016
rect 10919 10013 10931 10047
rect 10873 10007 10931 10013
rect 10965 10047 11023 10053
rect 10965 10013 10977 10047
rect 11011 10013 11023 10047
rect 10965 10007 11023 10013
rect 12342 10004 12348 10056
rect 12400 10044 12406 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12400 10016 13185 10044
rect 12400 10004 12406 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 15746 10004 15752 10056
rect 15804 10044 15810 10056
rect 16132 10053 16160 10084
rect 17126 10072 17132 10084
rect 17184 10112 17190 10124
rect 18046 10112 18052 10124
rect 17184 10084 18052 10112
rect 17184 10072 17190 10084
rect 18046 10072 18052 10084
rect 18104 10112 18110 10124
rect 18601 10115 18659 10121
rect 18601 10112 18613 10115
rect 18104 10084 18613 10112
rect 18104 10072 18110 10084
rect 18601 10081 18613 10084
rect 18647 10112 18659 10115
rect 19242 10112 19248 10124
rect 18647 10084 19248 10112
rect 18647 10081 18659 10084
rect 18601 10075 18659 10081
rect 19242 10072 19248 10084
rect 19300 10072 19306 10124
rect 16117 10047 16175 10053
rect 16117 10044 16129 10047
rect 15804 10016 16129 10044
rect 15804 10004 15810 10016
rect 16117 10013 16129 10016
rect 16163 10013 16175 10047
rect 16117 10007 16175 10013
rect 566 9936 572 9988
rect 624 9976 630 9988
rect 4522 9976 4528 9988
rect 624 9948 4528 9976
rect 624 9936 630 9948
rect 4522 9936 4528 9948
rect 4580 9936 4586 9988
rect 12710 9976 12716 9988
rect 5736 9948 6316 9976
rect 1762 9868 1768 9920
rect 1820 9908 1826 9920
rect 2225 9911 2283 9917
rect 2225 9908 2237 9911
rect 1820 9880 2237 9908
rect 1820 9868 1826 9880
rect 2225 9877 2237 9880
rect 2271 9877 2283 9911
rect 2225 9871 2283 9877
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 5736 9908 5764 9948
rect 6178 9908 6184 9920
rect 2832 9880 5764 9908
rect 6139 9880 6184 9908
rect 2832 9868 2838 9880
rect 6178 9868 6184 9880
rect 6236 9868 6242 9920
rect 6288 9908 6316 9948
rect 8036 9948 12716 9976
rect 8036 9908 8064 9948
rect 12710 9936 12716 9948
rect 12768 9936 12774 9988
rect 17862 9976 17868 9988
rect 17052 9948 17868 9976
rect 10410 9908 10416 9920
rect 6288 9880 8064 9908
rect 10371 9880 10416 9908
rect 10410 9868 10416 9880
rect 10468 9868 10474 9920
rect 10502 9868 10508 9920
rect 10560 9908 10566 9920
rect 11054 9908 11060 9920
rect 10560 9880 11060 9908
rect 10560 9868 10566 9880
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 12618 9908 12624 9920
rect 12579 9880 12624 9908
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 17052 9908 17080 9948
rect 17862 9936 17868 9948
rect 17920 9936 17926 9988
rect 12860 9880 17080 9908
rect 12860 9868 12866 9880
rect 19886 9868 19892 9920
rect 19944 9908 19950 9920
rect 19981 9911 20039 9917
rect 19981 9908 19993 9911
rect 19944 9880 19993 9908
rect 19944 9868 19950 9880
rect 19981 9877 19993 9880
rect 20027 9877 20039 9911
rect 19981 9871 20039 9877
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 2682 9664 2688 9716
rect 2740 9704 2746 9716
rect 3694 9704 3700 9716
rect 2740 9676 3556 9704
rect 3655 9676 3700 9704
rect 2740 9664 2746 9676
rect 1210 9596 1216 9648
rect 1268 9636 1274 9648
rect 1486 9636 1492 9648
rect 1268 9608 1492 9636
rect 1268 9596 1274 9608
rect 1486 9596 1492 9608
rect 1544 9596 1550 9648
rect 2498 9596 2504 9648
rect 2556 9636 2562 9648
rect 2869 9639 2927 9645
rect 2869 9636 2881 9639
rect 2556 9608 2881 9636
rect 2556 9596 2562 9608
rect 2869 9605 2881 9608
rect 2915 9605 2927 9639
rect 3528 9636 3556 9676
rect 3694 9664 3700 9676
rect 3752 9664 3758 9716
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 9122 9704 9128 9716
rect 4120 9676 8984 9704
rect 9083 9676 9128 9704
rect 4120 9664 4126 9676
rect 3970 9636 3976 9648
rect 3528 9608 3976 9636
rect 2869 9599 2927 9605
rect 2884 9568 2912 9599
rect 3970 9596 3976 9608
rect 4028 9596 4034 9648
rect 8956 9636 8984 9676
rect 9122 9664 9128 9676
rect 9180 9664 9186 9716
rect 12802 9704 12808 9716
rect 9232 9676 12808 9704
rect 9232 9636 9260 9676
rect 12802 9664 12808 9676
rect 12860 9664 12866 9716
rect 12894 9664 12900 9716
rect 12952 9704 12958 9716
rect 16482 9704 16488 9716
rect 12952 9676 16488 9704
rect 12952 9664 12958 9676
rect 16482 9664 16488 9676
rect 16540 9664 16546 9716
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 16632 9676 19012 9704
rect 16632 9664 16638 9676
rect 8956 9608 9260 9636
rect 10597 9639 10655 9645
rect 10597 9605 10609 9639
rect 10643 9636 10655 9639
rect 11514 9636 11520 9648
rect 10643 9608 11520 9636
rect 10643 9605 10655 9608
rect 10597 9599 10655 9605
rect 11514 9596 11520 9608
rect 11572 9596 11578 9648
rect 15289 9639 15347 9645
rect 15289 9636 15301 9639
rect 14936 9608 15301 9636
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 2884 9540 4261 9568
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 4249 9531 4307 9537
rect 6638 9528 6644 9580
rect 6696 9568 6702 9580
rect 7558 9568 7564 9580
rect 6696 9540 7564 9568
rect 6696 9528 6702 9540
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 10410 9528 10416 9580
rect 10468 9568 10474 9580
rect 11057 9571 11115 9577
rect 11057 9568 11069 9571
rect 10468 9540 11069 9568
rect 10468 9528 10474 9540
rect 11057 9537 11069 9540
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9537 11207 9571
rect 11149 9531 11207 9537
rect 1486 9500 1492 9512
rect 1447 9472 1492 9500
rect 1486 9460 1492 9472
rect 1544 9460 1550 9512
rect 3234 9460 3240 9512
rect 3292 9500 3298 9512
rect 4065 9503 4123 9509
rect 4065 9500 4077 9503
rect 3292 9472 4077 9500
rect 3292 9460 3298 9472
rect 4065 9469 4077 9472
rect 4111 9469 4123 9503
rect 4065 9463 4123 9469
rect 5166 9460 5172 9512
rect 5224 9500 5230 9512
rect 5261 9503 5319 9509
rect 5261 9500 5273 9503
rect 5224 9472 5273 9500
rect 5224 9460 5230 9472
rect 5261 9469 5273 9472
rect 5307 9469 5319 9503
rect 7742 9500 7748 9512
rect 7703 9472 7748 9500
rect 5261 9463 5319 9469
rect 7742 9460 7748 9472
rect 7800 9460 7806 9512
rect 8012 9503 8070 9509
rect 8012 9469 8024 9503
rect 8058 9500 8070 9503
rect 11164 9500 11192 9531
rect 8058 9472 11192 9500
rect 12621 9503 12679 9509
rect 8058 9469 8070 9472
rect 8012 9463 8070 9469
rect 11072 9444 11100 9472
rect 12621 9469 12633 9503
rect 12667 9500 12679 9503
rect 12802 9500 12808 9512
rect 12667 9472 12808 9500
rect 12667 9469 12679 9472
rect 12621 9463 12679 9469
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 13446 9460 13452 9512
rect 13504 9500 13510 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13504 9472 13921 9500
rect 13504 9460 13510 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 14458 9460 14464 9512
rect 14516 9500 14522 9512
rect 14936 9500 14964 9608
rect 15289 9605 15301 9608
rect 15335 9636 15347 9639
rect 18984 9636 19012 9676
rect 19978 9664 19984 9716
rect 20036 9704 20042 9716
rect 20438 9704 20444 9716
rect 20036 9676 20444 9704
rect 20036 9664 20042 9676
rect 20438 9664 20444 9676
rect 20496 9664 20502 9716
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 21082 9704 21088 9716
rect 20772 9676 21088 9704
rect 20772 9664 20778 9676
rect 21082 9664 21088 9676
rect 21140 9664 21146 9716
rect 21174 9664 21180 9716
rect 21232 9704 21238 9716
rect 21358 9704 21364 9716
rect 21232 9676 21364 9704
rect 21232 9664 21238 9676
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 19429 9639 19487 9645
rect 19429 9636 19441 9639
rect 15335 9608 16712 9636
rect 18984 9608 19441 9636
rect 15335 9605 15347 9608
rect 15289 9599 15347 9605
rect 15930 9528 15936 9580
rect 15988 9568 15994 9580
rect 16684 9577 16712 9608
rect 19429 9605 19441 9608
rect 19475 9605 19487 9639
rect 19429 9599 19487 9605
rect 16577 9571 16635 9577
rect 16577 9568 16589 9571
rect 15988 9540 16589 9568
rect 15988 9528 15994 9540
rect 16577 9537 16589 9540
rect 16623 9537 16635 9571
rect 16577 9531 16635 9537
rect 16669 9571 16727 9577
rect 16669 9537 16681 9571
rect 16715 9537 16727 9571
rect 18046 9568 18052 9580
rect 18007 9540 18052 9568
rect 16669 9531 16727 9537
rect 18046 9528 18052 9540
rect 18104 9528 18110 9580
rect 14516 9472 14964 9500
rect 14516 9460 14522 9472
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 16485 9503 16543 9509
rect 16485 9500 16497 9503
rect 15344 9472 16497 9500
rect 15344 9460 15350 9472
rect 16485 9469 16497 9472
rect 16531 9469 16543 9503
rect 20254 9500 20260 9512
rect 20215 9472 20260 9500
rect 16485 9463 16543 9469
rect 20254 9460 20260 9472
rect 20312 9460 20318 9512
rect 1756 9435 1814 9441
rect 1756 9401 1768 9435
rect 1802 9432 1814 9435
rect 2682 9432 2688 9444
rect 1802 9404 2688 9432
rect 1802 9401 1814 9404
rect 1756 9395 1814 9401
rect 2682 9392 2688 9404
rect 2740 9392 2746 9444
rect 5537 9435 5595 9441
rect 5537 9432 5549 9435
rect 3252 9404 5549 9432
rect 3252 9376 3280 9404
rect 5537 9401 5549 9404
rect 5583 9401 5595 9435
rect 5537 9395 5595 9401
rect 5902 9392 5908 9444
rect 5960 9432 5966 9444
rect 5960 9404 7420 9432
rect 5960 9392 5966 9404
rect 3234 9324 3240 9376
rect 3292 9324 3298 9376
rect 4157 9367 4215 9373
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 7282 9364 7288 9376
rect 4203 9336 7288 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 7392 9364 7420 9404
rect 7558 9392 7564 9444
rect 7616 9432 7622 9444
rect 10686 9432 10692 9444
rect 7616 9404 10692 9432
rect 7616 9392 7622 9404
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 11054 9392 11060 9444
rect 11112 9392 11118 9444
rect 12897 9435 12955 9441
rect 12897 9401 12909 9435
rect 12943 9401 12955 9435
rect 12897 9395 12955 9401
rect 14176 9435 14234 9441
rect 14176 9401 14188 9435
rect 14222 9432 14234 9435
rect 15194 9432 15200 9444
rect 14222 9404 15200 9432
rect 14222 9401 14234 9404
rect 14176 9395 14234 9401
rect 10410 9364 10416 9376
rect 7392 9336 10416 9364
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 10965 9367 11023 9373
rect 10965 9333 10977 9367
rect 11011 9364 11023 9367
rect 11882 9364 11888 9376
rect 11011 9336 11888 9364
rect 11011 9333 11023 9336
rect 10965 9327 11023 9333
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 12912 9364 12940 9395
rect 15194 9392 15200 9404
rect 15252 9432 15258 9444
rect 15838 9432 15844 9444
rect 15252 9404 15844 9432
rect 15252 9392 15258 9404
rect 15838 9392 15844 9404
rect 15896 9392 15902 9444
rect 17678 9392 17684 9444
rect 17736 9432 17742 9444
rect 18294 9435 18352 9441
rect 18294 9432 18306 9435
rect 17736 9404 18306 9432
rect 17736 9392 17742 9404
rect 18294 9401 18306 9404
rect 18340 9401 18352 9435
rect 18294 9395 18352 9401
rect 19978 9392 19984 9444
rect 20036 9432 20042 9444
rect 20533 9435 20591 9441
rect 20533 9432 20545 9435
rect 20036 9404 20545 9432
rect 20036 9392 20042 9404
rect 20533 9401 20545 9404
rect 20579 9401 20591 9435
rect 20533 9395 20591 9401
rect 15378 9364 15384 9376
rect 12912 9336 15384 9364
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 16114 9364 16120 9376
rect 16075 9336 16120 9364
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 17310 9364 17316 9376
rect 16816 9336 17316 9364
rect 16816 9324 16822 9336
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 1486 9160 1492 9172
rect 1412 9132 1492 9160
rect 1412 9024 1440 9132
rect 1486 9120 1492 9132
rect 1544 9120 1550 9172
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 3145 9163 3203 9169
rect 3145 9160 3157 9163
rect 2924 9132 3157 9160
rect 2924 9120 2930 9132
rect 3145 9129 3157 9132
rect 3191 9129 3203 9163
rect 4246 9160 4252 9172
rect 4207 9132 4252 9160
rect 3145 9123 3203 9129
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 5902 9160 5908 9172
rect 4908 9132 5908 9160
rect 2032 9027 2090 9033
rect 1412 8996 1808 9024
rect 1780 8965 1808 8996
rect 2032 8993 2044 9027
rect 2078 9024 2090 9027
rect 2498 9024 2504 9036
rect 2078 8996 2504 9024
rect 2078 8993 2090 8996
rect 2032 8987 2090 8993
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 4028 8996 4077 9024
rect 4028 8984 4034 8996
rect 4065 8993 4077 8996
rect 4111 9024 4123 9027
rect 4908 9024 4936 9132
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 6546 9160 6552 9172
rect 6507 9132 6552 9160
rect 6546 9120 6552 9132
rect 6604 9120 6610 9172
rect 8021 9163 8079 9169
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 8294 9160 8300 9172
rect 8067 9132 8300 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 9030 9160 9036 9172
rect 8444 9132 9036 9160
rect 8444 9120 8450 9132
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 9122 9120 9128 9172
rect 9180 9160 9186 9172
rect 9490 9160 9496 9172
rect 9180 9132 9496 9160
rect 9180 9120 9186 9132
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 10042 9120 10048 9172
rect 10100 9160 10106 9172
rect 10686 9160 10692 9172
rect 10100 9132 10692 9160
rect 10100 9120 10106 9132
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 11054 9160 11060 9172
rect 11015 9132 11060 9160
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11882 9160 11888 9172
rect 11843 9132 11888 9160
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 12253 9163 12311 9169
rect 12253 9129 12265 9163
rect 12299 9160 12311 9163
rect 13449 9163 13507 9169
rect 13449 9160 13461 9163
rect 12299 9132 13461 9160
rect 12299 9129 12311 9132
rect 12253 9123 12311 9129
rect 13449 9129 13461 9132
rect 13495 9129 13507 9163
rect 13449 9123 13507 9129
rect 15473 9163 15531 9169
rect 15473 9129 15485 9163
rect 15519 9160 15531 9163
rect 15654 9160 15660 9172
rect 15519 9132 15660 9160
rect 15519 9129 15531 9132
rect 15473 9123 15531 9129
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 17310 9120 17316 9172
rect 17368 9160 17374 9172
rect 17586 9160 17592 9172
rect 17368 9132 17592 9160
rect 17368 9120 17374 9132
rect 17586 9120 17592 9132
rect 17644 9120 17650 9172
rect 19150 9120 19156 9172
rect 19208 9160 19214 9172
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 19208 9132 19257 9160
rect 19208 9120 19214 9132
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 19610 9160 19616 9172
rect 19571 9132 19616 9160
rect 19245 9123 19303 9129
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 5166 9092 5172 9104
rect 5040 9064 5172 9092
rect 5040 9052 5046 9064
rect 5166 9052 5172 9064
rect 5224 9052 5230 9104
rect 5436 9095 5494 9101
rect 5436 9061 5448 9095
rect 5482 9092 5494 9095
rect 5534 9092 5540 9104
rect 5482 9064 5540 9092
rect 5482 9061 5494 9064
rect 5436 9055 5494 9061
rect 5534 9052 5540 9064
rect 5592 9052 5598 9104
rect 8570 9092 8576 9104
rect 7944 9064 8576 9092
rect 5718 9024 5724 9036
rect 4111 8996 4936 9024
rect 5184 8996 5724 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8925 1823 8959
rect 1765 8919 1823 8925
rect 1780 8820 1808 8919
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 2958 8956 2964 8968
rect 2832 8928 2964 8956
rect 2832 8916 2838 8928
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 4246 8916 4252 8968
rect 4304 8956 4310 8968
rect 4798 8956 4804 8968
rect 4304 8928 4804 8956
rect 4304 8916 4310 8928
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 5184 8965 5212 8996
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 7944 9033 7972 9064
rect 8570 9052 8576 9064
rect 8628 9052 8634 9104
rect 12066 9092 12072 9104
rect 8680 9064 12072 9092
rect 7929 9027 7987 9033
rect 7929 8993 7941 9027
rect 7975 8993 7987 9027
rect 8386 9024 8392 9036
rect 8347 8996 8392 9024
rect 7929 8987 7987 8993
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 8680 9024 8708 9064
rect 12066 9052 12072 9064
rect 12124 9052 12130 9104
rect 12345 9095 12403 9101
rect 12345 9061 12357 9095
rect 12391 9092 12403 9095
rect 12618 9092 12624 9104
rect 12391 9064 12624 9092
rect 12391 9061 12403 9064
rect 12345 9055 12403 9061
rect 12618 9052 12624 9064
rect 12676 9052 12682 9104
rect 12710 9052 12716 9104
rect 12768 9092 12774 9104
rect 13817 9095 13875 9101
rect 13817 9092 13829 9095
rect 12768 9064 13829 9092
rect 12768 9052 12774 9064
rect 13817 9061 13829 9064
rect 13863 9061 13875 9095
rect 15930 9092 15936 9104
rect 13817 9055 13875 9061
rect 13924 9064 15936 9092
rect 8588 8996 8708 9024
rect 8588 8968 8616 8996
rect 9306 8984 9312 9036
rect 9364 9024 9370 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 9364 8996 9689 9024
rect 9364 8984 9370 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 9944 9027 10002 9033
rect 9944 8993 9956 9027
rect 9990 9024 10002 9027
rect 9990 8996 10916 9024
rect 9990 8993 10002 8996
rect 9944 8987 10002 8993
rect 10888 8968 10916 8996
rect 11606 8984 11612 9036
rect 11664 9024 11670 9036
rect 13924 9033 13952 9064
rect 15930 9052 15936 9064
rect 15988 9052 15994 9104
rect 16482 9052 16488 9104
rect 16540 9092 16546 9104
rect 18230 9092 18236 9104
rect 16540 9064 18236 9092
rect 16540 9052 16546 9064
rect 18230 9052 18236 9064
rect 18288 9052 18294 9104
rect 19702 9052 19708 9104
rect 19760 9052 19766 9104
rect 13909 9027 13967 9033
rect 13909 9024 13921 9027
rect 11664 8996 13921 9024
rect 11664 8984 11670 8996
rect 13909 8993 13921 8996
rect 13955 8993 13967 9027
rect 15286 9024 15292 9036
rect 15247 8996 15292 9024
rect 13909 8987 13967 8993
rect 15286 8984 15292 8996
rect 15344 8984 15350 9036
rect 16752 9027 16810 9033
rect 16752 8993 16764 9027
rect 16798 9024 16810 9027
rect 17586 9024 17592 9036
rect 16798 8996 17592 9024
rect 16798 8993 16810 8996
rect 16752 8987 16810 8993
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 19720 9024 19748 9052
rect 19720 8996 19840 9024
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8925 5227 8959
rect 5169 8919 5227 8925
rect 2958 8820 2964 8832
rect 1780 8792 2964 8820
rect 2958 8780 2964 8792
rect 3016 8820 3022 8832
rect 5184 8820 5212 8919
rect 7374 8916 7380 8968
rect 7432 8956 7438 8968
rect 8481 8959 8539 8965
rect 8481 8956 8493 8959
rect 7432 8928 8493 8956
rect 7432 8916 7438 8928
rect 8481 8925 8493 8928
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 8570 8916 8576 8968
rect 8628 8916 8634 8968
rect 8665 8959 8723 8965
rect 8665 8925 8677 8959
rect 8711 8956 8723 8959
rect 9582 8956 9588 8968
rect 8711 8928 9588 8956
rect 8711 8925 8723 8928
rect 8665 8919 8723 8925
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 10870 8916 10876 8968
rect 10928 8956 10934 8968
rect 12437 8959 12495 8965
rect 12437 8956 12449 8959
rect 10928 8928 12449 8956
rect 10928 8916 10934 8928
rect 12437 8925 12449 8928
rect 12483 8925 12495 8959
rect 14001 8959 14059 8965
rect 14001 8956 14013 8959
rect 12437 8919 12495 8925
rect 13740 8928 14013 8956
rect 9030 8848 9036 8900
rect 9088 8888 9094 8900
rect 9088 8860 9260 8888
rect 9088 8848 9094 8860
rect 7742 8820 7748 8832
rect 3016 8792 5212 8820
rect 7655 8792 7748 8820
rect 3016 8780 3022 8792
rect 7742 8780 7748 8792
rect 7800 8820 7806 8832
rect 8754 8820 8760 8832
rect 7800 8792 8760 8820
rect 7800 8780 7806 8792
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9232 8820 9260 8860
rect 13740 8832 13768 8928
rect 14001 8925 14013 8928
rect 14047 8925 14059 8959
rect 14001 8919 14059 8925
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 16485 8959 16543 8965
rect 16485 8956 16497 8959
rect 15896 8928 16497 8956
rect 15896 8916 15902 8928
rect 16485 8925 16497 8928
rect 16531 8925 16543 8959
rect 19702 8956 19708 8968
rect 19663 8928 19708 8956
rect 16485 8919 16543 8925
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 18230 8848 18236 8900
rect 18288 8888 18294 8900
rect 19610 8888 19616 8900
rect 18288 8860 19616 8888
rect 18288 8848 18294 8860
rect 19610 8848 19616 8860
rect 19668 8848 19674 8900
rect 12710 8820 12716 8832
rect 9232 8792 12716 8820
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 13722 8780 13728 8832
rect 13780 8780 13786 8832
rect 14274 8780 14280 8832
rect 14332 8820 14338 8832
rect 15654 8820 15660 8832
rect 14332 8792 15660 8820
rect 14332 8780 14338 8792
rect 15654 8780 15660 8792
rect 15712 8780 15718 8832
rect 17678 8780 17684 8832
rect 17736 8820 17742 8832
rect 17865 8823 17923 8829
rect 17865 8820 17877 8823
rect 17736 8792 17877 8820
rect 17736 8780 17742 8792
rect 17865 8789 17877 8792
rect 17911 8789 17923 8823
rect 19812 8820 19840 8996
rect 19889 8959 19947 8965
rect 19889 8925 19901 8959
rect 19935 8956 19947 8959
rect 20070 8956 20076 8968
rect 19935 8928 20076 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 20070 8916 20076 8928
rect 20128 8916 20134 8968
rect 20070 8820 20076 8832
rect 19812 8792 20076 8820
rect 17865 8783 17923 8789
rect 20070 8780 20076 8792
rect 20128 8780 20134 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 2958 8576 2964 8628
rect 3016 8576 3022 8628
rect 3510 8576 3516 8628
rect 3568 8616 3574 8628
rect 4525 8619 4583 8625
rect 3568 8588 4200 8616
rect 3568 8576 3574 8588
rect 2976 8548 3004 8576
rect 2976 8520 3188 8548
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 2958 8480 2964 8492
rect 2087 8452 2964 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 3160 8489 3188 8520
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 1762 8412 1768 8424
rect 1723 8384 1768 8412
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 4172 8412 4200 8588
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 5534 8616 5540 8628
rect 4571 8588 5540 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 6788 8588 6837 8616
rect 6788 8576 6794 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 10318 8616 10324 8628
rect 6825 8579 6883 8585
rect 8404 8588 10324 8616
rect 7558 8508 7564 8560
rect 7616 8508 7622 8560
rect 5626 8480 5632 8492
rect 5587 8452 5632 8480
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 6880 8452 7389 8480
rect 6880 8440 6886 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 5353 8415 5411 8421
rect 5353 8412 5365 8415
rect 4172 8384 5365 8412
rect 5353 8381 5365 8384
rect 5399 8381 5411 8415
rect 5353 8375 5411 8381
rect 7098 8372 7104 8424
rect 7156 8412 7162 8424
rect 7193 8415 7251 8421
rect 7193 8412 7205 8415
rect 7156 8384 7205 8412
rect 7156 8372 7162 8384
rect 7193 8381 7205 8384
rect 7239 8381 7251 8415
rect 7193 8375 7251 8381
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 7576 8412 7604 8508
rect 8404 8489 8432 8588
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 10870 8616 10876 8628
rect 10827 8588 10876 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 15286 8616 15292 8628
rect 13832 8588 15292 8616
rect 12250 8508 12256 8560
rect 12308 8508 12314 8560
rect 12618 8508 12624 8560
rect 12676 8548 12682 8560
rect 12894 8548 12900 8560
rect 12676 8520 12900 8548
rect 12676 8508 12682 8520
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 8812 8452 9352 8480
rect 8812 8440 8818 8452
rect 9324 8424 9352 8452
rect 7331 8384 7604 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 9030 8412 9036 8424
rect 8628 8384 9036 8412
rect 8628 8372 8634 8384
rect 9030 8372 9036 8384
rect 9088 8372 9094 8424
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 12268 8421 12296 8508
rect 12713 8483 12771 8489
rect 12713 8449 12725 8483
rect 12759 8480 12771 8483
rect 13832 8480 13860 8588
rect 15286 8576 15292 8588
rect 15344 8576 15350 8628
rect 15654 8576 15660 8628
rect 15712 8616 15718 8628
rect 16025 8619 16083 8625
rect 16025 8616 16037 8619
rect 15712 8588 16037 8616
rect 15712 8576 15718 8588
rect 16025 8585 16037 8588
rect 16071 8585 16083 8619
rect 16025 8579 16083 8585
rect 18233 8619 18291 8625
rect 18233 8585 18245 8619
rect 18279 8616 18291 8619
rect 18874 8616 18880 8628
rect 18279 8588 18880 8616
rect 18279 8585 18291 8588
rect 18233 8579 18291 8585
rect 18874 8576 18880 8588
rect 18932 8576 18938 8628
rect 15197 8551 15255 8557
rect 15197 8517 15209 8551
rect 15243 8548 15255 8551
rect 15562 8548 15568 8560
rect 15243 8520 15568 8548
rect 15243 8517 15255 8520
rect 15197 8511 15255 8517
rect 15562 8508 15568 8520
rect 15620 8548 15626 8560
rect 15620 8520 16620 8548
rect 15620 8508 15626 8520
rect 12759 8452 13860 8480
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 16114 8440 16120 8492
rect 16172 8480 16178 8492
rect 16592 8489 16620 8520
rect 18046 8508 18052 8560
rect 18104 8548 18110 8560
rect 18104 8520 19196 8548
rect 18104 8508 18110 8520
rect 19168 8492 19196 8520
rect 16485 8483 16543 8489
rect 16485 8480 16497 8483
rect 16172 8452 16497 8480
rect 16172 8440 16178 8452
rect 16485 8449 16497 8452
rect 16531 8449 16543 8483
rect 16485 8443 16543 8449
rect 16577 8483 16635 8489
rect 16577 8449 16589 8483
rect 16623 8449 16635 8483
rect 19150 8480 19156 8492
rect 19063 8452 19156 8480
rect 16577 8443 16635 8449
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 9364 8384 9413 8412
rect 9364 8372 9370 8384
rect 9401 8381 9413 8384
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8381 12311 8415
rect 12253 8375 12311 8381
rect 12434 8372 12440 8424
rect 12492 8412 12498 8424
rect 13446 8412 13452 8424
rect 12492 8384 12537 8412
rect 12820 8384 13452 8412
rect 12492 8372 12498 8384
rect 2866 8304 2872 8356
rect 2924 8344 2930 8356
rect 3390 8347 3448 8353
rect 3390 8344 3402 8347
rect 2924 8316 3402 8344
rect 2924 8304 2930 8316
rect 3390 8313 3402 8316
rect 3436 8313 3448 8347
rect 3390 8307 3448 8313
rect 4062 8304 4068 8356
rect 4120 8344 4126 8356
rect 8754 8344 8760 8356
rect 4120 8316 8760 8344
rect 4120 8304 4126 8316
rect 8754 8304 8760 8316
rect 8812 8304 8818 8356
rect 9582 8304 9588 8356
rect 9640 8353 9646 8356
rect 9640 8347 9704 8353
rect 9640 8313 9658 8347
rect 9692 8344 9704 8347
rect 11330 8344 11336 8356
rect 9692 8316 11336 8344
rect 9692 8313 9704 8316
rect 9640 8307 9704 8313
rect 9640 8304 9646 8307
rect 11330 8304 11336 8316
rect 11388 8304 11394 8356
rect 12820 8344 12848 8384
rect 13446 8372 13452 8384
rect 13504 8412 13510 8424
rect 13817 8415 13875 8421
rect 13817 8412 13829 8415
rect 13504 8384 13829 8412
rect 13504 8372 13510 8384
rect 13817 8381 13829 8384
rect 13863 8381 13875 8415
rect 13817 8375 13875 8381
rect 14084 8415 14142 8421
rect 14084 8381 14096 8415
rect 14130 8412 14142 8415
rect 14458 8412 14464 8424
rect 14130 8384 14464 8412
rect 14130 8381 14142 8384
rect 14084 8375 14142 8381
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 17218 8412 17224 8424
rect 16776 8384 17224 8412
rect 12360 8316 12848 8344
rect 12360 8288 12388 8316
rect 12894 8304 12900 8356
rect 12952 8344 12958 8356
rect 13170 8344 13176 8356
rect 12952 8316 13176 8344
rect 12952 8304 12958 8316
rect 13170 8304 13176 8316
rect 13228 8304 13234 8356
rect 15286 8304 15292 8356
rect 15344 8344 15350 8356
rect 16393 8347 16451 8353
rect 16393 8344 16405 8347
rect 15344 8316 16405 8344
rect 15344 8304 15350 8316
rect 16393 8313 16405 8316
rect 16439 8313 16451 8347
rect 16393 8307 16451 8313
rect 8478 8236 8484 8288
rect 8536 8276 8542 8288
rect 9030 8276 9036 8288
rect 8536 8248 9036 8276
rect 8536 8236 8542 8248
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 12069 8279 12127 8285
rect 12069 8245 12081 8279
rect 12115 8276 12127 8279
rect 12342 8276 12348 8288
rect 12115 8248 12348 8276
rect 12115 8245 12127 8248
rect 12069 8239 12127 8245
rect 12342 8236 12348 8248
rect 12400 8236 12406 8288
rect 13262 8236 13268 8288
rect 13320 8276 13326 8288
rect 13446 8276 13452 8288
rect 13320 8248 13452 8276
rect 13320 8236 13326 8248
rect 13446 8236 13452 8248
rect 13504 8236 13510 8288
rect 14274 8236 14280 8288
rect 14332 8276 14338 8288
rect 16776 8276 16804 8384
rect 17218 8372 17224 8384
rect 17276 8412 17282 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17276 8384 18061 8412
rect 17276 8372 17282 8384
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 19420 8415 19478 8421
rect 19420 8381 19432 8415
rect 19466 8412 19478 8415
rect 20162 8412 20168 8424
rect 19466 8384 20168 8412
rect 19466 8381 19478 8384
rect 19420 8375 19478 8381
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 20530 8372 20536 8424
rect 20588 8412 20594 8424
rect 20898 8412 20904 8424
rect 20588 8384 20904 8412
rect 20588 8372 20594 8384
rect 20898 8372 20904 8384
rect 20956 8372 20962 8424
rect 14332 8248 16804 8276
rect 14332 8236 14338 8248
rect 17126 8236 17132 8288
rect 17184 8276 17190 8288
rect 17770 8276 17776 8288
rect 17184 8248 17776 8276
rect 17184 8236 17190 8248
rect 17770 8236 17776 8248
rect 17828 8236 17834 8288
rect 20162 8236 20168 8288
rect 20220 8276 20226 8288
rect 20346 8276 20352 8288
rect 20220 8248 20352 8276
rect 20220 8236 20226 8248
rect 20346 8236 20352 8248
rect 20404 8236 20410 8288
rect 20530 8276 20536 8288
rect 20491 8248 20536 8276
rect 20530 8236 20536 8248
rect 20588 8236 20594 8288
rect 20622 8236 20628 8288
rect 20680 8276 20686 8288
rect 21450 8276 21456 8288
rect 20680 8248 21456 8276
rect 20680 8236 20686 8248
rect 21450 8236 21456 8248
rect 21508 8236 21514 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 5445 8075 5503 8081
rect 5445 8041 5457 8075
rect 5491 8072 5503 8075
rect 6549 8075 6607 8081
rect 6549 8072 6561 8075
rect 5491 8044 6561 8072
rect 5491 8041 5503 8044
rect 5445 8035 5503 8041
rect 6549 8041 6561 8044
rect 6595 8041 6607 8075
rect 6549 8035 6607 8041
rect 9861 8075 9919 8081
rect 9861 8041 9873 8075
rect 9907 8072 9919 8075
rect 10502 8072 10508 8084
rect 9907 8044 10508 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 10778 8072 10784 8084
rect 10739 8044 10784 8072
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 10870 8032 10876 8084
rect 10928 8072 10934 8084
rect 14274 8072 14280 8084
rect 10928 8044 14280 8072
rect 10928 8032 10934 8044
rect 14274 8032 14280 8044
rect 14332 8032 14338 8084
rect 15396 8044 15976 8072
rect 1854 7964 1860 8016
rect 1912 8004 1918 8016
rect 2498 8004 2504 8016
rect 1912 7976 2504 8004
rect 1912 7964 1918 7976
rect 2498 7964 2504 7976
rect 2556 7964 2562 8016
rect 2682 7964 2688 8016
rect 2740 8004 2746 8016
rect 3602 8004 3608 8016
rect 2740 7976 3608 8004
rect 2740 7964 2746 7976
rect 3602 7964 3608 7976
rect 3660 7964 3666 8016
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 11054 8004 11060 8016
rect 4120 7976 8248 8004
rect 4120 7964 4126 7976
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2590 7936 2596 7948
rect 2179 7908 2596 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 2590 7896 2596 7908
rect 2648 7896 2654 7948
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 5353 7939 5411 7945
rect 5353 7936 5365 7939
rect 4948 7908 5365 7936
rect 4948 7896 4954 7908
rect 5353 7905 5365 7908
rect 5399 7905 5411 7939
rect 5353 7899 5411 7905
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 6880 7908 6929 7936
rect 6880 7896 6886 7908
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 1854 7828 1860 7880
rect 1912 7868 1918 7880
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 1912 7840 2329 7868
rect 1912 7828 1918 7840
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7868 5687 7871
rect 6178 7868 6184 7880
rect 5675 7840 6184 7868
rect 5675 7837 5687 7840
rect 5629 7831 5687 7837
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 7006 7868 7012 7880
rect 6967 7840 7012 7868
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 2130 7760 2136 7812
rect 2188 7800 2194 7812
rect 2406 7800 2412 7812
rect 2188 7772 2412 7800
rect 2188 7760 2194 7772
rect 2406 7760 2412 7772
rect 2464 7760 2470 7812
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 4120 7772 5120 7800
rect 4120 7760 4126 7772
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 4985 7735 5043 7741
rect 4985 7732 4997 7735
rect 1820 7704 4997 7732
rect 1820 7692 1826 7704
rect 4985 7701 4997 7704
rect 5031 7701 5043 7735
rect 5092 7732 5120 7772
rect 6546 7760 6552 7812
rect 6604 7800 6610 7812
rect 7116 7800 7144 7831
rect 6604 7772 7144 7800
rect 8220 7800 8248 7976
rect 8312 7976 11060 8004
rect 8312 7945 8340 7976
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 11149 8007 11207 8013
rect 11149 7973 11161 8007
rect 11195 8004 11207 8007
rect 11698 8004 11704 8016
rect 11195 7976 11704 8004
rect 11195 7973 11207 7976
rect 11149 7967 11207 7973
rect 11698 7964 11704 7976
rect 11756 8004 11762 8016
rect 12066 8004 12072 8016
rect 11756 7976 12072 8004
rect 11756 7964 11762 7976
rect 12066 7964 12072 7976
rect 12124 7964 12130 8016
rect 12250 8004 12256 8016
rect 12167 7976 12256 8004
rect 8297 7939 8355 7945
rect 8297 7905 8309 7939
rect 8343 7905 8355 7939
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 8297 7899 8355 7905
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10502 7936 10508 7948
rect 10008 7908 10508 7936
rect 10008 7896 10014 7908
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 11238 7936 11244 7948
rect 11151 7908 11244 7936
rect 11238 7896 11244 7908
rect 11296 7936 11302 7948
rect 11882 7936 11888 7948
rect 11296 7908 11888 7936
rect 11296 7896 11302 7908
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 12167 7936 12195 7976
rect 12250 7964 12256 7976
rect 12308 8004 12314 8016
rect 12612 8007 12670 8013
rect 12308 7976 12401 8004
rect 12308 7964 12314 7976
rect 11992 7908 12195 7936
rect 12367 7936 12395 7976
rect 12612 7973 12624 8007
rect 12658 8004 12670 8007
rect 15396 8004 15424 8044
rect 15562 8013 15568 8016
rect 15556 8004 15568 8013
rect 12658 7976 15424 8004
rect 15523 7976 15568 8004
rect 12658 7973 12670 7976
rect 12612 7967 12670 7973
rect 15556 7967 15568 7976
rect 15562 7964 15568 7967
rect 15620 7964 15626 8016
rect 15948 8004 15976 8044
rect 17402 8032 17408 8084
rect 17460 8072 17466 8084
rect 17497 8075 17555 8081
rect 17497 8072 17509 8075
rect 17460 8044 17509 8072
rect 17460 8032 17466 8044
rect 17497 8041 17509 8044
rect 17543 8041 17555 8075
rect 17497 8035 17555 8041
rect 17862 8032 17868 8084
rect 17920 8072 17926 8084
rect 18046 8072 18052 8084
rect 17920 8044 18052 8072
rect 17920 8032 17926 8044
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 19245 8075 19303 8081
rect 19245 8041 19257 8075
rect 19291 8072 19303 8075
rect 19702 8072 19708 8084
rect 19291 8044 19708 8072
rect 19291 8041 19303 8044
rect 19245 8035 19303 8041
rect 19702 8032 19708 8044
rect 19760 8032 19766 8084
rect 20346 8004 20352 8016
rect 15948 7976 20352 8004
rect 20346 7964 20352 7976
rect 20404 7964 20410 8016
rect 13722 7936 13728 7948
rect 12367 7908 13728 7936
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7868 8631 7871
rect 10134 7868 10140 7880
rect 8619 7840 10140 7868
rect 8619 7837 8631 7840
rect 8573 7831 8631 7837
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 11330 7868 11336 7880
rect 11291 7840 11336 7868
rect 11330 7828 11336 7840
rect 11388 7868 11394 7880
rect 11992 7868 12020 7908
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 15289 7939 15347 7945
rect 15289 7905 15301 7939
rect 15335 7936 15347 7939
rect 15838 7936 15844 7948
rect 15335 7908 15844 7936
rect 15335 7905 15347 7908
rect 15289 7899 15347 7905
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 16666 7896 16672 7948
rect 16724 7936 16730 7948
rect 17402 7936 17408 7948
rect 16724 7908 17408 7936
rect 16724 7896 16730 7908
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 17862 7936 17868 7948
rect 17823 7908 17868 7936
rect 17862 7896 17868 7908
rect 17920 7896 17926 7948
rect 18874 7896 18880 7948
rect 18932 7936 18938 7948
rect 19153 7939 19211 7945
rect 19153 7936 19165 7939
rect 18932 7908 19165 7936
rect 18932 7896 18938 7908
rect 19153 7905 19165 7908
rect 19199 7936 19211 7939
rect 19613 7939 19671 7945
rect 19613 7936 19625 7939
rect 19199 7908 19625 7936
rect 19199 7905 19211 7908
rect 19153 7899 19211 7905
rect 19613 7905 19625 7908
rect 19659 7936 19671 7939
rect 20622 7936 20628 7948
rect 19659 7908 20628 7936
rect 19659 7905 19671 7908
rect 19613 7899 19671 7905
rect 20622 7896 20628 7908
rect 20680 7896 20686 7948
rect 12342 7868 12348 7880
rect 11388 7840 12020 7868
rect 12303 7840 12348 7868
rect 11388 7828 11394 7840
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 9858 7800 9864 7812
rect 8220 7772 9864 7800
rect 6604 7760 6610 7772
rect 9858 7760 9864 7772
rect 9916 7800 9922 7812
rect 11698 7800 11704 7812
rect 9916 7772 11704 7800
rect 9916 7760 9922 7772
rect 11698 7760 11704 7772
rect 11756 7760 11762 7812
rect 13740 7809 13768 7896
rect 17770 7828 17776 7880
rect 17828 7868 17834 7880
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 17828 7840 17969 7868
rect 17828 7828 17834 7840
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7837 19763 7871
rect 19886 7868 19892 7880
rect 19847 7840 19892 7868
rect 19705 7831 19763 7837
rect 13725 7803 13783 7809
rect 13725 7769 13737 7803
rect 13771 7769 13783 7803
rect 13725 7763 13783 7769
rect 17494 7760 17500 7812
rect 17552 7800 17558 7812
rect 18064 7800 18092 7831
rect 17552 7772 18092 7800
rect 19720 7800 19748 7831
rect 19886 7828 19892 7840
rect 19944 7828 19950 7880
rect 20438 7800 20444 7812
rect 19720 7772 20444 7800
rect 17552 7760 17558 7772
rect 19904 7744 19932 7772
rect 20438 7760 20444 7772
rect 20496 7760 20502 7812
rect 10870 7732 10876 7744
rect 5092 7704 10876 7732
rect 4985 7695 5043 7701
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 12250 7692 12256 7744
rect 12308 7732 12314 7744
rect 12618 7732 12624 7744
rect 12308 7704 12624 7732
rect 12308 7692 12314 7704
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 16669 7735 16727 7741
rect 16669 7701 16681 7735
rect 16715 7732 16727 7735
rect 16758 7732 16764 7744
rect 16715 7704 16764 7732
rect 16715 7701 16727 7704
rect 16669 7695 16727 7701
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 19886 7692 19892 7744
rect 19944 7692 19950 7744
rect 20806 7692 20812 7744
rect 20864 7732 20870 7744
rect 21266 7732 21272 7744
rect 20864 7704 21272 7732
rect 20864 7692 20870 7704
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7528 3111 7531
rect 3326 7528 3332 7540
rect 3099 7500 3332 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 4890 7528 4896 7540
rect 4851 7500 4896 7528
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 6822 7528 6828 7540
rect 6783 7500 6828 7528
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 7760 7500 9137 7528
rect 3602 7392 3608 7404
rect 3563 7364 3608 7392
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 6546 7392 6552 7404
rect 5491 7364 6552 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 7374 7392 7380 7404
rect 7335 7364 7380 7392
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 1762 7324 1768 7336
rect 1723 7296 1768 7324
rect 1762 7284 1768 7296
rect 1820 7284 1826 7336
rect 4890 7284 4896 7336
rect 4948 7324 4954 7336
rect 5258 7324 5264 7336
rect 4948 7296 5264 7324
rect 4948 7284 4954 7296
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7324 7343 7327
rect 7760 7324 7788 7500
rect 9125 7497 9137 7500
rect 9171 7528 9183 7531
rect 12618 7528 12624 7540
rect 9171 7500 12624 7528
rect 9171 7497 9183 7500
rect 9125 7491 9183 7497
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 14277 7531 14335 7537
rect 14277 7497 14289 7531
rect 14323 7528 14335 7531
rect 15286 7528 15292 7540
rect 14323 7500 15292 7528
rect 14323 7497 14335 7500
rect 14277 7491 14335 7497
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 16393 7531 16451 7537
rect 16393 7497 16405 7531
rect 16439 7528 16451 7531
rect 16850 7528 16856 7540
rect 16439 7500 16856 7528
rect 16439 7497 16451 7500
rect 16393 7491 16451 7497
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 17218 7488 17224 7540
rect 17276 7528 17282 7540
rect 17276 7500 19012 7528
rect 17276 7488 17282 7500
rect 8478 7420 8484 7472
rect 8536 7460 8542 7472
rect 11238 7460 11244 7472
rect 8536 7432 11244 7460
rect 8536 7420 8542 7432
rect 11238 7420 11244 7432
rect 11296 7420 11302 7472
rect 18874 7460 18880 7472
rect 11440 7432 18880 7460
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 9861 7395 9919 7401
rect 7892 7364 9812 7392
rect 7892 7352 7898 7364
rect 9122 7324 9128 7336
rect 7331 7296 7788 7324
rect 9083 7296 9128 7324
rect 7331 7293 7343 7296
rect 7285 7287 7343 7293
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 9677 7327 9735 7333
rect 9677 7324 9689 7327
rect 9548 7296 9689 7324
rect 9548 7284 9554 7296
rect 9677 7293 9689 7296
rect 9723 7293 9735 7327
rect 9784 7324 9812 7364
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 9950 7392 9956 7404
rect 9907 7364 9956 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 11333 7395 11391 7401
rect 11333 7392 11345 7395
rect 11204 7364 11345 7392
rect 11204 7352 11210 7364
rect 11333 7361 11345 7364
rect 11379 7361 11391 7395
rect 11333 7355 11391 7361
rect 11440 7324 11468 7432
rect 18874 7420 18880 7432
rect 18932 7420 18938 7472
rect 13357 7395 13415 7401
rect 13357 7361 13369 7395
rect 13403 7392 13415 7395
rect 14274 7392 14280 7404
rect 13403 7364 14280 7392
rect 13403 7361 13415 7364
rect 13357 7355 13415 7361
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 14829 7395 14887 7401
rect 14829 7392 14841 7395
rect 14516 7364 14841 7392
rect 14516 7352 14522 7364
rect 14829 7361 14841 7364
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 16574 7352 16580 7404
rect 16632 7392 16638 7404
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 16632 7364 16957 7392
rect 16632 7352 16638 7364
rect 16945 7361 16957 7364
rect 16991 7392 17003 7395
rect 18506 7392 18512 7404
rect 16991 7364 18512 7392
rect 16991 7361 17003 7364
rect 16945 7355 17003 7361
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 9784 7296 11468 7324
rect 13081 7327 13139 7333
rect 9677 7287 9735 7293
rect 13081 7293 13093 7327
rect 13127 7324 13139 7327
rect 13170 7324 13176 7336
rect 13127 7296 13176 7324
rect 13127 7293 13139 7296
rect 13081 7287 13139 7293
rect 13170 7284 13176 7296
rect 13228 7284 13234 7336
rect 13262 7284 13268 7336
rect 13320 7324 13326 7336
rect 13538 7324 13544 7336
rect 13320 7296 13544 7324
rect 13320 7284 13326 7296
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 14645 7327 14703 7333
rect 14645 7293 14657 7327
rect 14691 7324 14703 7327
rect 14918 7324 14924 7336
rect 14691 7296 14924 7324
rect 14691 7293 14703 7296
rect 14645 7287 14703 7293
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 16390 7284 16396 7336
rect 16448 7324 16454 7336
rect 16853 7327 16911 7333
rect 16853 7324 16865 7327
rect 16448 7296 16865 7324
rect 16448 7284 16454 7296
rect 16853 7293 16865 7296
rect 16899 7293 16911 7327
rect 16853 7287 16911 7293
rect 18046 7284 18052 7336
rect 18104 7333 18110 7336
rect 18104 7327 18117 7333
rect 18105 7324 18117 7327
rect 18105 7296 18149 7324
rect 18105 7293 18117 7296
rect 18104 7287 18117 7293
rect 18104 7284 18110 7287
rect 18874 7284 18880 7336
rect 18932 7324 18938 7336
rect 18984 7324 19012 7500
rect 20346 7488 20352 7540
rect 20404 7528 20410 7540
rect 20717 7531 20775 7537
rect 20717 7528 20729 7531
rect 20404 7500 20729 7528
rect 20404 7488 20410 7500
rect 20717 7497 20729 7500
rect 20763 7497 20775 7531
rect 20717 7491 20775 7497
rect 20438 7420 20444 7472
rect 20496 7460 20502 7472
rect 20898 7460 20904 7472
rect 20496 7432 20904 7460
rect 20496 7420 20502 7432
rect 20898 7420 20904 7432
rect 20956 7420 20962 7472
rect 19150 7352 19156 7404
rect 19208 7392 19214 7404
rect 19337 7395 19395 7401
rect 19337 7392 19349 7395
rect 19208 7364 19349 7392
rect 19208 7352 19214 7364
rect 19337 7361 19349 7364
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 18932 7296 19012 7324
rect 19604 7327 19662 7333
rect 18932 7284 18938 7296
rect 19604 7293 19616 7327
rect 19650 7324 19662 7327
rect 20530 7324 20536 7336
rect 19650 7296 20536 7324
rect 19650 7293 19662 7296
rect 19604 7287 19662 7293
rect 20530 7284 20536 7296
rect 20588 7284 20594 7336
rect 2038 7256 2044 7268
rect 1999 7228 2044 7256
rect 2038 7216 2044 7228
rect 2096 7216 2102 7268
rect 3050 7216 3056 7268
rect 3108 7256 3114 7268
rect 3234 7256 3240 7268
rect 3108 7228 3240 7256
rect 3108 7216 3114 7228
rect 3234 7216 3240 7228
rect 3292 7256 3298 7268
rect 3513 7259 3571 7265
rect 3513 7256 3525 7259
rect 3292 7228 3525 7256
rect 3292 7216 3298 7228
rect 3513 7225 3525 7228
rect 3559 7225 3571 7259
rect 11241 7259 11299 7265
rect 11241 7256 11253 7259
rect 3513 7219 3571 7225
rect 9232 7228 11253 7256
rect 1026 7148 1032 7200
rect 1084 7188 1090 7200
rect 1762 7188 1768 7200
rect 1084 7160 1768 7188
rect 1084 7148 1090 7160
rect 1762 7148 1768 7160
rect 1820 7148 1826 7200
rect 2590 7148 2596 7200
rect 2648 7188 2654 7200
rect 3418 7188 3424 7200
rect 2648 7160 3424 7188
rect 2648 7148 2654 7160
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 5258 7188 5264 7200
rect 5219 7160 5264 7188
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 5350 7148 5356 7200
rect 5408 7188 5414 7200
rect 7190 7188 7196 7200
rect 5408 7160 5453 7188
rect 7151 7160 7196 7188
rect 5408 7148 5414 7160
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 9232 7197 9260 7228
rect 11241 7225 11253 7228
rect 11287 7225 11299 7259
rect 11241 7219 11299 7225
rect 11330 7216 11336 7268
rect 11388 7256 11394 7268
rect 11388 7228 15424 7256
rect 11388 7216 11394 7228
rect 9217 7191 9275 7197
rect 9217 7157 9229 7191
rect 9263 7157 9275 7191
rect 9582 7188 9588 7200
rect 9543 7160 9588 7188
rect 9217 7151 9275 7157
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 10781 7191 10839 7197
rect 10781 7157 10793 7191
rect 10827 7188 10839 7191
rect 11054 7188 11060 7200
rect 10827 7160 11060 7188
rect 10827 7157 10839 7160
rect 10781 7151 10839 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11149 7191 11207 7197
rect 11149 7157 11161 7191
rect 11195 7188 11207 7191
rect 11698 7188 11704 7200
rect 11195 7160 11704 7188
rect 11195 7157 11207 7160
rect 11149 7151 11207 7157
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 12710 7188 12716 7200
rect 12671 7160 12716 7188
rect 12710 7148 12716 7160
rect 12768 7148 12774 7200
rect 13173 7191 13231 7197
rect 13173 7157 13185 7191
rect 13219 7188 13231 7191
rect 13354 7188 13360 7200
rect 13219 7160 13360 7188
rect 13219 7157 13231 7160
rect 13173 7151 13231 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 14737 7191 14795 7197
rect 14737 7157 14749 7191
rect 14783 7188 14795 7191
rect 15286 7188 15292 7200
rect 14783 7160 15292 7188
rect 14783 7157 14795 7160
rect 14737 7151 14795 7157
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15396 7188 15424 7228
rect 16574 7216 16580 7268
rect 16632 7256 16638 7268
rect 16761 7259 16819 7265
rect 16761 7256 16773 7259
rect 16632 7228 16773 7256
rect 16632 7216 16638 7228
rect 16761 7225 16773 7228
rect 16807 7225 16819 7259
rect 18325 7259 18383 7265
rect 18325 7256 18337 7259
rect 16761 7219 16819 7225
rect 16868 7228 18337 7256
rect 16868 7188 16896 7228
rect 18325 7225 18337 7228
rect 18371 7225 18383 7259
rect 18325 7219 18383 7225
rect 15396 7160 16896 7188
rect 17954 7148 17960 7200
rect 18012 7188 18018 7200
rect 19886 7188 19892 7200
rect 18012 7160 19892 7188
rect 18012 7148 18018 7160
rect 19886 7148 19892 7160
rect 19944 7148 19950 7200
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 4709 6987 4767 6993
rect 4709 6953 4721 6987
rect 4755 6984 4767 6987
rect 5258 6984 5264 6996
rect 4755 6956 5264 6984
rect 4755 6953 4767 6956
rect 4709 6947 4767 6953
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 7006 6984 7012 6996
rect 6967 6956 7012 6984
rect 7006 6944 7012 6956
rect 7064 6944 7070 6996
rect 7377 6987 7435 6993
rect 7377 6953 7389 6987
rect 7423 6984 7435 6987
rect 8386 6984 8392 6996
rect 7423 6956 7972 6984
rect 7423 6953 7435 6956
rect 7377 6947 7435 6953
rect 5074 6916 5080 6928
rect 5035 6888 5080 6916
rect 5074 6876 5080 6888
rect 5132 6876 5138 6928
rect 6086 6876 6092 6928
rect 6144 6916 6150 6928
rect 7944 6916 7972 6956
rect 8128 6956 8392 6984
rect 8128 6916 8156 6956
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 9582 6944 9588 6996
rect 9640 6944 9646 6996
rect 11057 6987 11115 6993
rect 11057 6953 11069 6987
rect 11103 6984 11115 6987
rect 11146 6984 11152 6996
rect 11103 6956 11152 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 11146 6944 11152 6956
rect 11204 6944 11210 6996
rect 12710 6944 12716 6996
rect 12768 6984 12774 6996
rect 16666 6984 16672 6996
rect 12768 6956 16672 6984
rect 12768 6944 12774 6956
rect 16666 6944 16672 6956
rect 16724 6944 16730 6996
rect 17494 6944 17500 6996
rect 17552 6984 17558 6996
rect 18785 6987 18843 6993
rect 18785 6984 18797 6987
rect 17552 6956 18797 6984
rect 17552 6944 17558 6956
rect 18785 6953 18797 6956
rect 18831 6953 18843 6987
rect 18785 6947 18843 6953
rect 6144 6888 7696 6916
rect 7944 6888 8156 6916
rect 6144 6876 6150 6888
rect 1118 6808 1124 6860
rect 1176 6848 1182 6860
rect 1486 6848 1492 6860
rect 1176 6820 1492 6848
rect 1176 6808 1182 6820
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 2225 6851 2283 6857
rect 2225 6817 2237 6851
rect 2271 6848 2283 6851
rect 2314 6848 2320 6860
rect 2271 6820 2320 6848
rect 2271 6817 2283 6820
rect 2225 6811 2283 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 7466 6848 7472 6860
rect 7427 6820 7472 6848
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7668 6848 7696 6888
rect 8202 6876 8208 6928
rect 8260 6916 8266 6928
rect 9600 6916 9628 6944
rect 8260 6888 9628 6916
rect 8260 6876 8266 6888
rect 14274 6876 14280 6928
rect 14332 6916 14338 6928
rect 16454 6919 16512 6925
rect 16454 6916 16466 6919
rect 14332 6888 16466 6916
rect 14332 6876 14338 6888
rect 16454 6885 16466 6888
rect 16500 6916 16512 6919
rect 16758 6916 16764 6928
rect 16500 6888 16764 6916
rect 16500 6885 16512 6888
rect 16454 6879 16512 6885
rect 16758 6876 16764 6888
rect 16816 6916 16822 6928
rect 17218 6916 17224 6928
rect 16816 6888 17224 6916
rect 16816 6876 16822 6888
rect 17218 6876 17224 6888
rect 17276 6876 17282 6928
rect 18874 6876 18880 6928
rect 18932 6876 18938 6928
rect 8386 6848 8392 6860
rect 7668 6820 8392 6848
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 9030 6808 9036 6860
rect 9088 6848 9094 6860
rect 9766 6848 9772 6860
rect 9088 6820 9772 6848
rect 9088 6808 9094 6820
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 9950 6857 9956 6860
rect 9944 6848 9956 6857
rect 9911 6820 9956 6848
rect 9944 6811 9956 6820
rect 9950 6808 9956 6811
rect 10008 6808 10014 6860
rect 11238 6808 11244 6860
rect 11296 6848 11302 6860
rect 12342 6848 12348 6860
rect 11296 6820 12348 6848
rect 11296 6808 11302 6820
rect 12342 6808 12348 6820
rect 12400 6848 12406 6860
rect 12805 6851 12863 6857
rect 12805 6848 12817 6851
rect 12400 6820 12817 6848
rect 12400 6808 12406 6820
rect 12805 6817 12817 6820
rect 12851 6817 12863 6851
rect 13061 6851 13119 6857
rect 13061 6848 13073 6851
rect 12805 6811 12863 6817
rect 12912 6820 13073 6848
rect 2501 6783 2559 6789
rect 2501 6749 2513 6783
rect 2547 6780 2559 6783
rect 2774 6780 2780 6792
rect 2547 6752 2780 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2774 6740 2780 6752
rect 2832 6740 2838 6792
rect 3418 6740 3424 6792
rect 3476 6780 3482 6792
rect 4706 6780 4712 6792
rect 3476 6752 4712 6780
rect 3476 6740 3482 6752
rect 4706 6740 4712 6752
rect 4764 6780 4770 6792
rect 5169 6783 5227 6789
rect 5169 6780 5181 6783
rect 4764 6752 5181 6780
rect 4764 6740 4770 6752
rect 5169 6749 5181 6752
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 5626 6780 5632 6792
rect 5399 6752 5632 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 5626 6740 5632 6752
rect 5684 6740 5690 6792
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 5644 6712 5672 6740
rect 7374 6712 7380 6724
rect 5644 6684 7380 6712
rect 7374 6672 7380 6684
rect 7432 6712 7438 6724
rect 7576 6712 7604 6743
rect 7432 6684 7604 6712
rect 7432 6672 7438 6684
rect 1210 6604 1216 6656
rect 1268 6644 1274 6656
rect 8202 6644 8208 6656
rect 1268 6616 8208 6644
rect 1268 6604 1274 6616
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8588 6644 8616 6743
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 9306 6780 9312 6792
rect 8812 6752 9312 6780
rect 8812 6740 8818 6752
rect 9306 6740 9312 6752
rect 9364 6780 9370 6792
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9364 6752 9689 6780
rect 9364 6740 9370 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 12912 6780 12940 6820
rect 13061 6817 13073 6820
rect 13107 6817 13119 6851
rect 13061 6811 13119 6817
rect 15838 6808 15844 6860
rect 15896 6848 15902 6860
rect 16209 6851 16267 6857
rect 16209 6848 16221 6851
rect 15896 6820 16221 6848
rect 15896 6808 15902 6820
rect 16209 6817 16221 6820
rect 16255 6817 16267 6851
rect 16209 6811 16267 6817
rect 18506 6808 18512 6860
rect 18564 6848 18570 6860
rect 18892 6848 18920 6876
rect 18564 6820 19012 6848
rect 18564 6808 18570 6820
rect 18984 6789 19012 6820
rect 18877 6783 18935 6789
rect 18877 6780 18889 6783
rect 9677 6743 9735 6749
rect 12820 6752 12940 6780
rect 17788 6752 18889 6780
rect 12710 6672 12716 6724
rect 12768 6712 12774 6724
rect 12820 6712 12848 6752
rect 12768 6684 12848 6712
rect 14185 6715 14243 6721
rect 12768 6672 12774 6684
rect 14185 6681 14197 6715
rect 14231 6712 14243 6715
rect 15194 6712 15200 6724
rect 14231 6684 15200 6712
rect 14231 6681 14243 6684
rect 14185 6675 14243 6681
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 17586 6712 17592 6724
rect 17547 6684 17592 6712
rect 17586 6672 17592 6684
rect 17644 6672 17650 6724
rect 13538 6644 13544 6656
rect 8588 6616 13544 6644
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 14274 6604 14280 6656
rect 14332 6644 14338 6656
rect 17788 6644 17816 6752
rect 18877 6749 18889 6752
rect 18923 6749 18935 6783
rect 18877 6743 18935 6749
rect 18969 6783 19027 6789
rect 18969 6749 18981 6783
rect 19015 6749 19027 6783
rect 18969 6743 19027 6749
rect 17862 6672 17868 6724
rect 17920 6712 17926 6724
rect 18417 6715 18475 6721
rect 18417 6712 18429 6715
rect 17920 6684 18429 6712
rect 17920 6672 17926 6684
rect 18417 6681 18429 6684
rect 18463 6681 18475 6715
rect 18417 6675 18475 6681
rect 18233 6647 18291 6653
rect 18233 6644 18245 6647
rect 14332 6616 18245 6644
rect 14332 6604 14338 6616
rect 18233 6613 18245 6616
rect 18279 6613 18291 6647
rect 18233 6607 18291 6613
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 3421 6443 3479 6449
rect 3421 6409 3433 6443
rect 3467 6440 3479 6443
rect 3786 6440 3792 6452
rect 3467 6412 3792 6440
rect 3467 6409 3479 6412
rect 3421 6403 3479 6409
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 4985 6443 5043 6449
rect 4985 6409 4997 6443
rect 5031 6440 5043 6443
rect 5350 6440 5356 6452
rect 5031 6412 5356 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 7837 6443 7895 6449
rect 7837 6409 7849 6443
rect 7883 6440 7895 6443
rect 10226 6440 10232 6452
rect 7883 6412 10232 6440
rect 7883 6409 7895 6412
rect 7837 6403 7895 6409
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 14369 6443 14427 6449
rect 12492 6412 12537 6440
rect 12492 6400 12498 6412
rect 14369 6409 14381 6443
rect 14415 6440 14427 6443
rect 14642 6440 14648 6452
rect 14415 6412 14648 6440
rect 14415 6409 14427 6412
rect 14369 6403 14427 6409
rect 14642 6400 14648 6412
rect 14700 6400 14706 6452
rect 15838 6400 15844 6452
rect 15896 6440 15902 6452
rect 16393 6443 16451 6449
rect 16393 6440 16405 6443
rect 15896 6412 16405 6440
rect 15896 6400 15902 6412
rect 16393 6409 16405 6412
rect 16439 6409 16451 6443
rect 16393 6403 16451 6409
rect 17770 6400 17776 6452
rect 17828 6440 17834 6452
rect 18417 6443 18475 6449
rect 18417 6440 18429 6443
rect 17828 6412 18429 6440
rect 17828 6400 17834 6412
rect 18417 6409 18429 6412
rect 18463 6409 18475 6443
rect 18417 6403 18475 6409
rect 5810 6372 5816 6384
rect 2240 6344 5816 6372
rect 2240 6313 2268 6344
rect 5810 6332 5816 6344
rect 5868 6332 5874 6384
rect 8386 6372 8392 6384
rect 7116 6344 8392 6372
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 3602 6264 3608 6316
rect 3660 6304 3666 6316
rect 5445 6307 5503 6313
rect 5445 6304 5457 6307
rect 3660 6276 5457 6304
rect 3660 6264 3666 6276
rect 5445 6273 5457 6276
rect 5491 6273 5503 6307
rect 5626 6304 5632 6316
rect 5587 6276 5632 6304
rect 5445 6267 5503 6273
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 1946 6236 1952 6248
rect 1907 6208 1952 6236
rect 1946 6196 1952 6208
rect 2004 6196 2010 6248
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 3237 6239 3295 6245
rect 3237 6236 3249 6239
rect 3016 6208 3249 6236
rect 3016 6196 3022 6208
rect 3237 6205 3249 6208
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 4706 6196 4712 6248
rect 4764 6236 4770 6248
rect 7116 6236 7144 6344
rect 8386 6332 8392 6344
rect 8444 6332 8450 6384
rect 9858 6332 9864 6384
rect 9916 6372 9922 6384
rect 9916 6344 20484 6372
rect 9916 6332 9922 6344
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 12434 6304 12440 6316
rect 7248 6276 8892 6304
rect 7248 6264 7254 6276
rect 7650 6236 7656 6248
rect 4764 6208 7144 6236
rect 7611 6208 7656 6236
rect 4764 6196 4770 6208
rect 7650 6196 7656 6208
rect 7708 6196 7714 6248
rect 8754 6236 8760 6248
rect 8715 6208 8760 6236
rect 8754 6196 8760 6208
rect 8812 6196 8818 6248
rect 8864 6236 8892 6276
rect 10152 6276 12440 6304
rect 10152 6236 10180 6276
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 12710 6264 12716 6316
rect 12768 6304 12774 6316
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12768 6276 13001 6304
rect 12768 6264 12774 6276
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 15013 6307 15071 6313
rect 15013 6273 15025 6307
rect 15059 6304 15071 6307
rect 15194 6304 15200 6316
rect 15059 6276 15200 6304
rect 15059 6273 15071 6276
rect 15013 6267 15071 6273
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17678 6304 17684 6316
rect 17083 6276 17684 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17678 6264 17684 6276
rect 17736 6264 17742 6316
rect 18874 6264 18880 6316
rect 18932 6304 18938 6316
rect 18969 6307 19027 6313
rect 18969 6304 18981 6307
rect 18932 6276 18981 6304
rect 18932 6264 18938 6276
rect 18969 6273 18981 6276
rect 19015 6273 19027 6307
rect 18969 6267 19027 6273
rect 8864 6208 10180 6236
rect 10226 6196 10232 6248
rect 10284 6236 10290 6248
rect 10410 6236 10416 6248
rect 10284 6208 10416 6236
rect 10284 6196 10290 6208
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 10652 6208 10977 6236
rect 10652 6196 10658 6208
rect 10965 6205 10977 6208
rect 11011 6205 11023 6239
rect 10965 6199 11023 6205
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 11112 6208 11652 6236
rect 11112 6196 11118 6208
rect 5350 6168 5356 6180
rect 5263 6140 5356 6168
rect 5350 6128 5356 6140
rect 5408 6168 5414 6180
rect 5534 6168 5540 6180
rect 5408 6140 5540 6168
rect 5408 6128 5414 6140
rect 5534 6128 5540 6140
rect 5592 6128 5598 6180
rect 5626 6128 5632 6180
rect 5684 6168 5690 6180
rect 9030 6177 9036 6180
rect 9024 6168 9036 6177
rect 5684 6140 8791 6168
rect 8991 6140 9036 6168
rect 5684 6128 5690 6140
rect 3786 6060 3792 6112
rect 3844 6100 3850 6112
rect 8294 6100 8300 6112
rect 3844 6072 8300 6100
rect 3844 6060 3850 6072
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 8386 6060 8392 6112
rect 8444 6100 8450 6112
rect 8662 6100 8668 6112
rect 8444 6072 8668 6100
rect 8444 6060 8450 6072
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 8763 6100 8791 6140
rect 9024 6131 9036 6140
rect 9030 6128 9036 6131
rect 9088 6128 9094 6180
rect 9122 6128 9128 6180
rect 9180 6168 9186 6180
rect 11241 6171 11299 6177
rect 11241 6168 11253 6171
rect 9180 6140 11253 6168
rect 9180 6128 9186 6140
rect 11241 6137 11253 6140
rect 11287 6137 11299 6171
rect 11624 6168 11652 6208
rect 13538 6196 13544 6248
rect 13596 6236 13602 6248
rect 14737 6239 14795 6245
rect 14737 6236 14749 6239
rect 13596 6208 14749 6236
rect 13596 6196 13602 6208
rect 14737 6205 14749 6208
rect 14783 6205 14795 6239
rect 14737 6199 14795 6205
rect 15746 6196 15752 6248
rect 15804 6236 15810 6248
rect 16850 6236 16856 6248
rect 15804 6208 16856 6236
rect 15804 6196 15810 6208
rect 16850 6196 16856 6208
rect 16908 6196 16914 6248
rect 18782 6236 18788 6248
rect 18743 6208 18788 6236
rect 18782 6196 18788 6208
rect 18840 6196 18846 6248
rect 19886 6196 19892 6248
rect 19944 6236 19950 6248
rect 20070 6236 20076 6248
rect 19944 6208 20076 6236
rect 19944 6196 19950 6208
rect 20070 6196 20076 6208
rect 20128 6196 20134 6248
rect 20456 6245 20484 6344
rect 20530 6264 20536 6316
rect 20588 6304 20594 6316
rect 20625 6307 20683 6313
rect 20625 6304 20637 6307
rect 20588 6276 20637 6304
rect 20588 6264 20594 6276
rect 20625 6273 20637 6276
rect 20671 6273 20683 6307
rect 20625 6267 20683 6273
rect 20441 6239 20499 6245
rect 20441 6205 20453 6239
rect 20487 6205 20499 6239
rect 20441 6199 20499 6205
rect 12897 6171 12955 6177
rect 12897 6168 12909 6171
rect 11624 6140 12909 6168
rect 11241 6131 11299 6137
rect 12897 6137 12909 6140
rect 12943 6137 12955 6171
rect 12897 6131 12955 6137
rect 15930 6128 15936 6180
rect 15988 6168 15994 6180
rect 17402 6168 17408 6180
rect 15988 6140 17408 6168
rect 15988 6128 15994 6140
rect 17402 6128 17408 6140
rect 17460 6128 17466 6180
rect 17494 6128 17500 6180
rect 17552 6168 17558 6180
rect 18874 6168 18880 6180
rect 17552 6140 18880 6168
rect 17552 6128 17558 6140
rect 18874 6128 18880 6140
rect 18932 6128 18938 6180
rect 9858 6100 9864 6112
rect 8763 6072 9864 6100
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 9950 6060 9956 6112
rect 10008 6100 10014 6112
rect 10137 6103 10195 6109
rect 10137 6100 10149 6103
rect 10008 6072 10149 6100
rect 10008 6060 10014 6072
rect 10137 6069 10149 6072
rect 10183 6100 10195 6103
rect 10410 6100 10416 6112
rect 10183 6072 10416 6100
rect 10183 6069 10195 6072
rect 10137 6063 10195 6069
rect 10410 6060 10416 6072
rect 10468 6060 10474 6112
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 11112 6072 12817 6100
rect 11112 6060 11118 6072
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 12805 6063 12863 6069
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 13872 6072 14841 6100
rect 13872 6060 13878 6072
rect 14829 6069 14841 6072
rect 14875 6069 14887 6103
rect 16758 6100 16764 6112
rect 16719 6072 16764 6100
rect 14829 6063 14887 6069
rect 16758 6060 16764 6072
rect 16816 6060 16822 6112
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 16908 6072 16953 6100
rect 16908 6060 16914 6072
rect 18782 6060 18788 6112
rect 18840 6100 18846 6112
rect 19150 6100 19156 6112
rect 18840 6072 19156 6100
rect 18840 6060 18846 6072
rect 19150 6060 19156 6072
rect 19208 6060 19214 6112
rect 20070 6100 20076 6112
rect 20031 6072 20076 6100
rect 20070 6060 20076 6072
rect 20128 6060 20134 6112
rect 20530 6060 20536 6112
rect 20588 6100 20594 6112
rect 20588 6072 20633 6100
rect 20588 6060 20594 6072
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 1949 5899 2007 5905
rect 1949 5865 1961 5899
rect 1995 5896 2007 5899
rect 2866 5896 2872 5908
rect 1995 5868 2872 5896
rect 1995 5865 2007 5868
rect 1949 5859 2007 5865
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3053 5899 3111 5905
rect 3053 5865 3065 5899
rect 3099 5896 3111 5899
rect 3510 5896 3516 5908
rect 3099 5868 3516 5896
rect 3099 5865 3111 5868
rect 3053 5859 3111 5865
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 4249 5899 4307 5905
rect 4249 5865 4261 5899
rect 4295 5896 4307 5899
rect 4338 5896 4344 5908
rect 4295 5868 4344 5896
rect 4295 5865 4307 5868
rect 4249 5859 4307 5865
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 5224 5868 5365 5896
rect 5224 5856 5230 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 6454 5896 6460 5908
rect 6415 5868 6460 5896
rect 5353 5859 5411 5865
rect 6454 5856 6460 5868
rect 6512 5856 6518 5908
rect 8662 5896 8668 5908
rect 7392 5868 8668 5896
rect 7190 5828 7196 5840
rect 5184 5800 7196 5828
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 2038 5760 2044 5772
rect 1811 5732 2044 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 2038 5720 2044 5732
rect 2096 5720 2102 5772
rect 2869 5763 2927 5769
rect 2869 5729 2881 5763
rect 2915 5729 2927 5763
rect 2869 5723 2927 5729
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 4706 5760 4712 5772
rect 4111 5732 4712 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 2884 5624 2912 5723
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 5184 5769 5212 5800
rect 7190 5788 7196 5800
rect 7248 5788 7254 5840
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5729 5227 5763
rect 5169 5723 5227 5729
rect 6273 5763 6331 5769
rect 6273 5729 6285 5763
rect 6319 5760 6331 5763
rect 6362 5760 6368 5772
rect 6319 5732 6368 5760
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 6362 5720 6368 5732
rect 6420 5720 6426 5772
rect 7392 5769 7420 5868
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 9677 5899 9735 5905
rect 9677 5896 9689 5899
rect 8763 5868 9689 5896
rect 8763 5828 8791 5868
rect 9677 5865 9689 5868
rect 9723 5865 9735 5899
rect 9677 5859 9735 5865
rect 9769 5899 9827 5905
rect 9769 5865 9781 5899
rect 9815 5896 9827 5899
rect 10686 5896 10692 5908
rect 9815 5868 10692 5896
rect 9815 5865 9827 5868
rect 9769 5859 9827 5865
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 12710 5896 12716 5908
rect 11440 5868 12572 5896
rect 12671 5868 12716 5896
rect 7484 5800 8791 5828
rect 7383 5763 7441 5769
rect 7383 5729 7395 5763
rect 7429 5729 7441 5763
rect 7383 5723 7441 5729
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 7484 5692 7512 5800
rect 9306 5788 9312 5840
rect 9364 5828 9370 5840
rect 9364 5800 11100 5828
rect 9364 5788 9370 5800
rect 8478 5760 8484 5772
rect 8439 5732 8484 5760
rect 8478 5720 8484 5732
rect 8536 5720 8542 5772
rect 8662 5720 8668 5772
rect 8720 5760 8726 5772
rect 9122 5760 9128 5772
rect 8720 5732 9128 5760
rect 8720 5720 8726 5732
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 10137 5763 10195 5769
rect 10137 5760 10149 5763
rect 9723 5732 10149 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 10137 5729 10149 5732
rect 10183 5729 10195 5763
rect 11072 5760 11100 5800
rect 11146 5788 11152 5840
rect 11204 5828 11210 5840
rect 11440 5828 11468 5868
rect 11204 5800 11468 5828
rect 11204 5788 11210 5800
rect 11514 5788 11520 5840
rect 11572 5837 11578 5840
rect 11572 5831 11636 5837
rect 11572 5797 11590 5831
rect 11624 5797 11636 5831
rect 12544 5828 12572 5868
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 13538 5896 13544 5908
rect 13499 5868 13544 5896
rect 13538 5856 13544 5868
rect 13596 5896 13602 5908
rect 14001 5899 14059 5905
rect 14001 5896 14013 5899
rect 13596 5868 14013 5896
rect 13596 5856 13602 5868
rect 14001 5865 14013 5868
rect 14047 5865 14059 5899
rect 14001 5859 14059 5865
rect 14093 5899 14151 5905
rect 14093 5865 14105 5899
rect 14139 5896 14151 5899
rect 14642 5896 14648 5908
rect 14139 5868 14648 5896
rect 14139 5865 14151 5868
rect 14093 5859 14151 5865
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 15286 5896 15292 5908
rect 15247 5868 15292 5896
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 16758 5856 16764 5908
rect 16816 5896 16822 5908
rect 17497 5899 17555 5905
rect 17497 5896 17509 5899
rect 16816 5868 17509 5896
rect 16816 5856 16822 5868
rect 17497 5865 17509 5868
rect 17543 5865 17555 5899
rect 17497 5859 17555 5865
rect 17957 5899 18015 5905
rect 17957 5865 17969 5899
rect 18003 5896 18015 5899
rect 19061 5899 19119 5905
rect 19061 5896 19073 5899
rect 18003 5868 19073 5896
rect 18003 5865 18015 5868
rect 17957 5859 18015 5865
rect 19061 5865 19073 5868
rect 19107 5865 19119 5899
rect 19061 5859 19119 5865
rect 19242 5856 19248 5908
rect 19300 5896 19306 5908
rect 19429 5899 19487 5905
rect 19429 5896 19441 5899
rect 19300 5868 19441 5896
rect 19300 5856 19306 5868
rect 19429 5865 19441 5868
rect 19475 5865 19487 5899
rect 19429 5859 19487 5865
rect 19150 5828 19156 5840
rect 12544 5800 19156 5828
rect 11572 5791 11636 5797
rect 11572 5788 11578 5791
rect 19150 5788 19156 5800
rect 19208 5828 19214 5840
rect 19521 5831 19579 5837
rect 19521 5828 19533 5831
rect 19208 5800 19533 5828
rect 19208 5788 19214 5800
rect 19521 5797 19533 5800
rect 19567 5797 19579 5831
rect 19521 5791 19579 5797
rect 11072 5732 12388 5760
rect 10137 5723 10195 5729
rect 3752 5664 7512 5692
rect 7576 5664 8791 5692
rect 3752 5652 3758 5664
rect 6086 5624 6092 5636
rect 2884 5596 6092 5624
rect 6086 5584 6092 5596
rect 6144 5584 6150 5636
rect 7576 5633 7604 5664
rect 7561 5627 7619 5633
rect 7561 5593 7573 5627
rect 7607 5593 7619 5627
rect 8763 5624 8791 5664
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 9364 5664 10180 5692
rect 9364 5652 9370 5664
rect 10152 5624 10180 5664
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10410 5692 10416 5704
rect 10284 5664 10329 5692
rect 10371 5664 10416 5692
rect 10284 5652 10290 5664
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 11330 5692 11336 5704
rect 11291 5664 11336 5692
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 11146 5624 11152 5636
rect 8763 5596 10088 5624
rect 10152 5596 11152 5624
rect 7561 5587 7619 5593
rect 6638 5516 6644 5568
rect 6696 5556 6702 5568
rect 8018 5556 8024 5568
rect 6696 5528 8024 5556
rect 6696 5516 6702 5528
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 8662 5556 8668 5568
rect 8623 5528 8668 5556
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 9122 5516 9128 5568
rect 9180 5556 9186 5568
rect 9858 5556 9864 5568
rect 9180 5528 9864 5556
rect 9180 5516 9186 5528
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 10060 5556 10088 5596
rect 11146 5584 11152 5596
rect 11204 5584 11210 5636
rect 12360 5624 12388 5732
rect 12618 5720 12624 5772
rect 12676 5760 12682 5772
rect 15654 5760 15660 5772
rect 12676 5732 15660 5760
rect 12676 5720 12682 5732
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 15749 5763 15807 5769
rect 15749 5729 15761 5763
rect 15795 5760 15807 5763
rect 17770 5760 17776 5772
rect 15795 5732 17776 5760
rect 15795 5729 15807 5732
rect 15749 5723 15807 5729
rect 17770 5720 17776 5732
rect 17828 5720 17834 5772
rect 17865 5763 17923 5769
rect 17865 5729 17877 5763
rect 17911 5760 17923 5763
rect 17954 5760 17960 5772
rect 17911 5732 17960 5760
rect 17911 5729 17923 5732
rect 17865 5723 17923 5729
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5692 14335 5695
rect 14366 5692 14372 5704
rect 14323 5664 14372 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 14366 5652 14372 5664
rect 14424 5652 14430 5704
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 15841 5695 15899 5701
rect 15841 5692 15853 5695
rect 15252 5664 15853 5692
rect 15252 5652 15258 5664
rect 15841 5661 15853 5664
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 17586 5652 17592 5704
rect 17644 5692 17650 5704
rect 18049 5695 18107 5701
rect 18049 5692 18061 5695
rect 17644 5664 18061 5692
rect 17644 5652 17650 5664
rect 18049 5661 18061 5664
rect 18095 5661 18107 5695
rect 18049 5655 18107 5661
rect 18874 5652 18880 5704
rect 18932 5692 18938 5704
rect 19613 5695 19671 5701
rect 19613 5692 19625 5695
rect 18932 5664 19625 5692
rect 18932 5652 18938 5664
rect 19613 5661 19625 5664
rect 19659 5661 19671 5695
rect 19613 5655 19671 5661
rect 13633 5627 13691 5633
rect 13633 5624 13645 5627
rect 12360 5596 13645 5624
rect 13633 5593 13645 5596
rect 13679 5593 13691 5627
rect 13633 5587 13691 5593
rect 10778 5556 10784 5568
rect 10060 5528 10784 5556
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 18966 5556 18972 5568
rect 13596 5528 18972 5556
rect 13596 5516 13602 5528
rect 18966 5516 18972 5528
rect 19024 5516 19030 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 1578 5312 1584 5364
rect 1636 5352 1642 5364
rect 1949 5355 2007 5361
rect 1949 5352 1961 5355
rect 1636 5324 1961 5352
rect 1636 5312 1642 5324
rect 1949 5321 1961 5324
rect 1995 5321 2007 5355
rect 1949 5315 2007 5321
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3142 5352 3148 5364
rect 3099 5324 3148 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3142 5312 3148 5324
rect 3200 5312 3206 5364
rect 4154 5352 4160 5364
rect 4115 5324 4160 5352
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 5261 5355 5319 5361
rect 5261 5321 5273 5355
rect 5307 5352 5319 5355
rect 5442 5352 5448 5364
rect 5307 5324 5448 5352
rect 5307 5321 5319 5324
rect 5261 5315 5319 5321
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5352 7159 5355
rect 7558 5352 7564 5364
rect 7147 5324 7564 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7558 5312 7564 5324
rect 7616 5312 7622 5364
rect 8202 5352 8208 5364
rect 8163 5324 8208 5352
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 9125 5355 9183 5361
rect 9125 5321 9137 5355
rect 9171 5352 9183 5355
rect 9490 5352 9496 5364
rect 9171 5324 9496 5352
rect 9171 5321 9183 5324
rect 9125 5315 9183 5321
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 10781 5355 10839 5361
rect 10781 5321 10793 5355
rect 10827 5352 10839 5355
rect 11054 5352 11060 5364
rect 10827 5324 11060 5352
rect 10827 5321 10839 5324
rect 10781 5315 10839 5321
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11698 5312 11704 5364
rect 11756 5352 11762 5364
rect 12437 5355 12495 5361
rect 12437 5352 12449 5355
rect 11756 5324 12449 5352
rect 11756 5312 11762 5324
rect 12437 5321 12449 5324
rect 12483 5321 12495 5355
rect 12437 5315 12495 5321
rect 14001 5355 14059 5361
rect 14001 5321 14013 5355
rect 14047 5352 14059 5355
rect 14182 5352 14188 5364
rect 14047 5324 14188 5352
rect 14047 5321 14059 5324
rect 14001 5315 14059 5321
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 16393 5355 16451 5361
rect 16393 5321 16405 5355
rect 16439 5352 16451 5355
rect 16850 5352 16856 5364
rect 16439 5324 16856 5352
rect 16439 5321 16451 5324
rect 16393 5315 16451 5321
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 18049 5355 18107 5361
rect 18049 5352 18061 5355
rect 18012 5324 18061 5352
rect 18012 5312 18018 5324
rect 18049 5321 18061 5324
rect 18095 5321 18107 5355
rect 18049 5315 18107 5321
rect 19981 5355 20039 5361
rect 19981 5321 19993 5355
rect 20027 5352 20039 5355
rect 20254 5352 20260 5364
rect 20027 5324 20260 5352
rect 20027 5321 20039 5324
rect 19981 5315 20039 5321
rect 20254 5312 20260 5324
rect 20312 5312 20318 5364
rect 9306 5284 9312 5296
rect 7116 5256 9312 5284
rect 7116 5228 7144 5256
rect 9306 5244 9312 5256
rect 9364 5244 9370 5296
rect 10318 5244 10324 5296
rect 10376 5284 10382 5296
rect 10376 5256 16896 5284
rect 10376 5244 10382 5256
rect 7098 5216 7104 5228
rect 1780 5188 7104 5216
rect 1780 5157 1808 5188
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 8570 5176 8576 5228
rect 8628 5216 8634 5228
rect 9030 5216 9036 5228
rect 8628 5188 9036 5216
rect 8628 5176 8634 5188
rect 9030 5176 9036 5188
rect 9088 5216 9094 5228
rect 9677 5219 9735 5225
rect 9677 5216 9689 5219
rect 9088 5188 9689 5216
rect 9088 5176 9094 5188
rect 9677 5185 9689 5188
rect 9723 5185 9735 5219
rect 9677 5179 9735 5185
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 11241 5219 11299 5225
rect 11241 5216 11253 5219
rect 10744 5188 11253 5216
rect 10744 5176 10750 5188
rect 11241 5185 11253 5188
rect 11287 5185 11299 5219
rect 11241 5179 11299 5185
rect 11330 5176 11336 5228
rect 11388 5216 11394 5228
rect 11388 5188 11433 5216
rect 11388 5176 11394 5188
rect 11698 5176 11704 5228
rect 11756 5216 11762 5228
rect 12989 5219 13047 5225
rect 12989 5216 13001 5219
rect 11756 5188 13001 5216
rect 11756 5176 11762 5188
rect 12989 5185 13001 5188
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 14366 5176 14372 5228
rect 14424 5216 14430 5228
rect 14553 5219 14611 5225
rect 14553 5216 14565 5219
rect 14424 5188 14565 5216
rect 14424 5176 14430 5188
rect 14553 5185 14565 5188
rect 14599 5185 14611 5219
rect 14553 5179 14611 5185
rect 16666 5176 16672 5228
rect 16724 5216 16730 5228
rect 16724 5188 16804 5216
rect 16724 5176 16730 5188
rect 1771 5151 1829 5157
rect 1771 5117 1783 5151
rect 1817 5117 1829 5151
rect 2866 5148 2872 5160
rect 2827 5120 2872 5148
rect 1771 5111 1829 5117
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 3973 5151 4031 5157
rect 3973 5117 3985 5151
rect 4019 5148 4031 5151
rect 4154 5148 4160 5160
rect 4019 5120 4160 5148
rect 4019 5117 4031 5120
rect 3973 5111 4031 5117
rect 4154 5108 4160 5120
rect 4212 5108 4218 5160
rect 4982 5108 4988 5160
rect 5040 5148 5046 5160
rect 5077 5151 5135 5157
rect 5077 5148 5089 5151
rect 5040 5120 5089 5148
rect 5040 5108 5046 5120
rect 5077 5117 5089 5120
rect 5123 5117 5135 5151
rect 5077 5111 5135 5117
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5117 6975 5151
rect 8018 5148 8024 5160
rect 7979 5120 8024 5148
rect 6917 5111 6975 5117
rect 6932 5080 6960 5111
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 9585 5151 9643 5157
rect 9585 5117 9597 5151
rect 9631 5148 9643 5151
rect 12618 5148 12624 5160
rect 9631 5120 12624 5148
rect 9631 5117 9643 5120
rect 9585 5111 9643 5117
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 13170 5148 13176 5160
rect 12943 5120 13176 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 13170 5108 13176 5120
rect 13228 5108 13234 5160
rect 13998 5108 14004 5160
rect 14056 5148 14062 5160
rect 16776 5157 16804 5188
rect 14461 5151 14519 5157
rect 14461 5148 14473 5151
rect 14056 5120 14473 5148
rect 14056 5108 14062 5120
rect 14461 5117 14473 5120
rect 14507 5117 14519 5151
rect 14461 5111 14519 5117
rect 16761 5151 16819 5157
rect 16761 5117 16773 5151
rect 16807 5117 16819 5151
rect 16868 5148 16896 5256
rect 17218 5244 17224 5296
rect 17276 5284 17282 5296
rect 18874 5284 18880 5296
rect 17276 5256 18880 5284
rect 17276 5244 17282 5256
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5216 17095 5219
rect 17586 5216 17592 5228
rect 17083 5188 17592 5216
rect 17083 5185 17095 5188
rect 17037 5179 17095 5185
rect 17586 5176 17592 5188
rect 17644 5176 17650 5228
rect 18616 5225 18644 5256
rect 18874 5244 18880 5256
rect 18932 5244 18938 5296
rect 20346 5244 20352 5296
rect 20404 5284 20410 5296
rect 20404 5256 20576 5284
rect 20404 5244 20410 5256
rect 18601 5219 18659 5225
rect 18601 5185 18613 5219
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 20070 5176 20076 5228
rect 20128 5216 20134 5228
rect 20548 5225 20576 5256
rect 20441 5219 20499 5225
rect 20441 5216 20453 5219
rect 20128 5188 20453 5216
rect 20128 5176 20134 5188
rect 20441 5185 20453 5188
rect 20487 5185 20499 5219
rect 20441 5179 20499 5185
rect 20533 5219 20591 5225
rect 20533 5185 20545 5219
rect 20579 5185 20591 5219
rect 20533 5179 20591 5185
rect 20349 5151 20407 5157
rect 20349 5148 20361 5151
rect 16868 5120 20361 5148
rect 16761 5111 16819 5117
rect 20349 5117 20361 5120
rect 20395 5117 20407 5151
rect 20349 5111 20407 5117
rect 9306 5080 9312 5092
rect 6932 5052 9312 5080
rect 9306 5040 9312 5052
rect 9364 5040 9370 5092
rect 9493 5083 9551 5089
rect 9493 5049 9505 5083
rect 9539 5080 9551 5083
rect 9766 5080 9772 5092
rect 9539 5052 9772 5080
rect 9539 5049 9551 5052
rect 9493 5043 9551 5049
rect 9766 5040 9772 5052
rect 9824 5040 9830 5092
rect 12434 5080 12440 5092
rect 10980 5052 12440 5080
rect 8202 4972 8208 5024
rect 8260 5012 8266 5024
rect 10980 5012 11008 5052
rect 12434 5040 12440 5052
rect 12492 5040 12498 5092
rect 18417 5083 18475 5089
rect 18417 5080 18429 5083
rect 12544 5052 18429 5080
rect 8260 4984 11008 5012
rect 8260 4972 8266 4984
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 11149 5015 11207 5021
rect 11149 5012 11161 5015
rect 11112 4984 11161 5012
rect 11112 4972 11118 4984
rect 11149 4981 11161 4984
rect 11195 4981 11207 5015
rect 11149 4975 11207 4981
rect 12342 4972 12348 5024
rect 12400 5012 12406 5024
rect 12544 5012 12572 5052
rect 18417 5049 18429 5052
rect 18463 5049 18475 5083
rect 18417 5043 18475 5049
rect 12400 4984 12572 5012
rect 12805 5015 12863 5021
rect 12400 4972 12406 4984
rect 12805 4981 12817 5015
rect 12851 5012 12863 5015
rect 14182 5012 14188 5024
rect 12851 4984 14188 5012
rect 12851 4981 12863 4984
rect 12805 4975 12863 4981
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 14274 4972 14280 5024
rect 14332 5012 14338 5024
rect 14369 5015 14427 5021
rect 14369 5012 14381 5015
rect 14332 4984 14381 5012
rect 14332 4972 14338 4984
rect 14369 4981 14381 4984
rect 14415 4981 14427 5015
rect 14369 4975 14427 4981
rect 16850 4972 16856 5024
rect 16908 5012 16914 5024
rect 16908 4984 16953 5012
rect 16908 4972 16914 4984
rect 17126 4972 17132 5024
rect 17184 5012 17190 5024
rect 18509 5015 18567 5021
rect 18509 5012 18521 5015
rect 17184 4984 18521 5012
rect 17184 4972 17190 4984
rect 18509 4981 18521 4984
rect 18555 4981 18567 5015
rect 18509 4975 18567 4981
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 1949 4811 2007 4817
rect 1949 4808 1961 4811
rect 1728 4780 1961 4808
rect 1728 4768 1734 4780
rect 1949 4777 1961 4780
rect 1995 4777 2007 4811
rect 1949 4771 2007 4777
rect 4249 4811 4307 4817
rect 4249 4777 4261 4811
rect 4295 4808 4307 4811
rect 4798 4808 4804 4820
rect 4295 4780 4804 4808
rect 4295 4777 4307 4780
rect 4249 4771 4307 4777
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 5994 4768 6000 4820
rect 6052 4808 6058 4820
rect 6365 4811 6423 4817
rect 6365 4808 6377 4811
rect 6052 4780 6377 4808
rect 6052 4768 6058 4780
rect 6365 4777 6377 4780
rect 6411 4777 6423 4811
rect 6365 4771 6423 4777
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 7742 4808 7748 4820
rect 7607 4780 7748 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 8386 4768 8392 4820
rect 8444 4808 8450 4820
rect 8665 4811 8723 4817
rect 8665 4808 8677 4811
rect 8444 4780 8677 4808
rect 8444 4768 8450 4780
rect 8665 4777 8677 4780
rect 8711 4777 8723 4811
rect 8665 4771 8723 4777
rect 10137 4811 10195 4817
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10318 4808 10324 4820
rect 10183 4780 10324 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10318 4768 10324 4780
rect 10376 4768 10382 4820
rect 11054 4808 11060 4820
rect 11015 4780 11060 4808
rect 11054 4768 11060 4780
rect 11112 4768 11118 4820
rect 11514 4808 11520 4820
rect 11427 4780 11520 4808
rect 11514 4768 11520 4780
rect 11572 4808 11578 4820
rect 11572 4780 11744 4808
rect 11572 4768 11578 4780
rect 3970 4700 3976 4752
rect 4028 4740 4034 4752
rect 11716 4740 11744 4780
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 12621 4811 12679 4817
rect 12621 4808 12633 4811
rect 12400 4780 12633 4808
rect 12400 4768 12406 4780
rect 12621 4777 12633 4780
rect 12667 4777 12679 4811
rect 13446 4808 13452 4820
rect 12621 4771 12679 4777
rect 12820 4780 13452 4808
rect 12820 4740 12848 4780
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 14001 4811 14059 4817
rect 14001 4777 14013 4811
rect 14047 4808 14059 4811
rect 14642 4808 14648 4820
rect 14047 4780 14648 4808
rect 14047 4777 14059 4780
rect 14001 4771 14059 4777
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 15470 4808 15476 4820
rect 15431 4780 15476 4808
rect 15470 4768 15476 4780
rect 15528 4768 15534 4820
rect 16485 4811 16543 4817
rect 16485 4777 16497 4811
rect 16531 4808 16543 4811
rect 16850 4808 16856 4820
rect 16531 4780 16856 4808
rect 16531 4777 16543 4780
rect 16485 4771 16543 4777
rect 16850 4768 16856 4780
rect 16908 4768 16914 4820
rect 18509 4811 18567 4817
rect 18509 4777 18521 4811
rect 18555 4808 18567 4811
rect 18782 4808 18788 4820
rect 18555 4780 18788 4808
rect 18555 4777 18567 4780
rect 18509 4771 18567 4777
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 19889 4811 19947 4817
rect 19889 4808 19901 4811
rect 19392 4780 19901 4808
rect 19392 4768 19398 4780
rect 19889 4777 19901 4780
rect 19935 4777 19947 4811
rect 19889 4771 19947 4777
rect 4028 4712 5212 4740
rect 11716 4712 12848 4740
rect 4028 4700 4034 4712
rect 1765 4675 1823 4681
rect 1765 4641 1777 4675
rect 1811 4672 1823 4675
rect 1854 4672 1860 4684
rect 1811 4644 1860 4672
rect 1811 4641 1823 4644
rect 1765 4635 1823 4641
rect 1854 4632 1860 4644
rect 1912 4632 1918 4684
rect 2869 4675 2927 4681
rect 2869 4641 2881 4675
rect 2915 4672 2927 4675
rect 3326 4672 3332 4684
rect 2915 4644 3332 4672
rect 2915 4641 2927 4644
rect 2869 4635 2927 4641
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 4065 4675 4123 4681
rect 4065 4641 4077 4675
rect 4111 4672 4123 4675
rect 4246 4672 4252 4684
rect 4111 4644 4252 4672
rect 4111 4641 4123 4644
rect 4065 4635 4123 4641
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 5184 4681 5212 4712
rect 13354 4700 13360 4752
rect 13412 4740 13418 4752
rect 14093 4743 14151 4749
rect 14093 4740 14105 4743
rect 13412 4712 14105 4740
rect 13412 4700 13418 4712
rect 14093 4709 14105 4712
rect 14139 4709 14151 4743
rect 14093 4703 14151 4709
rect 14182 4700 14188 4752
rect 14240 4740 14246 4752
rect 16666 4740 16672 4752
rect 14240 4712 16672 4740
rect 14240 4700 14246 4712
rect 16666 4700 16672 4712
rect 16724 4700 16730 4752
rect 16945 4743 17003 4749
rect 16945 4740 16957 4743
rect 16767 4712 16957 4740
rect 5169 4675 5227 4681
rect 5169 4641 5181 4675
rect 5215 4641 5227 4675
rect 5169 4635 5227 4641
rect 7377 4675 7435 4681
rect 7377 4641 7389 4675
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4672 8539 4675
rect 9398 4672 9404 4684
rect 8527 4644 9404 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 3970 4564 3976 4616
rect 4028 4604 4034 4616
rect 7392 4604 7420 4635
rect 9398 4632 9404 4644
rect 9456 4632 9462 4684
rect 9950 4672 9956 4684
rect 9911 4644 9956 4672
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 11054 4632 11060 4684
rect 11112 4672 11118 4684
rect 11425 4675 11483 4681
rect 11425 4672 11437 4675
rect 11112 4644 11437 4672
rect 11112 4632 11118 4644
rect 11425 4641 11437 4644
rect 11471 4641 11483 4675
rect 15289 4675 15347 4681
rect 11425 4635 11483 4641
rect 12360 4644 14688 4672
rect 11514 4604 11520 4616
rect 4028 4576 11520 4604
rect 4028 4564 4034 4576
rect 11514 4564 11520 4576
rect 11572 4564 11578 4616
rect 11698 4604 11704 4616
rect 11659 4576 11704 4604
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 14 4496 20 4548
rect 72 4536 78 4548
rect 3053 4539 3111 4545
rect 3053 4536 3065 4539
rect 72 4508 3065 4536
rect 72 4496 78 4508
rect 3053 4505 3065 4508
rect 3099 4505 3111 4539
rect 3053 4499 3111 4505
rect 5353 4539 5411 4545
rect 5353 4505 5365 4539
rect 5399 4536 5411 4539
rect 12360 4536 12388 4644
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 14550 4604 14556 4616
rect 14323 4576 14556 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 14550 4564 14556 4576
rect 14608 4564 14614 4616
rect 14660 4604 14688 4644
rect 15289 4641 15301 4675
rect 15335 4672 15347 4675
rect 15378 4672 15384 4684
rect 15335 4644 15384 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 15378 4632 15384 4644
rect 15436 4632 15442 4684
rect 16390 4632 16396 4684
rect 16448 4672 16454 4684
rect 16767 4672 16795 4712
rect 16945 4709 16957 4712
rect 16991 4740 17003 4743
rect 17678 4740 17684 4752
rect 16991 4712 17684 4740
rect 16991 4709 17003 4712
rect 16945 4703 17003 4709
rect 17678 4700 17684 4712
rect 17736 4700 17742 4752
rect 18138 4700 18144 4752
rect 18196 4740 18202 4752
rect 18196 4712 18736 4740
rect 18196 4700 18202 4712
rect 16448 4644 16795 4672
rect 16448 4632 16454 4644
rect 16850 4632 16856 4684
rect 16908 4672 16914 4684
rect 17494 4672 17500 4684
rect 16908 4644 16953 4672
rect 17052 4644 17500 4672
rect 16908 4632 16914 4644
rect 17052 4604 17080 4644
rect 17494 4632 17500 4644
rect 17552 4632 17558 4684
rect 17586 4632 17592 4684
rect 17644 4672 17650 4684
rect 18601 4675 18659 4681
rect 18601 4672 18613 4675
rect 17644 4644 18613 4672
rect 17644 4632 17650 4644
rect 18601 4641 18613 4644
rect 18647 4641 18659 4675
rect 18601 4635 18659 4641
rect 14660 4576 17080 4604
rect 17129 4607 17187 4613
rect 17129 4573 17141 4607
rect 17175 4604 17187 4607
rect 17218 4604 17224 4616
rect 17175 4576 17224 4604
rect 17175 4573 17187 4576
rect 17129 4567 17187 4573
rect 17218 4564 17224 4576
rect 17276 4564 17282 4616
rect 18708 4613 18736 4712
rect 19518 4700 19524 4752
rect 19576 4740 19582 4752
rect 20254 4740 20260 4752
rect 19576 4712 20260 4740
rect 19576 4700 19582 4712
rect 20254 4700 20260 4712
rect 20312 4700 20318 4752
rect 19426 4632 19432 4684
rect 19484 4672 19490 4684
rect 19705 4675 19763 4681
rect 19705 4672 19717 4675
rect 19484 4644 19717 4672
rect 19484 4632 19490 4644
rect 19705 4641 19717 4644
rect 19751 4641 19763 4675
rect 19705 4635 19763 4641
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4573 18751 4607
rect 18693 4567 18751 4573
rect 19518 4564 19524 4616
rect 19576 4604 19582 4616
rect 20714 4604 20720 4616
rect 19576 4576 20720 4604
rect 19576 4564 19582 4576
rect 20714 4564 20720 4576
rect 20772 4564 20778 4616
rect 5399 4508 12388 4536
rect 5399 4505 5411 4508
rect 5353 4499 5411 4505
rect 12434 4496 12440 4548
rect 12492 4536 12498 4548
rect 18782 4536 18788 4548
rect 12492 4508 18788 4536
rect 12492 4496 12498 4508
rect 18782 4496 18788 4508
rect 18840 4496 18846 4548
rect 3786 4428 3792 4480
rect 3844 4468 3850 4480
rect 9030 4468 9036 4480
rect 3844 4440 9036 4468
rect 3844 4428 3850 4440
rect 9030 4428 9036 4440
rect 9088 4468 9094 4480
rect 9582 4468 9588 4480
rect 9088 4440 9588 4468
rect 9088 4428 9094 4440
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 14274 4428 14280 4480
rect 14332 4468 14338 4480
rect 17126 4468 17132 4480
rect 14332 4440 17132 4468
rect 14332 4428 14338 4440
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 18141 4471 18199 4477
rect 18141 4437 18153 4471
rect 18187 4468 18199 4471
rect 19610 4468 19616 4480
rect 18187 4440 19616 4468
rect 18187 4437 18199 4440
rect 18141 4431 18199 4437
rect 19610 4428 19616 4440
rect 19668 4428 19674 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 10042 4264 10048 4276
rect 7852 4236 10048 4264
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 4798 4128 4804 4140
rect 1544 4100 4804 4128
rect 1544 4088 1550 4100
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 5074 4128 5080 4140
rect 5035 4100 5080 4128
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 6917 4131 6975 4137
rect 6917 4097 6929 4131
rect 6963 4128 6975 4131
rect 7852 4128 7880 4236
rect 10042 4224 10048 4236
rect 10100 4224 10106 4276
rect 10318 4264 10324 4276
rect 10279 4236 10324 4264
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 12342 4224 12348 4276
rect 12400 4264 12406 4276
rect 15194 4264 15200 4276
rect 12400 4236 15200 4264
rect 12400 4224 12406 4236
rect 15194 4224 15200 4236
rect 15252 4224 15258 4276
rect 16850 4224 16856 4276
rect 16908 4264 16914 4276
rect 17126 4264 17132 4276
rect 16908 4236 17132 4264
rect 16908 4224 16914 4236
rect 17126 4224 17132 4236
rect 17184 4224 17190 4276
rect 17494 4224 17500 4276
rect 17552 4264 17558 4276
rect 21358 4264 21364 4276
rect 17552 4236 21364 4264
rect 17552 4224 17558 4236
rect 21358 4224 21364 4236
rect 21416 4224 21422 4276
rect 9858 4156 9864 4208
rect 9916 4196 9922 4208
rect 14274 4196 14280 4208
rect 9916 4168 14280 4196
rect 9916 4156 9922 4168
rect 14274 4156 14280 4168
rect 14332 4156 14338 4208
rect 14550 4156 14556 4208
rect 14608 4196 14614 4208
rect 14608 4168 14688 4196
rect 14608 4156 14614 4168
rect 12342 4128 12348 4140
rect 6963 4100 7880 4128
rect 7944 4100 12348 4128
rect 6963 4097 6975 4100
rect 6917 4091 6975 4097
rect 1771 4063 1829 4069
rect 1771 4029 1783 4063
rect 1817 4029 1829 4063
rect 1771 4023 1829 4029
rect 1780 3992 1808 4023
rect 2774 4020 2780 4072
rect 2832 4060 2838 4072
rect 2869 4063 2927 4069
rect 2869 4060 2881 4063
rect 2832 4032 2881 4060
rect 2832 4020 2838 4032
rect 2869 4029 2881 4032
rect 2915 4029 2927 4063
rect 2869 4023 2927 4029
rect 3878 4020 3884 4072
rect 3936 4060 3942 4072
rect 7944 4069 7972 4100
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 12986 4128 12992 4140
rect 12947 4100 12992 4128
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 13173 4131 13231 4137
rect 13173 4097 13185 4131
rect 13219 4128 13231 4131
rect 13722 4128 13728 4140
rect 13219 4100 13728 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 14660 4137 14688 4168
rect 16298 4156 16304 4208
rect 16356 4156 16362 4208
rect 17034 4156 17040 4208
rect 17092 4196 17098 4208
rect 17092 4168 18644 4196
rect 17092 4156 17098 4168
rect 14645 4131 14703 4137
rect 14645 4097 14657 4131
rect 14691 4097 14703 4131
rect 16316 4128 16344 4156
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16316 4100 16681 4128
rect 14645 4091 14703 4097
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 17402 4088 17408 4140
rect 17460 4128 17466 4140
rect 18616 4137 18644 4168
rect 18509 4131 18567 4137
rect 18509 4128 18521 4131
rect 17460 4100 18521 4128
rect 17460 4088 17466 4100
rect 18509 4097 18521 4100
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4097 18659 4131
rect 18601 4091 18659 4097
rect 18782 4088 18788 4140
rect 18840 4128 18846 4140
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 18840 4100 20085 4128
rect 18840 4088 18846 4100
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20254 4128 20260 4140
rect 20215 4100 20260 4128
rect 20073 4091 20131 4097
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 3973 4063 4031 4069
rect 3973 4060 3985 4063
rect 3936 4032 3985 4060
rect 3936 4020 3942 4032
rect 3973 4029 3985 4032
rect 4019 4029 4031 4063
rect 3973 4023 4031 4029
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4029 7987 4063
rect 9030 4060 9036 4072
rect 8991 4032 9036 4060
rect 7929 4023 7987 4029
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4060 10195 4063
rect 10778 4060 10784 4072
rect 10183 4032 10784 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 11229 4063 11287 4069
rect 11229 4029 11241 4063
rect 11275 4060 11287 4063
rect 12250 4060 12256 4072
rect 11275 4032 12256 4060
rect 11275 4029 11287 4032
rect 11229 4023 11287 4029
rect 12250 4020 12256 4032
rect 12308 4020 12314 4072
rect 14461 4063 14519 4069
rect 14461 4029 14473 4063
rect 14507 4060 14519 4063
rect 14734 4060 14740 4072
rect 14507 4032 14740 4060
rect 14507 4029 14519 4032
rect 14461 4023 14519 4029
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 16114 4020 16120 4072
rect 16172 4020 16178 4072
rect 16298 4020 16304 4072
rect 16356 4060 16362 4072
rect 17589 4063 17647 4069
rect 17589 4060 17601 4063
rect 16356 4032 17601 4060
rect 16356 4020 16362 4032
rect 17589 4029 17601 4032
rect 17635 4060 17647 4063
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 17635 4032 18429 4060
rect 17635 4029 17647 4032
rect 17589 4023 17647 4029
rect 18417 4029 18429 4032
rect 18463 4060 18475 4063
rect 18877 4063 18935 4069
rect 18877 4060 18889 4063
rect 18463 4032 18889 4060
rect 18463 4029 18475 4032
rect 18417 4023 18475 4029
rect 18877 4029 18889 4032
rect 18923 4029 18935 4063
rect 18877 4023 18935 4029
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 20438 4060 20444 4072
rect 19392 4032 20444 4060
rect 19392 4020 19398 4032
rect 20438 4020 20444 4032
rect 20496 4020 20502 4072
rect 10042 3992 10048 4004
rect 1780 3964 10048 3992
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 10502 3992 10508 4004
rect 10152 3964 10508 3992
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 1949 3927 2007 3933
rect 1949 3924 1961 3927
rect 1452 3896 1961 3924
rect 1452 3884 1458 3896
rect 1949 3893 1961 3896
rect 1995 3893 2007 3927
rect 3050 3924 3056 3936
rect 3011 3896 3056 3924
rect 1949 3887 2007 3893
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 4154 3924 4160 3936
rect 4115 3896 4160 3924
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8202 3924 8208 3936
rect 8159 3896 8208 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9217 3927 9275 3933
rect 9217 3924 9229 3927
rect 8996 3896 9229 3924
rect 8996 3884 9002 3896
rect 9217 3893 9229 3896
rect 9263 3893 9275 3927
rect 9217 3887 9275 3893
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 10152 3924 10180 3964
rect 10502 3952 10508 3964
rect 10560 3952 10566 4004
rect 16132 3992 16160 4020
rect 11440 3964 16160 3992
rect 16485 3995 16543 4001
rect 11440 3933 11468 3964
rect 16485 3961 16497 3995
rect 16531 3992 16543 3995
rect 17494 3992 17500 4004
rect 16531 3964 17500 3992
rect 16531 3961 16543 3964
rect 16485 3955 16543 3961
rect 17494 3952 17500 3964
rect 17552 3952 17558 4004
rect 17862 3952 17868 4004
rect 17920 3992 17926 4004
rect 19981 3995 20039 4001
rect 19981 3992 19993 3995
rect 17920 3964 19993 3992
rect 17920 3952 17926 3964
rect 19981 3961 19993 3964
rect 20027 3961 20039 3995
rect 19981 3955 20039 3961
rect 9732 3896 10180 3924
rect 11425 3927 11483 3933
rect 9732 3884 9738 3896
rect 11425 3893 11437 3927
rect 11471 3893 11483 3927
rect 11425 3887 11483 3893
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12529 3927 12587 3933
rect 12529 3924 12541 3927
rect 12492 3896 12541 3924
rect 12492 3884 12498 3896
rect 12529 3893 12541 3896
rect 12575 3893 12587 3927
rect 12894 3924 12900 3936
rect 12855 3896 12900 3924
rect 12529 3887 12587 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 13906 3884 13912 3936
rect 13964 3924 13970 3936
rect 14093 3927 14151 3933
rect 14093 3924 14105 3927
rect 13964 3896 14105 3924
rect 13964 3884 13970 3896
rect 14093 3893 14105 3896
rect 14139 3893 14151 3927
rect 14093 3887 14151 3893
rect 14553 3927 14611 3933
rect 14553 3893 14565 3927
rect 14599 3924 14611 3927
rect 15562 3924 15568 3936
rect 14599 3896 15568 3924
rect 14599 3893 14611 3896
rect 14553 3887 14611 3893
rect 15562 3884 15568 3896
rect 15620 3884 15626 3936
rect 16022 3884 16028 3936
rect 16080 3924 16086 3936
rect 16117 3927 16175 3933
rect 16117 3924 16129 3927
rect 16080 3896 16129 3924
rect 16080 3884 16086 3896
rect 16117 3893 16129 3896
rect 16163 3893 16175 3927
rect 16117 3887 16175 3893
rect 16390 3884 16396 3936
rect 16448 3924 16454 3936
rect 16577 3927 16635 3933
rect 16577 3924 16589 3927
rect 16448 3896 16589 3924
rect 16448 3884 16454 3896
rect 16577 3893 16589 3896
rect 16623 3893 16635 3927
rect 16577 3887 16635 3893
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 16816 3896 18061 3924
rect 16816 3884 16822 3896
rect 18049 3893 18061 3896
rect 18095 3893 18107 3927
rect 18049 3887 18107 3893
rect 19058 3884 19064 3936
rect 19116 3924 19122 3936
rect 19613 3927 19671 3933
rect 19613 3924 19625 3927
rect 19116 3896 19625 3924
rect 19116 3884 19122 3896
rect 19613 3893 19625 3896
rect 19659 3893 19671 3927
rect 19613 3887 19671 3893
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 2041 3723 2099 3729
rect 2041 3689 2053 3723
rect 2087 3720 2099 3723
rect 2130 3720 2136 3732
rect 2087 3692 2136 3720
rect 2087 3689 2099 3692
rect 2041 3683 2099 3689
rect 2130 3680 2136 3692
rect 2188 3680 2194 3732
rect 2961 3723 3019 3729
rect 2961 3689 2973 3723
rect 3007 3720 3019 3723
rect 4890 3720 4896 3732
rect 3007 3692 4896 3720
rect 3007 3689 3019 3692
rect 2961 3683 3019 3689
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 5902 3680 5908 3732
rect 5960 3720 5966 3732
rect 9674 3720 9680 3732
rect 5960 3692 9680 3720
rect 5960 3680 5966 3692
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 10042 3720 10048 3732
rect 10003 3692 10048 3720
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 11149 3723 11207 3729
rect 11149 3689 11161 3723
rect 11195 3720 11207 3723
rect 11974 3720 11980 3732
rect 11195 3692 11980 3720
rect 11195 3689 11207 3692
rect 11149 3683 11207 3689
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 12069 3723 12127 3729
rect 12069 3689 12081 3723
rect 12115 3720 12127 3723
rect 12158 3720 12164 3732
rect 12115 3692 12164 3720
rect 12115 3689 12127 3692
rect 12069 3683 12127 3689
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 12492 3692 12537 3720
rect 12492 3680 12498 3692
rect 12894 3680 12900 3732
rect 12952 3720 12958 3732
rect 13633 3723 13691 3729
rect 13633 3720 13645 3723
rect 12952 3692 13645 3720
rect 12952 3680 12958 3692
rect 13633 3689 13645 3692
rect 13679 3689 13691 3723
rect 13998 3720 14004 3732
rect 13959 3692 14004 3720
rect 13633 3683 13691 3689
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 16393 3723 16451 3729
rect 16393 3689 16405 3723
rect 16439 3720 16451 3723
rect 16758 3720 16764 3732
rect 16439 3692 16764 3720
rect 16439 3689 16451 3692
rect 16393 3683 16451 3689
rect 16758 3680 16764 3692
rect 16816 3680 16822 3732
rect 16850 3680 16856 3732
rect 16908 3720 16914 3732
rect 17770 3720 17776 3732
rect 16908 3692 17776 3720
rect 16908 3680 16914 3692
rect 17770 3680 17776 3692
rect 17828 3680 17834 3732
rect 18049 3723 18107 3729
rect 18049 3689 18061 3723
rect 18095 3720 18107 3723
rect 18138 3720 18144 3732
rect 18095 3692 18144 3720
rect 18095 3689 18107 3692
rect 18049 3683 18107 3689
rect 18138 3680 18144 3692
rect 18196 3680 18202 3732
rect 19610 3720 19616 3732
rect 19571 3692 19616 3720
rect 19610 3680 19616 3692
rect 19668 3680 19674 3732
rect 8573 3655 8631 3661
rect 8573 3621 8585 3655
rect 8619 3652 8631 3655
rect 8662 3652 8668 3664
rect 8619 3624 8668 3652
rect 8619 3621 8631 3624
rect 8573 3615 8631 3621
rect 8662 3612 8668 3624
rect 8720 3612 8726 3664
rect 10870 3652 10876 3664
rect 9692 3624 10876 3652
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 2222 3584 2228 3596
rect 1903 3556 2228 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 4062 3584 4068 3596
rect 4023 3556 4068 3584
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 6595 3556 9597 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 9585 3553 9597 3556
rect 9631 3553 9643 3587
rect 9585 3547 9643 3553
rect 7561 3519 7619 3525
rect 7561 3485 7573 3519
rect 7607 3516 7619 3519
rect 9692 3516 9720 3624
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 12529 3655 12587 3661
rect 12529 3621 12541 3655
rect 12575 3652 12587 3655
rect 12618 3652 12624 3664
rect 12575 3624 12624 3652
rect 12575 3621 12587 3624
rect 12529 3615 12587 3621
rect 12618 3612 12624 3624
rect 12676 3612 12682 3664
rect 13814 3612 13820 3664
rect 13872 3652 13878 3664
rect 14093 3655 14151 3661
rect 14093 3652 14105 3655
rect 13872 3624 14105 3652
rect 13872 3612 13878 3624
rect 14093 3621 14105 3624
rect 14139 3652 14151 3655
rect 14366 3652 14372 3664
rect 14139 3624 14372 3652
rect 14139 3621 14151 3624
rect 14093 3615 14151 3621
rect 14366 3612 14372 3624
rect 14424 3612 14430 3664
rect 16114 3612 16120 3664
rect 16172 3652 16178 3664
rect 16172 3624 16252 3652
rect 16172 3612 16178 3624
rect 9858 3544 9864 3596
rect 9916 3584 9922 3596
rect 9916 3556 9961 3584
rect 9916 3544 9922 3556
rect 10686 3544 10692 3596
rect 10744 3584 10750 3596
rect 10965 3587 11023 3593
rect 10965 3584 10977 3587
rect 10744 3556 10977 3584
rect 10744 3544 10750 3556
rect 10965 3553 10977 3556
rect 11011 3553 11023 3587
rect 10965 3547 11023 3553
rect 13722 3544 13728 3596
rect 13780 3584 13786 3596
rect 14642 3584 14648 3596
rect 13780 3556 14648 3584
rect 13780 3544 13786 3556
rect 14642 3544 14648 3556
rect 14700 3544 14706 3596
rect 16224 3584 16252 3624
rect 17310 3612 17316 3664
rect 17368 3652 17374 3664
rect 17368 3624 18184 3652
rect 17368 3612 17374 3624
rect 17957 3587 18015 3593
rect 16224 3556 16620 3584
rect 7607 3488 9720 3516
rect 9769 3519 9827 3525
rect 7607 3485 7619 3488
rect 7561 3479 7619 3485
rect 9769 3485 9781 3519
rect 9815 3516 9827 3519
rect 10594 3516 10600 3528
rect 9815 3488 10600 3516
rect 9815 3485 9827 3488
rect 9769 3479 9827 3485
rect 10594 3476 10600 3488
rect 10652 3476 10658 3528
rect 12713 3519 12771 3525
rect 12713 3485 12725 3519
rect 12759 3516 12771 3519
rect 12802 3516 12808 3528
rect 12759 3488 12808 3516
rect 12759 3485 12771 3488
rect 12713 3479 12771 3485
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 14182 3476 14188 3528
rect 14240 3516 14246 3528
rect 16482 3516 16488 3528
rect 14240 3488 14285 3516
rect 16443 3488 16488 3516
rect 14240 3476 14246 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 16592 3525 16620 3556
rect 17957 3553 17969 3587
rect 18003 3584 18015 3587
rect 18046 3584 18052 3596
rect 18003 3556 18052 3584
rect 18003 3553 18015 3556
rect 17957 3547 18015 3553
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 18156 3525 18184 3624
rect 19150 3612 19156 3664
rect 19208 3652 19214 3664
rect 19521 3655 19579 3661
rect 19521 3652 19533 3655
rect 19208 3624 19533 3652
rect 19208 3612 19214 3624
rect 19521 3621 19533 3624
rect 19567 3621 19579 3655
rect 19521 3615 19579 3621
rect 18322 3544 18328 3596
rect 18380 3584 18386 3596
rect 19978 3584 19984 3596
rect 18380 3556 19984 3584
rect 18380 3544 18386 3556
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 16577 3519 16635 3525
rect 16577 3485 16589 3519
rect 16623 3485 16635 3519
rect 16577 3479 16635 3485
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 18874 3476 18880 3528
rect 18932 3516 18938 3528
rect 19334 3516 19340 3528
rect 18932 3488 19340 3516
rect 18932 3476 18938 3488
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 19797 3519 19855 3525
rect 19797 3485 19809 3519
rect 19843 3516 19855 3519
rect 20254 3516 20260 3528
rect 19843 3488 20260 3516
rect 19843 3485 19855 3488
rect 19797 3479 19855 3485
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 4246 3448 4252 3460
rect 4207 3420 4252 3448
rect 4246 3408 4252 3420
rect 4304 3408 4310 3460
rect 5626 3448 5632 3460
rect 4356 3420 5632 3448
rect 3970 3340 3976 3392
rect 4028 3380 4034 3392
rect 4356 3380 4384 3420
rect 5626 3408 5632 3420
rect 5684 3408 5690 3460
rect 5810 3408 5816 3460
rect 5868 3448 5874 3460
rect 16025 3451 16083 3457
rect 16025 3448 16037 3451
rect 5868 3420 16037 3448
rect 5868 3408 5874 3420
rect 16025 3417 16037 3420
rect 16071 3417 16083 3451
rect 16025 3411 16083 3417
rect 17494 3408 17500 3460
rect 17552 3448 17558 3460
rect 17589 3451 17647 3457
rect 17589 3448 17601 3451
rect 17552 3420 17601 3448
rect 17552 3408 17558 3420
rect 17589 3417 17601 3420
rect 17635 3417 17647 3451
rect 20714 3448 20720 3460
rect 17589 3411 17647 3417
rect 17696 3420 20720 3448
rect 4028 3352 4384 3380
rect 4028 3340 4034 3352
rect 4798 3340 4804 3392
rect 4856 3380 4862 3392
rect 11974 3380 11980 3392
rect 4856 3352 11980 3380
rect 4856 3340 4862 3352
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 12434 3340 12440 3392
rect 12492 3380 12498 3392
rect 17696 3380 17724 3420
rect 20714 3408 20720 3420
rect 20772 3408 20778 3460
rect 19150 3380 19156 3392
rect 12492 3352 17724 3380
rect 19111 3352 19156 3380
rect 12492 3340 12498 3352
rect 19150 3340 19156 3352
rect 19208 3340 19214 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 1302 3136 1308 3188
rect 1360 3176 1366 3188
rect 1949 3179 2007 3185
rect 1949 3176 1961 3179
rect 1360 3148 1961 3176
rect 1360 3136 1366 3148
rect 1949 3145 1961 3148
rect 1995 3145 2007 3179
rect 1949 3139 2007 3145
rect 2498 3136 2504 3188
rect 2556 3176 2562 3188
rect 5810 3176 5816 3188
rect 2556 3148 5816 3176
rect 2556 3136 2562 3148
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 5905 3179 5963 3185
rect 5905 3145 5917 3179
rect 5951 3176 5963 3179
rect 10321 3179 10379 3185
rect 5951 3148 9168 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 8570 3108 8576 3120
rect 8531 3080 8576 3108
rect 8570 3068 8576 3080
rect 8628 3068 8634 3120
rect 9140 3108 9168 3148
rect 10321 3145 10333 3179
rect 10367 3176 10379 3179
rect 10962 3176 10968 3188
rect 10367 3148 10968 3176
rect 10367 3145 10379 3148
rect 10321 3139 10379 3145
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 11425 3179 11483 3185
rect 11425 3145 11437 3179
rect 11471 3176 11483 3179
rect 11790 3176 11796 3188
rect 11471 3148 11796 3176
rect 11471 3145 11483 3148
rect 11425 3139 11483 3145
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 16298 3176 16304 3188
rect 12032 3148 16304 3176
rect 12032 3136 12038 3148
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 16393 3179 16451 3185
rect 16393 3145 16405 3179
rect 16439 3176 16451 3179
rect 16482 3176 16488 3188
rect 16439 3148 16488 3176
rect 16439 3145 16451 3148
rect 16393 3139 16451 3145
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 16666 3136 16672 3188
rect 16724 3176 16730 3188
rect 20162 3176 20168 3188
rect 16724 3148 20168 3176
rect 16724 3136 16730 3148
rect 20162 3136 20168 3148
rect 20220 3136 20226 3188
rect 12434 3108 12440 3120
rect 9140 3080 12440 3108
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 12618 3068 12624 3120
rect 12676 3108 12682 3120
rect 18049 3111 18107 3117
rect 18049 3108 18061 3111
rect 12676 3080 18061 3108
rect 12676 3068 12682 3080
rect 18049 3077 18061 3080
rect 18095 3077 18107 3111
rect 18049 3071 18107 3077
rect 9306 3000 9312 3052
rect 9364 3040 9370 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 9364 3012 13001 3040
rect 9364 3000 9370 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 14550 3040 14556 3052
rect 14511 3012 14556 3040
rect 12989 3003 13047 3009
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 14642 3000 14648 3052
rect 14700 3040 14706 3052
rect 17034 3040 17040 3052
rect 14700 3012 14745 3040
rect 16995 3012 17040 3040
rect 14700 3000 14706 3012
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 18598 3040 18604 3052
rect 18559 3012 18604 3040
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 1762 2972 1768 2984
rect 1723 2944 1768 2972
rect 1762 2932 1768 2944
rect 1820 2932 1826 2984
rect 2866 2972 2872 2984
rect 2827 2944 2872 2972
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 8754 2972 8760 2984
rect 7239 2944 8760 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 8754 2932 8760 2944
rect 8812 2932 8818 2984
rect 10134 2972 10140 2984
rect 10095 2944 10140 2972
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 11238 2972 11244 2984
rect 11199 2944 11244 2972
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 12710 2932 12716 2984
rect 12768 2972 12774 2984
rect 12805 2975 12863 2981
rect 12805 2972 12817 2975
rect 12768 2944 12817 2972
rect 12768 2932 12774 2944
rect 12805 2941 12817 2944
rect 12851 2941 12863 2975
rect 12805 2935 12863 2941
rect 14274 2932 14280 2984
rect 14332 2972 14338 2984
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 14332 2944 14473 2972
rect 14332 2932 14338 2944
rect 14461 2941 14473 2944
rect 14507 2941 14519 2975
rect 14568 2972 14596 3000
rect 15470 2972 15476 2984
rect 14568 2944 15476 2972
rect 14461 2935 14519 2941
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 16758 2972 16764 2984
rect 16719 2944 16764 2972
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 18509 2975 18567 2981
rect 18509 2941 18521 2975
rect 18555 2972 18567 2975
rect 19150 2972 19156 2984
rect 18555 2944 19156 2972
rect 18555 2941 18567 2944
rect 18509 2935 18567 2941
rect 19150 2932 19156 2944
rect 19208 2932 19214 2984
rect 19613 2975 19671 2981
rect 19613 2941 19625 2975
rect 19659 2972 19671 2975
rect 19702 2972 19708 2984
rect 19659 2944 19708 2972
rect 19659 2941 19671 2944
rect 19613 2935 19671 2941
rect 19702 2932 19708 2944
rect 19760 2932 19766 2984
rect 7098 2864 7104 2916
rect 7156 2904 7162 2916
rect 7438 2907 7496 2913
rect 7438 2904 7450 2907
rect 7156 2876 7450 2904
rect 7156 2864 7162 2876
rect 7438 2873 7450 2876
rect 7484 2873 7496 2907
rect 7438 2867 7496 2873
rect 7558 2864 7564 2916
rect 7616 2904 7622 2916
rect 10502 2904 10508 2916
rect 7616 2876 10508 2904
rect 7616 2864 7622 2876
rect 10502 2864 10508 2876
rect 10560 2864 10566 2916
rect 10594 2864 10600 2916
rect 10652 2904 10658 2916
rect 14182 2904 14188 2916
rect 10652 2876 14188 2904
rect 10652 2864 10658 2876
rect 14182 2864 14188 2876
rect 14240 2864 14246 2916
rect 16853 2907 16911 2913
rect 16853 2873 16865 2907
rect 16899 2904 16911 2907
rect 16942 2904 16948 2916
rect 16899 2876 16948 2904
rect 16899 2873 16911 2876
rect 16853 2867 16911 2873
rect 16942 2864 16948 2876
rect 17000 2864 17006 2916
rect 18417 2907 18475 2913
rect 18417 2873 18429 2907
rect 18463 2904 18475 2907
rect 19058 2904 19064 2916
rect 18463 2876 19064 2904
rect 18463 2873 18475 2876
rect 18417 2867 18475 2873
rect 19058 2864 19064 2876
rect 19116 2864 19122 2916
rect 3050 2836 3056 2848
rect 3011 2808 3056 2836
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 7282 2796 7288 2848
rect 7340 2836 7346 2848
rect 11238 2836 11244 2848
rect 7340 2808 11244 2836
rect 7340 2796 7346 2808
rect 11238 2796 11244 2808
rect 11296 2796 11302 2848
rect 14093 2839 14151 2845
rect 14093 2805 14105 2839
rect 14139 2836 14151 2839
rect 16574 2836 16580 2848
rect 14139 2808 16580 2836
rect 14139 2805 14151 2808
rect 14093 2799 14151 2805
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 19242 2796 19248 2848
rect 19300 2836 19306 2848
rect 19797 2839 19855 2845
rect 19797 2836 19809 2839
rect 19300 2808 19809 2836
rect 19300 2796 19306 2808
rect 19797 2805 19809 2808
rect 19843 2805 19855 2839
rect 19797 2799 19855 2805
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 4062 2592 4068 2644
rect 4120 2632 4126 2644
rect 5350 2632 5356 2644
rect 4120 2604 5356 2632
rect 4120 2592 4126 2604
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 9122 2632 9128 2644
rect 8711 2604 9128 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 10413 2635 10471 2641
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 11054 2632 11060 2644
rect 10459 2604 11060 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 11609 2635 11667 2641
rect 11609 2601 11621 2635
rect 11655 2632 11667 2635
rect 13262 2632 13268 2644
rect 11655 2604 13268 2632
rect 11655 2601 11667 2604
rect 11609 2595 11667 2601
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 13814 2632 13820 2644
rect 13775 2604 13820 2632
rect 13814 2592 13820 2604
rect 13872 2592 13878 2644
rect 14182 2632 14188 2644
rect 14143 2604 14188 2632
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 16390 2592 16396 2644
rect 16448 2632 16454 2644
rect 16485 2635 16543 2641
rect 16485 2632 16497 2635
rect 16448 2604 16497 2632
rect 16448 2592 16454 2604
rect 16485 2601 16497 2604
rect 16531 2601 16543 2635
rect 16485 2595 16543 2601
rect 16945 2635 17003 2641
rect 16945 2601 16957 2635
rect 16991 2632 17003 2635
rect 17126 2632 17132 2644
rect 16991 2604 17132 2632
rect 16991 2601 17003 2604
rect 16945 2595 17003 2601
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 19613 2635 19671 2641
rect 19613 2601 19625 2635
rect 19659 2632 19671 2635
rect 19794 2632 19800 2644
rect 19659 2604 19800 2632
rect 19659 2601 19671 2604
rect 19613 2595 19671 2601
rect 19794 2592 19800 2604
rect 19852 2592 19858 2644
rect 13538 2524 13544 2576
rect 13596 2564 13602 2576
rect 15473 2567 15531 2573
rect 13596 2536 15240 2564
rect 13596 2524 13602 2536
rect 1854 2496 1860 2508
rect 1815 2468 1860 2496
rect 1854 2456 1860 2468
rect 1912 2456 1918 2508
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2465 11483 2499
rect 11425 2459 11483 2465
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 12713 2499 12771 2505
rect 12713 2496 12725 2499
rect 12667 2468 12725 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 12713 2465 12725 2468
rect 12759 2465 12771 2499
rect 15212 2496 15240 2536
rect 15473 2533 15485 2567
rect 15519 2564 15531 2567
rect 17862 2564 17868 2576
rect 15519 2536 17868 2564
rect 15519 2533 15531 2536
rect 15473 2527 15531 2533
rect 17862 2524 17868 2536
rect 17920 2524 17926 2576
rect 16853 2499 16911 2505
rect 16853 2496 16865 2499
rect 15212 2468 16865 2496
rect 12713 2459 12771 2465
rect 16853 2465 16865 2468
rect 16899 2465 16911 2499
rect 16853 2459 16911 2465
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 5442 2428 5448 2440
rect 2832 2400 5448 2428
rect 2832 2388 2838 2400
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 11440 2428 11468 2459
rect 18046 2456 18052 2508
rect 18104 2496 18110 2508
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18104 2468 18337 2496
rect 18104 2456 18110 2468
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 19426 2496 19432 2508
rect 19387 2468 19432 2496
rect 18325 2459 18383 2465
rect 19426 2456 19432 2468
rect 19484 2456 19490 2508
rect 11440 2400 14228 2428
rect 7837 2363 7895 2369
rect 7837 2329 7849 2363
rect 7883 2360 7895 2363
rect 13722 2360 13728 2372
rect 7883 2332 13728 2360
rect 7883 2329 7895 2332
rect 7837 2323 7895 2329
rect 13722 2320 13728 2332
rect 13780 2320 13786 2372
rect 2038 2292 2044 2304
rect 1999 2264 2044 2292
rect 2038 2252 2044 2264
rect 2096 2252 2102 2304
rect 6914 2252 6920 2304
rect 6972 2292 6978 2304
rect 12621 2295 12679 2301
rect 12621 2292 12633 2295
rect 6972 2264 12633 2292
rect 6972 2252 6978 2264
rect 12621 2261 12633 2264
rect 12667 2261 12679 2295
rect 12621 2255 12679 2261
rect 12897 2295 12955 2301
rect 12897 2261 12909 2295
rect 12943 2292 12955 2295
rect 13446 2292 13452 2304
rect 12943 2264 13452 2292
rect 12943 2261 12955 2264
rect 12897 2255 12955 2261
rect 13446 2252 13452 2264
rect 13504 2252 13510 2304
rect 14200 2292 14228 2400
rect 14274 2388 14280 2440
rect 14332 2428 14338 2440
rect 14461 2431 14519 2437
rect 14332 2400 14377 2428
rect 14332 2388 14338 2400
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 14642 2428 14648 2440
rect 14507 2400 14648 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 14642 2388 14648 2400
rect 14700 2388 14706 2440
rect 17129 2431 17187 2437
rect 17129 2397 17141 2431
rect 17175 2428 17187 2431
rect 17310 2428 17316 2440
rect 17175 2400 17316 2428
rect 17175 2397 17187 2400
rect 17129 2391 17187 2397
rect 17310 2388 17316 2400
rect 17368 2388 17374 2440
rect 16206 2320 16212 2372
rect 16264 2360 16270 2372
rect 18509 2363 18567 2369
rect 18509 2360 18521 2363
rect 16264 2332 18521 2360
rect 16264 2320 16270 2332
rect 18509 2329 18521 2332
rect 18555 2329 18567 2363
rect 18509 2323 18567 2329
rect 18690 2292 18696 2304
rect 14200 2264 18696 2292
rect 18690 2252 18696 2264
rect 18748 2252 18754 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 2038 2048 2044 2100
rect 2096 2088 2102 2100
rect 13725 2091 13783 2097
rect 13725 2088 13737 2091
rect 2096 2060 13737 2088
rect 2096 2048 2102 2060
rect 13725 2057 13737 2060
rect 13771 2057 13783 2091
rect 13725 2051 13783 2057
rect 7466 1980 7472 2032
rect 7524 2020 7530 2032
rect 14274 2020 14280 2032
rect 7524 1992 14280 2020
rect 7524 1980 7530 1992
rect 14274 1980 14280 1992
rect 14332 1980 14338 2032
rect 14366 1980 14372 2032
rect 14424 2020 14430 2032
rect 18506 2020 18512 2032
rect 14424 1992 18512 2020
rect 14424 1980 14430 1992
rect 18506 1980 18512 1992
rect 18564 1980 18570 2032
rect 13998 1844 14004 1896
rect 14056 1884 14062 1896
rect 18690 1884 18696 1896
rect 14056 1856 18696 1884
rect 14056 1844 14062 1856
rect 18690 1844 18696 1856
rect 18748 1844 18754 1896
rect 13722 1776 13728 1828
rect 13780 1816 13786 1828
rect 19518 1816 19524 1828
rect 13780 1788 19524 1816
rect 13780 1776 13786 1788
rect 19518 1776 19524 1788
rect 19576 1776 19582 1828
rect 8846 1708 8852 1760
rect 8904 1748 8910 1760
rect 18046 1748 18052 1760
rect 8904 1720 18052 1748
rect 8904 1708 8910 1720
rect 18046 1708 18052 1720
rect 18104 1708 18110 1760
rect 13725 1683 13783 1689
rect 13725 1649 13737 1683
rect 13771 1680 13783 1683
rect 21450 1680 21456 1692
rect 13771 1652 21456 1680
rect 13771 1649 13783 1652
rect 13725 1643 13783 1649
rect 21450 1640 21456 1652
rect 21508 1640 21514 1692
rect 10502 1572 10508 1624
rect 10560 1612 10566 1624
rect 16114 1612 16120 1624
rect 10560 1584 16120 1612
rect 10560 1572 10566 1584
rect 16114 1572 16120 1584
rect 16172 1572 16178 1624
rect 13078 1300 13084 1352
rect 13136 1340 13142 1352
rect 18138 1340 18144 1352
rect 13136 1312 18144 1340
rect 13136 1300 13142 1312
rect 18138 1300 18144 1312
rect 18196 1300 18202 1352
rect 2314 1232 2320 1284
rect 2372 1272 2378 1284
rect 5902 1272 5908 1284
rect 2372 1244 5908 1272
rect 2372 1232 2378 1244
rect 5902 1232 5908 1244
rect 5960 1232 5966 1284
<< via1 >>
rect 3516 21632 3568 21684
rect 5172 21632 5224 21684
rect 15200 21156 15252 21208
rect 17960 21156 18012 21208
rect 17960 20952 18012 21004
rect 18236 20952 18288 21004
rect 4804 20884 4856 20936
rect 5356 20884 5408 20936
rect 3700 20816 3752 20868
rect 6276 20816 6328 20868
rect 3516 20748 3568 20800
rect 4896 20748 4948 20800
rect 8668 20748 8720 20800
rect 18052 20748 18104 20800
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 5264 20544 5316 20596
rect 8760 20544 8812 20596
rect 9312 20544 9364 20596
rect 13912 20544 13964 20596
rect 15200 20544 15252 20596
rect 17868 20544 17920 20596
rect 2688 20408 2740 20460
rect 3056 20408 3108 20460
rect 6828 20340 6880 20392
rect 18696 20476 18748 20528
rect 7288 20408 7340 20460
rect 11060 20408 11112 20460
rect 13268 20451 13320 20460
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 13360 20408 13412 20460
rect 17132 20451 17184 20460
rect 9036 20340 9088 20392
rect 3976 20272 4028 20324
rect 4988 20272 5040 20324
rect 12164 20340 12216 20392
rect 14372 20340 14424 20392
rect 15200 20340 15252 20392
rect 17132 20417 17141 20451
rect 17141 20417 17175 20451
rect 17175 20417 17184 20451
rect 17132 20408 17184 20417
rect 17316 20451 17368 20460
rect 17316 20417 17325 20451
rect 17325 20417 17359 20451
rect 17359 20417 17368 20451
rect 17316 20408 17368 20417
rect 19892 20408 19944 20460
rect 10416 20272 10468 20324
rect 17040 20315 17092 20324
rect 17040 20281 17049 20315
rect 17049 20281 17083 20315
rect 17083 20281 17092 20315
rect 17040 20272 17092 20281
rect 2228 20204 2280 20256
rect 2780 20247 2832 20256
rect 2780 20213 2789 20247
rect 2789 20213 2823 20247
rect 2823 20213 2832 20247
rect 2780 20204 2832 20213
rect 3884 20204 3936 20256
rect 4712 20204 4764 20256
rect 5264 20204 5316 20256
rect 7656 20204 7708 20256
rect 8208 20204 8260 20256
rect 8484 20247 8536 20256
rect 8484 20213 8493 20247
rect 8493 20213 8527 20247
rect 8527 20213 8536 20247
rect 8484 20204 8536 20213
rect 8760 20204 8812 20256
rect 10692 20247 10744 20256
rect 10692 20213 10701 20247
rect 10701 20213 10735 20247
rect 10735 20213 10744 20247
rect 10692 20204 10744 20213
rect 10968 20204 11020 20256
rect 12348 20204 12400 20256
rect 13176 20204 13228 20256
rect 16672 20247 16724 20256
rect 16672 20213 16681 20247
rect 16681 20213 16715 20247
rect 16715 20213 16724 20247
rect 16672 20204 16724 20213
rect 18972 20247 19024 20256
rect 18972 20213 18981 20247
rect 18981 20213 19015 20247
rect 19015 20213 19024 20247
rect 18972 20204 19024 20213
rect 19064 20204 19116 20256
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 4160 20000 4212 20052
rect 4712 20043 4764 20052
rect 4712 20009 4721 20043
rect 4721 20009 4755 20043
rect 4755 20009 4764 20043
rect 4712 20000 4764 20009
rect 5448 20000 5500 20052
rect 10416 20000 10468 20052
rect 16672 20000 16724 20052
rect 8944 19932 8996 19984
rect 9036 19932 9088 19984
rect 5724 19864 5776 19916
rect 1860 19796 1912 19848
rect 3056 19839 3108 19848
rect 3056 19805 3065 19839
rect 3065 19805 3099 19839
rect 3099 19805 3108 19839
rect 3056 19796 3108 19805
rect 4896 19839 4948 19848
rect 4896 19805 4905 19839
rect 4905 19805 4939 19839
rect 4939 19805 4948 19839
rect 6368 19839 6420 19848
rect 4896 19796 4948 19805
rect 6368 19805 6377 19839
rect 6377 19805 6411 19839
rect 6411 19805 6420 19839
rect 6368 19796 6420 19805
rect 6828 19864 6880 19916
rect 7288 19796 7340 19848
rect 2872 19660 2924 19712
rect 5448 19660 5500 19712
rect 7288 19660 7340 19712
rect 12440 19932 12492 19984
rect 13912 19932 13964 19984
rect 9496 19796 9548 19848
rect 11060 19796 11112 19848
rect 14372 19864 14424 19916
rect 15292 19907 15344 19916
rect 15292 19873 15301 19907
rect 15301 19873 15335 19907
rect 15335 19873 15344 19907
rect 15292 19864 15344 19873
rect 17132 19839 17184 19848
rect 13268 19728 13320 19780
rect 17132 19805 17141 19839
rect 17141 19805 17175 19839
rect 17175 19805 17184 19839
rect 17132 19796 17184 19805
rect 17316 19839 17368 19848
rect 17316 19805 17325 19839
rect 17325 19805 17359 19839
rect 17359 19805 17368 19839
rect 17316 19796 17368 19805
rect 19892 19839 19944 19848
rect 14096 19728 14148 19780
rect 19892 19805 19901 19839
rect 19901 19805 19935 19839
rect 19935 19805 19944 19839
rect 19892 19796 19944 19805
rect 10876 19660 10928 19712
rect 11060 19703 11112 19712
rect 11060 19669 11069 19703
rect 11069 19669 11103 19703
rect 11103 19669 11112 19703
rect 11060 19660 11112 19669
rect 11888 19703 11940 19712
rect 11888 19669 11897 19703
rect 11897 19669 11931 19703
rect 11931 19669 11940 19703
rect 11888 19660 11940 19669
rect 18052 19660 18104 19712
rect 19248 19703 19300 19712
rect 19248 19669 19257 19703
rect 19257 19669 19291 19703
rect 19291 19669 19300 19703
rect 19248 19660 19300 19669
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 2688 19320 2740 19372
rect 5540 19456 5592 19508
rect 8300 19456 8352 19508
rect 16948 19499 17000 19508
rect 16948 19465 16957 19499
rect 16957 19465 16991 19499
rect 16991 19465 17000 19499
rect 16948 19456 17000 19465
rect 17224 19456 17276 19508
rect 3332 19363 3384 19372
rect 3332 19329 3341 19363
rect 3341 19329 3375 19363
rect 3375 19329 3384 19363
rect 3332 19320 3384 19329
rect 7748 19388 7800 19440
rect 8392 19388 8444 19440
rect 8668 19388 8720 19440
rect 17960 19388 18012 19440
rect 18144 19388 18196 19440
rect 6920 19252 6972 19304
rect 7288 19295 7340 19304
rect 7288 19261 7297 19295
rect 7297 19261 7331 19295
rect 7331 19261 7340 19295
rect 7288 19252 7340 19261
rect 7656 19252 7708 19304
rect 8208 19252 8260 19304
rect 8576 19252 8628 19304
rect 9496 19295 9548 19304
rect 9496 19261 9505 19295
rect 9505 19261 9539 19295
rect 9539 19261 9548 19295
rect 9496 19252 9548 19261
rect 16672 19320 16724 19372
rect 18696 19320 18748 19372
rect 18972 19320 19024 19372
rect 20168 19320 20220 19372
rect 3056 19184 3108 19236
rect 3700 19184 3752 19236
rect 1768 19159 1820 19168
rect 1768 19125 1777 19159
rect 1777 19125 1811 19159
rect 1811 19125 1820 19159
rect 1768 19116 1820 19125
rect 2136 19159 2188 19168
rect 2136 19125 2145 19159
rect 2145 19125 2179 19159
rect 2179 19125 2188 19159
rect 2136 19116 2188 19125
rect 2688 19116 2740 19168
rect 3148 19116 3200 19168
rect 5724 19184 5776 19236
rect 8484 19184 8536 19236
rect 11060 19184 11112 19236
rect 11520 19252 11572 19304
rect 19248 19295 19300 19304
rect 11980 19184 12032 19236
rect 14556 19184 14608 19236
rect 15476 19184 15528 19236
rect 19248 19261 19257 19295
rect 19257 19261 19291 19295
rect 19291 19261 19300 19295
rect 19248 19252 19300 19261
rect 20076 19252 20128 19304
rect 4252 19116 4304 19168
rect 4896 19116 4948 19168
rect 5816 19159 5868 19168
rect 5816 19125 5825 19159
rect 5825 19125 5859 19159
rect 5859 19125 5868 19159
rect 5816 19116 5868 19125
rect 6828 19159 6880 19168
rect 6828 19125 6837 19159
rect 6837 19125 6871 19159
rect 6871 19125 6880 19159
rect 6828 19116 6880 19125
rect 7196 19159 7248 19168
rect 7196 19125 7205 19159
rect 7205 19125 7239 19159
rect 7239 19125 7248 19159
rect 7196 19116 7248 19125
rect 10784 19116 10836 19168
rect 10968 19116 11020 19168
rect 11704 19116 11756 19168
rect 11796 19116 11848 19168
rect 14004 19116 14056 19168
rect 14648 19116 14700 19168
rect 16580 19184 16632 19236
rect 19800 19184 19852 19236
rect 16304 19116 16356 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 1400 18955 1452 18964
rect 1400 18921 1409 18955
rect 1409 18921 1443 18955
rect 1443 18921 1452 18955
rect 1400 18912 1452 18921
rect 4068 18912 4120 18964
rect 4160 18912 4212 18964
rect 8208 18912 8260 18964
rect 1584 18844 1636 18896
rect 5816 18844 5868 18896
rect 6828 18844 6880 18896
rect 10416 18912 10468 18964
rect 10692 18955 10744 18964
rect 10692 18921 10701 18955
rect 10701 18921 10735 18955
rect 10735 18921 10744 18955
rect 10692 18912 10744 18921
rect 12532 18912 12584 18964
rect 15200 18912 15252 18964
rect 17040 18912 17092 18964
rect 17316 18912 17368 18964
rect 4160 18776 4212 18828
rect 8760 18844 8812 18896
rect 9680 18776 9732 18828
rect 11888 18844 11940 18896
rect 11612 18776 11664 18828
rect 11704 18776 11756 18828
rect 14096 18819 14148 18828
rect 14096 18785 14105 18819
rect 14105 18785 14139 18819
rect 14139 18785 14148 18819
rect 14096 18776 14148 18785
rect 14464 18776 14516 18828
rect 15476 18776 15528 18828
rect 15568 18776 15620 18828
rect 16948 18776 17000 18828
rect 17960 18776 18012 18828
rect 2780 18640 2832 18692
rect 4804 18708 4856 18760
rect 4988 18708 5040 18760
rect 5172 18708 5224 18760
rect 6828 18751 6880 18760
rect 6828 18717 6837 18751
rect 6837 18717 6871 18751
rect 6871 18717 6880 18751
rect 6828 18708 6880 18717
rect 7656 18708 7708 18760
rect 8668 18708 8720 18760
rect 10600 18708 10652 18760
rect 10784 18751 10836 18760
rect 10784 18717 10793 18751
rect 10793 18717 10827 18751
rect 10827 18717 10836 18751
rect 10784 18708 10836 18717
rect 11060 18708 11112 18760
rect 11520 18708 11572 18760
rect 2596 18572 2648 18624
rect 5172 18572 5224 18624
rect 6644 18640 6696 18692
rect 7380 18640 7432 18692
rect 8208 18640 8260 18692
rect 8484 18640 8536 18692
rect 8852 18640 8904 18692
rect 13268 18640 13320 18692
rect 9588 18572 9640 18624
rect 10600 18572 10652 18624
rect 18788 18572 18840 18624
rect 19892 18615 19944 18624
rect 19892 18581 19901 18615
rect 19901 18581 19935 18615
rect 19935 18581 19944 18615
rect 19892 18572 19944 18581
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 2228 18275 2280 18284
rect 2228 18241 2237 18275
rect 2237 18241 2271 18275
rect 2271 18241 2280 18275
rect 2228 18232 2280 18241
rect 4804 18368 4856 18420
rect 11704 18368 11756 18420
rect 12440 18411 12492 18420
rect 12440 18377 12449 18411
rect 12449 18377 12483 18411
rect 12483 18377 12492 18411
rect 12440 18368 12492 18377
rect 13544 18368 13596 18420
rect 15660 18368 15712 18420
rect 17132 18368 17184 18420
rect 10416 18300 10468 18352
rect 10968 18300 11020 18352
rect 3332 18275 3384 18284
rect 3332 18241 3341 18275
rect 3341 18241 3375 18275
rect 3375 18241 3384 18275
rect 3332 18232 3384 18241
rect 6552 18232 6604 18284
rect 1768 18164 1820 18216
rect 3976 18164 4028 18216
rect 3056 18096 3108 18148
rect 4252 18096 4304 18148
rect 5632 18164 5684 18216
rect 5724 18164 5776 18216
rect 204 18028 256 18080
rect 1308 18028 1360 18080
rect 5540 18028 5592 18080
rect 6920 18164 6972 18216
rect 7196 18096 7248 18148
rect 9220 18096 9272 18148
rect 9496 18164 9548 18216
rect 10784 18164 10836 18216
rect 12900 18232 12952 18284
rect 13268 18232 13320 18284
rect 10968 18164 11020 18216
rect 14648 18275 14700 18284
rect 14648 18241 14657 18275
rect 14657 18241 14691 18275
rect 14691 18241 14700 18275
rect 14648 18232 14700 18241
rect 16948 18275 17000 18284
rect 16948 18241 16957 18275
rect 16957 18241 16991 18275
rect 16991 18241 17000 18275
rect 16948 18232 17000 18241
rect 17960 18232 18012 18284
rect 13544 18096 13596 18148
rect 13636 18096 13688 18148
rect 17776 18096 17828 18148
rect 19892 18164 19944 18216
rect 18972 18096 19024 18148
rect 8208 18071 8260 18080
rect 8208 18037 8217 18071
rect 8217 18037 8251 18071
rect 8251 18037 8260 18071
rect 8208 18028 8260 18037
rect 9128 18028 9180 18080
rect 10324 18028 10376 18080
rect 10692 18028 10744 18080
rect 13820 18028 13872 18080
rect 13912 18028 13964 18080
rect 14556 18028 14608 18080
rect 16948 18028 17000 18080
rect 20168 18071 20220 18080
rect 20168 18037 20177 18071
rect 20177 18037 20211 18071
rect 20211 18037 20220 18071
rect 20168 18028 20220 18037
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 4160 17824 4212 17876
rect 7196 17824 7248 17876
rect 9680 17867 9732 17876
rect 3884 17756 3936 17808
rect 4344 17688 4396 17740
rect 4804 17756 4856 17808
rect 5356 17756 5408 17808
rect 6184 17756 6236 17808
rect 6276 17756 6328 17808
rect 6736 17756 6788 17808
rect 8208 17756 8260 17808
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 10232 17824 10284 17876
rect 11704 17824 11756 17876
rect 13268 17824 13320 17876
rect 8116 17688 8168 17740
rect 9956 17688 10008 17740
rect 2412 17620 2464 17672
rect 2504 17620 2556 17672
rect 3056 17663 3108 17672
rect 3056 17629 3065 17663
rect 3065 17629 3099 17663
rect 3099 17629 3108 17663
rect 3056 17620 3108 17629
rect 3332 17620 3384 17672
rect 6552 17620 6604 17672
rect 7656 17620 7708 17672
rect 10140 17620 10192 17672
rect 10416 17756 10468 17808
rect 12716 17756 12768 17808
rect 12900 17756 12952 17808
rect 15200 17756 15252 17808
rect 11888 17731 11940 17740
rect 11888 17697 11922 17731
rect 11922 17697 11940 17731
rect 11888 17688 11940 17697
rect 12348 17688 12400 17740
rect 11060 17620 11112 17672
rect 12808 17688 12860 17740
rect 14372 17688 14424 17740
rect 15936 17756 15988 17808
rect 17592 17756 17644 17808
rect 17960 17688 18012 17740
rect 18604 17688 18656 17740
rect 15016 17620 15068 17672
rect 15200 17620 15252 17672
rect 8484 17552 8536 17604
rect 11520 17552 11572 17604
rect 12624 17552 12676 17604
rect 18788 17552 18840 17604
rect 20536 17620 20588 17672
rect 20812 17620 20864 17672
rect 20444 17552 20496 17604
rect 6828 17484 6880 17536
rect 8116 17484 8168 17536
rect 10232 17484 10284 17536
rect 12532 17484 12584 17536
rect 15200 17484 15252 17536
rect 17684 17527 17736 17536
rect 17684 17493 17693 17527
rect 17693 17493 17727 17527
rect 17727 17493 17736 17527
rect 17684 17484 17736 17493
rect 19156 17484 19208 17536
rect 20812 17484 20864 17536
rect 21824 17484 21876 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 3332 17280 3384 17332
rect 3700 17323 3752 17332
rect 3700 17289 3709 17323
rect 3709 17289 3743 17323
rect 3743 17289 3752 17323
rect 3700 17280 3752 17289
rect 4344 17280 4396 17332
rect 5356 17280 5408 17332
rect 7656 17280 7708 17332
rect 3792 17212 3844 17264
rect 9312 17280 9364 17332
rect 9588 17280 9640 17332
rect 12532 17280 12584 17332
rect 17960 17280 18012 17332
rect 18972 17280 19024 17332
rect 20444 17323 20496 17332
rect 20444 17289 20453 17323
rect 20453 17289 20487 17323
rect 20487 17289 20496 17323
rect 20444 17280 20496 17289
rect 20904 17280 20956 17332
rect 21180 17280 21232 17332
rect 10140 17212 10192 17264
rect 10232 17212 10284 17264
rect 13820 17212 13872 17264
rect 7380 17144 7432 17196
rect 10692 17187 10744 17196
rect 10692 17153 10701 17187
rect 10701 17153 10735 17187
rect 10735 17153 10744 17187
rect 10692 17144 10744 17153
rect 13360 17144 13412 17196
rect 15016 17144 15068 17196
rect 2412 17076 2464 17128
rect 13728 17076 13780 17128
rect 14004 17119 14056 17128
rect 14004 17085 14013 17119
rect 14013 17085 14047 17119
rect 14047 17085 14056 17119
rect 14004 17076 14056 17085
rect 14096 17076 14148 17128
rect 17868 17144 17920 17196
rect 18604 17144 18656 17196
rect 20904 17144 20956 17196
rect 22284 17144 22336 17196
rect 18696 17076 18748 17128
rect 20168 17076 20220 17128
rect 3056 17008 3108 17060
rect 8300 17008 8352 17060
rect 9404 17008 9456 17060
rect 4804 16940 4856 16992
rect 7012 16940 7064 16992
rect 7196 16940 7248 16992
rect 11704 17008 11756 17060
rect 10324 16940 10376 16992
rect 10876 16940 10928 16992
rect 12532 16940 12584 16992
rect 12716 17008 12768 17060
rect 14188 17008 14240 17060
rect 14648 16940 14700 16992
rect 15936 16940 15988 16992
rect 16212 16940 16264 16992
rect 16304 16940 16356 16992
rect 17960 16940 18012 16992
rect 18604 16940 18656 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 2504 16736 2556 16788
rect 4160 16736 4212 16788
rect 10968 16736 11020 16788
rect 11980 16779 12032 16788
rect 11980 16745 11989 16779
rect 11989 16745 12023 16779
rect 12023 16745 12032 16779
rect 11980 16736 12032 16745
rect 12808 16779 12860 16788
rect 12808 16745 12817 16779
rect 12817 16745 12851 16779
rect 12851 16745 12860 16779
rect 12808 16736 12860 16745
rect 2872 16668 2924 16720
rect 1492 16600 1544 16652
rect 5356 16668 5408 16720
rect 6276 16668 6328 16720
rect 13728 16736 13780 16788
rect 19156 16779 19208 16788
rect 19156 16745 19165 16779
rect 19165 16745 19199 16779
rect 19199 16745 19208 16779
rect 19156 16736 19208 16745
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4068 16600 4120 16609
rect 3700 16532 3752 16584
rect 5724 16532 5776 16584
rect 8300 16600 8352 16652
rect 9220 16600 9272 16652
rect 9588 16600 9640 16652
rect 7380 16575 7432 16584
rect 1860 16464 1912 16516
rect 3792 16464 3844 16516
rect 5448 16464 5500 16516
rect 7380 16541 7389 16575
rect 7389 16541 7423 16575
rect 7423 16541 7432 16575
rect 7380 16532 7432 16541
rect 5356 16439 5408 16448
rect 5356 16405 5365 16439
rect 5365 16405 5399 16439
rect 5399 16405 5408 16439
rect 5356 16396 5408 16405
rect 5540 16396 5592 16448
rect 8116 16396 8168 16448
rect 11244 16396 11296 16448
rect 13544 16668 13596 16720
rect 14188 16668 14240 16720
rect 16488 16668 16540 16720
rect 11980 16600 12032 16652
rect 12072 16532 12124 16584
rect 13820 16600 13872 16652
rect 14740 16600 14792 16652
rect 15568 16600 15620 16652
rect 17132 16600 17184 16652
rect 12256 16464 12308 16516
rect 15292 16532 15344 16584
rect 14832 16464 14884 16516
rect 15844 16464 15896 16516
rect 17684 16668 17736 16720
rect 19156 16532 19208 16584
rect 12440 16396 12492 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 3056 16235 3108 16244
rect 3056 16201 3065 16235
rect 3065 16201 3099 16235
rect 3099 16201 3108 16235
rect 3056 16192 3108 16201
rect 7564 16192 7616 16244
rect 8576 16192 8628 16244
rect 11888 16192 11940 16244
rect 9588 16167 9640 16176
rect 9588 16133 9597 16167
rect 9597 16133 9631 16167
rect 9631 16133 9640 16167
rect 9588 16124 9640 16133
rect 10232 16124 10284 16176
rect 3332 15988 3384 16040
rect 10324 16056 10376 16108
rect 15568 16056 15620 16108
rect 15752 16099 15804 16108
rect 15752 16065 15761 16099
rect 15761 16065 15795 16099
rect 15795 16065 15804 16099
rect 15752 16056 15804 16065
rect 19524 16056 19576 16108
rect 20536 16056 20588 16108
rect 5356 15988 5408 16040
rect 8116 15988 8168 16040
rect 8300 15988 8352 16040
rect 10692 15988 10744 16040
rect 12624 15988 12676 16040
rect 3884 15920 3936 15972
rect 4068 15920 4120 15972
rect 1584 15852 1636 15904
rect 2320 15852 2372 15904
rect 4620 15895 4672 15904
rect 4620 15861 4629 15895
rect 4629 15861 4663 15895
rect 4663 15861 4672 15895
rect 4620 15852 4672 15861
rect 5540 15920 5592 15972
rect 7564 15920 7616 15972
rect 10416 15920 10468 15972
rect 10876 15920 10928 15972
rect 12072 15920 12124 15972
rect 14096 15988 14148 16040
rect 18788 16031 18840 16040
rect 18788 15997 18822 16031
rect 18822 15997 18840 16031
rect 18788 15988 18840 15997
rect 14004 15920 14056 15972
rect 16396 15920 16448 15972
rect 14556 15852 14608 15904
rect 15200 15852 15252 15904
rect 15936 15852 15988 15904
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 18788 15852 18840 15904
rect 19340 15920 19392 15972
rect 19156 15852 19208 15904
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 4620 15648 4672 15700
rect 2780 15555 2832 15564
rect 2780 15521 2789 15555
rect 2789 15521 2823 15555
rect 2823 15521 2832 15555
rect 2780 15512 2832 15521
rect 3332 15512 3384 15564
rect 5448 15512 5500 15564
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 8300 15648 8352 15700
rect 8852 15648 8904 15700
rect 9496 15648 9548 15700
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 12440 15648 12492 15700
rect 14004 15648 14056 15700
rect 14372 15691 14424 15700
rect 14372 15657 14381 15691
rect 14381 15657 14415 15691
rect 14415 15657 14424 15691
rect 14372 15648 14424 15657
rect 15292 15648 15344 15700
rect 6828 15580 6880 15632
rect 10784 15580 10836 15632
rect 11152 15580 11204 15632
rect 11888 15580 11940 15632
rect 7104 15512 7156 15564
rect 8944 15512 8996 15564
rect 11520 15512 11572 15564
rect 12072 15512 12124 15564
rect 13084 15512 13136 15564
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 10692 15444 10744 15496
rect 12164 15444 12216 15496
rect 18052 15580 18104 15632
rect 15568 15512 15620 15564
rect 17684 15512 17736 15564
rect 19340 15512 19392 15564
rect 7472 15376 7524 15428
rect 13544 15444 13596 15496
rect 14372 15444 14424 15496
rect 20260 15444 20312 15496
rect 1952 15308 2004 15360
rect 3884 15308 3936 15360
rect 6184 15308 6236 15360
rect 9312 15308 9364 15360
rect 11060 15308 11112 15360
rect 16396 15308 16448 15360
rect 19616 15308 19668 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 2780 15104 2832 15156
rect 6092 15104 6144 15156
rect 6552 15104 6604 15156
rect 7748 15036 7800 15088
rect 3884 15011 3936 15020
rect 3884 14977 3893 15011
rect 3893 14977 3927 15011
rect 3927 14977 3936 15011
rect 3884 14968 3936 14977
rect 5448 15011 5500 15020
rect 5448 14977 5457 15011
rect 5457 14977 5491 15011
rect 5491 14977 5500 15011
rect 5448 14968 5500 14977
rect 7380 15011 7432 15020
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7380 14968 7432 14977
rect 6552 14900 6604 14952
rect 7104 14900 7156 14952
rect 16304 15147 16356 15156
rect 16304 15113 16313 15147
rect 16313 15113 16347 15147
rect 16347 15113 16356 15147
rect 16304 15104 16356 15113
rect 11152 15036 11204 15088
rect 12256 15036 12308 15088
rect 14096 15036 14148 15088
rect 14372 15036 14424 15088
rect 18788 15036 18840 15088
rect 8852 14968 8904 15020
rect 10692 14968 10744 15020
rect 9588 14900 9640 14952
rect 11244 14943 11296 14952
rect 11244 14909 11253 14943
rect 11253 14909 11287 14943
rect 11287 14909 11296 14943
rect 11244 14900 11296 14909
rect 12440 14968 12492 15020
rect 13544 14968 13596 15020
rect 2320 14764 2372 14816
rect 3700 14807 3752 14816
rect 3700 14773 3709 14807
rect 3709 14773 3743 14807
rect 3743 14773 3752 14807
rect 3700 14764 3752 14773
rect 4988 14764 5040 14816
rect 5540 14764 5592 14816
rect 11060 14832 11112 14884
rect 8392 14764 8444 14816
rect 11336 14764 11388 14816
rect 12440 14764 12492 14816
rect 13176 14832 13228 14884
rect 13452 14764 13504 14816
rect 18788 14900 18840 14952
rect 19156 14943 19208 14952
rect 19156 14909 19190 14943
rect 19190 14909 19208 14943
rect 19156 14900 19208 14909
rect 16948 14832 17000 14884
rect 17316 14764 17368 14816
rect 20260 14807 20312 14816
rect 20260 14773 20269 14807
rect 20269 14773 20303 14807
rect 20303 14773 20312 14807
rect 20260 14764 20312 14773
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 2872 14603 2924 14612
rect 2872 14569 2881 14603
rect 2881 14569 2915 14603
rect 2915 14569 2924 14603
rect 2872 14560 2924 14569
rect 3700 14560 3752 14612
rect 6552 14560 6604 14612
rect 14004 14560 14056 14612
rect 14372 14560 14424 14612
rect 19340 14560 19392 14612
rect 19616 14603 19668 14612
rect 19616 14569 19625 14603
rect 19625 14569 19659 14603
rect 19659 14569 19668 14603
rect 19616 14560 19668 14569
rect 7472 14492 7524 14544
rect 9036 14492 9088 14544
rect 12716 14492 12768 14544
rect 15568 14492 15620 14544
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 3792 14424 3844 14476
rect 5448 14424 5500 14476
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 2688 14356 2740 14408
rect 3424 14356 3476 14408
rect 4896 14356 4948 14408
rect 5356 14356 5408 14408
rect 2504 14288 2556 14340
rect 3700 14288 3752 14340
rect 4988 14288 5040 14340
rect 9496 14424 9548 14476
rect 9680 14467 9732 14476
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 11152 14424 11204 14476
rect 12440 14424 12492 14476
rect 13360 14424 13412 14476
rect 14096 14467 14148 14476
rect 14096 14433 14105 14467
rect 14105 14433 14139 14467
rect 14139 14433 14148 14467
rect 14096 14424 14148 14433
rect 15752 14424 15804 14476
rect 17040 14424 17092 14476
rect 8852 14356 8904 14408
rect 11060 14356 11112 14408
rect 11612 14356 11664 14408
rect 14372 14356 14424 14408
rect 14556 14356 14608 14408
rect 19708 14399 19760 14408
rect 19708 14365 19717 14399
rect 19717 14365 19751 14399
rect 19751 14365 19760 14399
rect 19708 14356 19760 14365
rect 20168 14356 20220 14408
rect 9496 14288 9548 14340
rect 6000 14220 6052 14272
rect 7380 14220 7432 14272
rect 11244 14220 11296 14272
rect 13452 14288 13504 14340
rect 13728 14288 13780 14340
rect 17684 14331 17736 14340
rect 17684 14297 17693 14331
rect 17693 14297 17727 14331
rect 17727 14297 17736 14331
rect 17684 14288 17736 14297
rect 13176 14220 13228 14272
rect 13360 14220 13412 14272
rect 16120 14220 16172 14272
rect 18144 14220 18196 14272
rect 18788 14220 18840 14272
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 6092 14016 6144 14068
rect 6552 14016 6604 14068
rect 4896 13948 4948 14000
rect 5080 13948 5132 14000
rect 5540 13948 5592 14000
rect 7840 14016 7892 14068
rect 9036 14059 9088 14068
rect 9036 14025 9045 14059
rect 9045 14025 9079 14059
rect 9079 14025 9088 14059
rect 9036 14016 9088 14025
rect 14004 14059 14056 14068
rect 9312 13948 9364 14000
rect 2228 13855 2280 13864
rect 2228 13821 2237 13855
rect 2237 13821 2271 13855
rect 2271 13821 2280 13855
rect 2228 13812 2280 13821
rect 3332 13855 3384 13864
rect 3332 13821 3341 13855
rect 3341 13821 3375 13855
rect 3375 13821 3384 13855
rect 3332 13812 3384 13821
rect 3424 13812 3476 13864
rect 4068 13812 4120 13864
rect 6184 13880 6236 13932
rect 10692 13948 10744 14000
rect 11704 13948 11756 14000
rect 12164 13948 12216 14000
rect 11336 13923 11388 13932
rect 11336 13889 11345 13923
rect 11345 13889 11379 13923
rect 11379 13889 11388 13923
rect 11336 13880 11388 13889
rect 5908 13812 5960 13864
rect 7380 13812 7432 13864
rect 12716 13880 12768 13932
rect 14004 14025 14013 14059
rect 14013 14025 14047 14059
rect 14047 14025 14056 14059
rect 14004 14016 14056 14025
rect 15568 14059 15620 14068
rect 15568 14025 15577 14059
rect 15577 14025 15611 14059
rect 15611 14025 15620 14059
rect 15568 14016 15620 14025
rect 16120 14016 16172 14068
rect 17960 14016 18012 14068
rect 13452 13948 13504 14000
rect 18788 13948 18840 14000
rect 13176 13880 13228 13932
rect 15568 13880 15620 13932
rect 16028 13880 16080 13932
rect 17500 13880 17552 13932
rect 12900 13855 12952 13864
rect 2504 13744 2556 13796
rect 2872 13744 2924 13796
rect 5540 13676 5592 13728
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 13820 13812 13872 13864
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 18144 13812 18196 13864
rect 8300 13744 8352 13796
rect 10508 13744 10560 13796
rect 11152 13787 11204 13796
rect 11152 13753 11161 13787
rect 11161 13753 11195 13787
rect 11195 13753 11204 13787
rect 11152 13744 11204 13753
rect 11888 13744 11940 13796
rect 12716 13744 12768 13796
rect 20260 13812 20312 13864
rect 19524 13744 19576 13796
rect 8760 13676 8812 13728
rect 9036 13676 9088 13728
rect 9588 13676 9640 13728
rect 9864 13676 9916 13728
rect 12992 13676 13044 13728
rect 16396 13719 16448 13728
rect 16396 13685 16405 13719
rect 16405 13685 16439 13719
rect 16439 13685 16448 13719
rect 16396 13676 16448 13685
rect 16764 13719 16816 13728
rect 16764 13685 16773 13719
rect 16773 13685 16807 13719
rect 16807 13685 16816 13719
rect 16764 13676 16816 13685
rect 20168 13719 20220 13728
rect 20168 13685 20177 13719
rect 20177 13685 20211 13719
rect 20211 13685 20220 13719
rect 20168 13676 20220 13685
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 6092 13515 6144 13524
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 7104 13472 7156 13524
rect 10692 13472 10744 13524
rect 10968 13472 11020 13524
rect 2596 13404 2648 13456
rect 3332 13404 3384 13456
rect 6000 13447 6052 13456
rect 6000 13413 6009 13447
rect 6009 13413 6043 13447
rect 6043 13413 6052 13447
rect 6000 13404 6052 13413
rect 3056 13336 3108 13388
rect 3148 13336 3200 13388
rect 4344 13336 4396 13388
rect 5724 13336 5776 13388
rect 6000 13268 6052 13320
rect 11336 13404 11388 13456
rect 11520 13447 11572 13456
rect 11520 13413 11554 13447
rect 11554 13413 11572 13447
rect 11520 13404 11572 13413
rect 6276 13311 6328 13320
rect 6276 13277 6285 13311
rect 6285 13277 6319 13311
rect 6319 13277 6328 13311
rect 6276 13268 6328 13277
rect 9864 13336 9916 13388
rect 10692 13336 10744 13388
rect 16396 13472 16448 13524
rect 18052 13404 18104 13456
rect 7656 13200 7708 13252
rect 8760 13268 8812 13320
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 9036 13200 9088 13252
rect 9312 13200 9364 13252
rect 12624 13336 12676 13388
rect 13544 13336 13596 13388
rect 11060 13268 11112 13320
rect 17408 13336 17460 13388
rect 17684 13379 17736 13388
rect 17684 13345 17693 13379
rect 17693 13345 17727 13379
rect 17727 13345 17736 13379
rect 17684 13336 17736 13345
rect 17960 13379 18012 13388
rect 17960 13345 17994 13379
rect 17994 13345 18012 13379
rect 17960 13336 18012 13345
rect 18788 13336 18840 13388
rect 14004 13311 14056 13320
rect 2872 13132 2924 13184
rect 4068 13175 4120 13184
rect 4068 13141 4077 13175
rect 4077 13141 4111 13175
rect 4111 13141 4120 13175
rect 4068 13132 4120 13141
rect 5816 13132 5868 13184
rect 8300 13132 8352 13184
rect 14004 13277 14013 13311
rect 14013 13277 14047 13311
rect 14047 13277 14056 13311
rect 14004 13268 14056 13277
rect 12440 13132 12492 13184
rect 13176 13132 13228 13184
rect 13452 13175 13504 13184
rect 13452 13141 13461 13175
rect 13461 13141 13495 13175
rect 13495 13141 13504 13175
rect 13452 13132 13504 13141
rect 15200 13132 15252 13184
rect 17960 13132 18012 13184
rect 19340 13132 19392 13184
rect 19616 13132 19668 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 5724 12928 5776 12980
rect 2596 12792 2648 12844
rect 6276 12792 6328 12844
rect 10232 12928 10284 12980
rect 10692 12971 10744 12980
rect 10692 12937 10701 12971
rect 10701 12937 10735 12971
rect 10735 12937 10744 12971
rect 10692 12928 10744 12937
rect 11796 12928 11848 12980
rect 12072 12928 12124 12980
rect 14096 12928 14148 12980
rect 17040 12928 17092 12980
rect 18788 12928 18840 12980
rect 10416 12860 10468 12912
rect 11888 12860 11940 12912
rect 14464 12860 14516 12912
rect 18328 12860 18380 12912
rect 19340 12860 19392 12912
rect 11244 12835 11296 12844
rect 2412 12724 2464 12776
rect 4252 12724 4304 12776
rect 5080 12724 5132 12776
rect 5448 12767 5500 12776
rect 5448 12733 5457 12767
rect 5457 12733 5491 12767
rect 5491 12733 5500 12767
rect 5448 12724 5500 12733
rect 5540 12767 5592 12776
rect 5540 12733 5549 12767
rect 5549 12733 5583 12767
rect 5583 12733 5592 12767
rect 5540 12724 5592 12733
rect 8760 12767 8812 12776
rect 8760 12733 8794 12767
rect 8794 12733 8812 12767
rect 11244 12801 11253 12835
rect 11253 12801 11287 12835
rect 11287 12801 11296 12835
rect 11244 12792 11296 12801
rect 12624 12792 12676 12844
rect 12716 12792 12768 12844
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 15752 12835 15804 12844
rect 15752 12801 15761 12835
rect 15761 12801 15795 12835
rect 15795 12801 15804 12835
rect 15752 12792 15804 12801
rect 11060 12767 11112 12776
rect 1860 12699 1912 12708
rect 1860 12665 1869 12699
rect 1869 12665 1903 12699
rect 1903 12665 1912 12699
rect 1860 12656 1912 12665
rect 2504 12588 2556 12640
rect 3056 12588 3108 12640
rect 4712 12656 4764 12708
rect 6736 12656 6788 12708
rect 8760 12724 8812 12733
rect 11060 12733 11069 12767
rect 11069 12733 11103 12767
rect 11103 12733 11112 12767
rect 11060 12724 11112 12733
rect 9680 12656 9732 12708
rect 9772 12656 9824 12708
rect 13452 12724 13504 12776
rect 18696 12724 18748 12776
rect 18880 12724 18932 12776
rect 19156 12724 19208 12776
rect 11428 12656 11480 12708
rect 13268 12656 13320 12708
rect 15292 12656 15344 12708
rect 18236 12656 18288 12708
rect 18604 12656 18656 12708
rect 19984 12656 20036 12708
rect 10508 12588 10560 12640
rect 10692 12588 10744 12640
rect 12440 12631 12492 12640
rect 12440 12597 12449 12631
rect 12449 12597 12483 12631
rect 12483 12597 12492 12631
rect 12808 12631 12860 12640
rect 12440 12588 12492 12597
rect 12808 12597 12817 12631
rect 12817 12597 12851 12631
rect 12851 12597 12860 12631
rect 12808 12588 12860 12597
rect 12992 12588 13044 12640
rect 14096 12588 14148 12640
rect 18512 12588 18564 12640
rect 19524 12588 19576 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 4068 12384 4120 12436
rect 6276 12427 6328 12436
rect 6276 12393 6285 12427
rect 6285 12393 6319 12427
rect 6319 12393 6328 12427
rect 6276 12384 6328 12393
rect 7196 12384 7248 12436
rect 7472 12384 7524 12436
rect 11060 12384 11112 12436
rect 11336 12384 11388 12436
rect 12072 12384 12124 12436
rect 14004 12384 14056 12436
rect 3424 12316 3476 12368
rect 6552 12316 6604 12368
rect 8392 12359 8444 12368
rect 8392 12325 8401 12359
rect 8401 12325 8435 12359
rect 8435 12325 8444 12359
rect 8392 12316 8444 12325
rect 8668 12316 8720 12368
rect 9496 12316 9548 12368
rect 2228 12248 2280 12300
rect 3332 12248 3384 12300
rect 7196 12248 7248 12300
rect 7748 12248 7800 12300
rect 8208 12248 8260 12300
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 10048 12316 10100 12368
rect 10232 12316 10284 12368
rect 10784 12316 10836 12368
rect 11704 12316 11756 12368
rect 2872 12223 2924 12232
rect 2872 12189 2881 12223
rect 2881 12189 2915 12223
rect 2915 12189 2924 12223
rect 2872 12180 2924 12189
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 9128 12180 9180 12232
rect 12256 12180 12308 12232
rect 13820 12248 13872 12300
rect 14832 12248 14884 12300
rect 15844 12316 15896 12368
rect 17224 12316 17276 12368
rect 19064 12384 19116 12436
rect 20076 12384 20128 12436
rect 19340 12316 19392 12368
rect 16120 12291 16172 12300
rect 16120 12257 16129 12291
rect 16129 12257 16163 12291
rect 16163 12257 16172 12291
rect 16120 12248 16172 12257
rect 3424 12112 3476 12164
rect 3700 12112 3752 12164
rect 4620 12112 4672 12164
rect 7656 12112 7708 12164
rect 8668 12112 8720 12164
rect 11152 12112 11204 12164
rect 11336 12112 11388 12164
rect 12624 12112 12676 12164
rect 4068 12044 4120 12096
rect 6920 12044 6972 12096
rect 10048 12044 10100 12096
rect 15752 12180 15804 12232
rect 13084 12044 13136 12096
rect 13176 12044 13228 12096
rect 13728 12044 13780 12096
rect 14096 12044 14148 12096
rect 14556 12044 14608 12096
rect 14832 12087 14884 12096
rect 14832 12053 14841 12087
rect 14841 12053 14875 12087
rect 14875 12053 14884 12087
rect 14832 12044 14884 12053
rect 15844 12044 15896 12096
rect 16120 12044 16172 12096
rect 18512 12248 18564 12300
rect 20628 12248 20680 12300
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 19984 12087 20036 12096
rect 19984 12053 19993 12087
rect 19993 12053 20027 12087
rect 20027 12053 20036 12087
rect 19984 12044 20036 12053
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 2228 11883 2280 11892
rect 2228 11849 2237 11883
rect 2237 11849 2271 11883
rect 2271 11849 2280 11883
rect 2228 11840 2280 11849
rect 2504 11704 2556 11756
rect 3148 11704 3200 11756
rect 8208 11840 8260 11892
rect 9312 11883 9364 11892
rect 9312 11849 9321 11883
rect 9321 11849 9355 11883
rect 9355 11849 9364 11883
rect 9312 11840 9364 11849
rect 11060 11840 11112 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 16764 11840 16816 11892
rect 17960 11840 18012 11892
rect 18696 11840 18748 11892
rect 19708 11840 19760 11892
rect 4252 11704 4304 11756
rect 6644 11704 6696 11756
rect 9772 11704 9824 11756
rect 9956 11747 10008 11756
rect 9956 11713 9965 11747
rect 9965 11713 9999 11747
rect 9999 11713 10008 11747
rect 9956 11704 10008 11713
rect 10048 11704 10100 11756
rect 6920 11636 6972 11688
rect 2964 11568 3016 11620
rect 3976 11568 4028 11620
rect 5264 11568 5316 11620
rect 5540 11568 5592 11620
rect 6644 11568 6696 11620
rect 10232 11636 10284 11688
rect 10416 11679 10468 11688
rect 10416 11645 10450 11679
rect 10450 11645 10468 11679
rect 10416 11636 10468 11645
rect 3700 11500 3752 11552
rect 7748 11500 7800 11552
rect 9220 11500 9272 11552
rect 13084 11636 13136 11688
rect 13452 11636 13504 11688
rect 12716 11611 12768 11620
rect 12716 11577 12750 11611
rect 12750 11577 12768 11611
rect 12716 11568 12768 11577
rect 13728 11568 13780 11620
rect 9864 11500 9916 11552
rect 11612 11543 11664 11552
rect 11612 11509 11621 11543
rect 11621 11509 11655 11543
rect 11655 11509 11664 11543
rect 11612 11500 11664 11509
rect 13084 11500 13136 11552
rect 15016 11679 15068 11688
rect 15016 11645 15025 11679
rect 15025 11645 15059 11679
rect 15059 11645 15068 11679
rect 15016 11636 15068 11645
rect 16580 11636 16632 11688
rect 17040 11636 17092 11688
rect 14280 11568 14332 11620
rect 14556 11568 14608 11620
rect 16488 11568 16540 11620
rect 19984 11704 20036 11756
rect 20260 11747 20312 11756
rect 20260 11713 20269 11747
rect 20269 11713 20303 11747
rect 20303 11713 20312 11747
rect 20260 11704 20312 11713
rect 20352 11568 20404 11620
rect 14464 11500 14516 11552
rect 16672 11500 16724 11552
rect 17040 11500 17092 11552
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 19156 11500 19208 11552
rect 20076 11543 20128 11552
rect 20076 11509 20085 11543
rect 20085 11509 20119 11543
rect 20119 11509 20128 11543
rect 20076 11500 20128 11509
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 6552 11296 6604 11348
rect 6828 11296 6880 11348
rect 7104 11296 7156 11348
rect 8576 11296 8628 11348
rect 9772 11296 9824 11348
rect 12256 11296 12308 11348
rect 16488 11296 16540 11348
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 19432 11296 19484 11348
rect 19708 11296 19760 11348
rect 4528 11228 4580 11280
rect 10232 11228 10284 11280
rect 14004 11228 14056 11280
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 4712 11160 4764 11212
rect 6184 11160 6236 11212
rect 6920 11160 6972 11212
rect 1860 11092 1912 11144
rect 2412 11092 2464 11144
rect 3148 11092 3200 11144
rect 4712 11024 4764 11076
rect 2412 10999 2464 11008
rect 2412 10965 2421 10999
rect 2421 10965 2455 10999
rect 2455 10965 2464 10999
rect 2412 10956 2464 10965
rect 5540 10956 5592 11008
rect 5724 10956 5776 11008
rect 8668 11160 8720 11212
rect 9956 11160 10008 11212
rect 12440 11160 12492 11212
rect 15200 11160 15252 11212
rect 16672 11228 16724 11280
rect 17500 11228 17552 11280
rect 17868 11228 17920 11280
rect 19984 11228 20036 11280
rect 7748 11024 7800 11076
rect 9496 11092 9548 11144
rect 11152 11092 11204 11144
rect 8760 11024 8812 11076
rect 12256 11024 12308 11076
rect 13820 11092 13872 11144
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 19248 11160 19300 11212
rect 15292 11067 15344 11076
rect 15292 11033 15301 11067
rect 15301 11033 15335 11067
rect 15335 11033 15344 11067
rect 15292 11024 15344 11033
rect 17132 11024 17184 11076
rect 19432 11092 19484 11144
rect 20260 11092 20312 11144
rect 7564 10999 7616 11008
rect 7564 10965 7573 10999
rect 7573 10965 7607 10999
rect 7607 10965 7616 10999
rect 7564 10956 7616 10965
rect 8576 10956 8628 11008
rect 9312 10956 9364 11008
rect 15384 10956 15436 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 1124 10752 1176 10804
rect 1492 10752 1544 10804
rect 8484 10752 8536 10804
rect 9128 10752 9180 10804
rect 9496 10752 9548 10804
rect 10416 10752 10468 10804
rect 12808 10752 12860 10804
rect 2688 10684 2740 10736
rect 4068 10684 4120 10736
rect 2504 10616 2556 10668
rect 3148 10616 3200 10668
rect 3976 10616 4028 10668
rect 2412 10548 2464 10600
rect 3332 10548 3384 10600
rect 3700 10548 3752 10600
rect 8576 10684 8628 10736
rect 5724 10616 5776 10668
rect 5540 10548 5592 10600
rect 7564 10616 7616 10668
rect 8484 10616 8536 10668
rect 12716 10684 12768 10736
rect 17684 10752 17736 10804
rect 20076 10752 20128 10804
rect 20628 10752 20680 10804
rect 13084 10616 13136 10668
rect 8392 10548 8444 10600
rect 8760 10548 8812 10600
rect 10140 10548 10192 10600
rect 14280 10616 14332 10668
rect 14464 10659 14516 10668
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 14832 10616 14884 10668
rect 15752 10684 15804 10736
rect 18236 10684 18288 10736
rect 9128 10523 9180 10532
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 3240 10455 3292 10464
rect 3240 10421 3249 10455
rect 3249 10421 3283 10455
rect 3283 10421 3292 10455
rect 3240 10412 3292 10421
rect 3700 10455 3752 10464
rect 3700 10421 3709 10455
rect 3709 10421 3743 10455
rect 3743 10421 3752 10455
rect 9128 10489 9140 10523
rect 9140 10489 9180 10523
rect 9128 10480 9180 10489
rect 9680 10480 9732 10532
rect 12348 10480 12400 10532
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 19248 10548 19300 10600
rect 14464 10480 14516 10532
rect 15568 10480 15620 10532
rect 16488 10480 16540 10532
rect 19892 10480 19944 10532
rect 21088 10480 21140 10532
rect 22744 10480 22796 10532
rect 3700 10412 3752 10421
rect 7104 10412 7156 10464
rect 7288 10455 7340 10464
rect 7288 10421 7297 10455
rect 7297 10421 7331 10455
rect 7331 10421 7340 10455
rect 7288 10412 7340 10421
rect 7472 10412 7524 10464
rect 9312 10412 9364 10464
rect 12440 10412 12492 10464
rect 13084 10412 13136 10464
rect 13268 10412 13320 10464
rect 14004 10455 14056 10464
rect 14004 10421 14013 10455
rect 14013 10421 14047 10455
rect 14047 10421 14056 10455
rect 14004 10412 14056 10421
rect 15752 10412 15804 10464
rect 17132 10455 17184 10464
rect 17132 10421 17141 10455
rect 17141 10421 17175 10455
rect 17175 10421 17184 10455
rect 17132 10412 17184 10421
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 1676 10208 1728 10260
rect 3976 10208 4028 10260
rect 8484 10251 8536 10260
rect 8484 10217 8493 10251
rect 8493 10217 8527 10251
rect 8527 10217 8536 10251
rect 8484 10208 8536 10217
rect 8668 10208 8720 10260
rect 12348 10251 12400 10260
rect 2780 10140 2832 10192
rect 3424 10140 3476 10192
rect 3700 10072 3752 10124
rect 5540 10140 5592 10192
rect 5724 10140 5776 10192
rect 7748 10140 7800 10192
rect 10876 10140 10928 10192
rect 12348 10217 12357 10251
rect 12357 10217 12391 10251
rect 12391 10217 12400 10251
rect 12348 10208 12400 10217
rect 12440 10208 12492 10260
rect 13820 10208 13872 10260
rect 16120 10208 16172 10260
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 12900 10140 12952 10192
rect 13268 10140 13320 10192
rect 15568 10140 15620 10192
rect 15752 10140 15804 10192
rect 16580 10140 16632 10192
rect 18696 10140 18748 10192
rect 6552 10072 6604 10124
rect 6644 10072 6696 10124
rect 10784 10115 10836 10124
rect 10784 10081 10793 10115
rect 10793 10081 10827 10115
rect 10827 10081 10836 10115
rect 10784 10072 10836 10081
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 8300 10004 8352 10056
rect 12624 10072 12676 10124
rect 14004 10072 14056 10124
rect 12348 10004 12400 10056
rect 15752 10004 15804 10056
rect 17132 10072 17184 10124
rect 18052 10072 18104 10124
rect 19248 10072 19300 10124
rect 572 9936 624 9988
rect 4528 9936 4580 9988
rect 1768 9868 1820 9920
rect 2780 9868 2832 9920
rect 6184 9911 6236 9920
rect 6184 9877 6193 9911
rect 6193 9877 6227 9911
rect 6227 9877 6236 9911
rect 6184 9868 6236 9877
rect 12716 9936 12768 9988
rect 10416 9911 10468 9920
rect 10416 9877 10425 9911
rect 10425 9877 10459 9911
rect 10459 9877 10468 9911
rect 10416 9868 10468 9877
rect 10508 9868 10560 9920
rect 11060 9868 11112 9920
rect 12624 9911 12676 9920
rect 12624 9877 12633 9911
rect 12633 9877 12667 9911
rect 12667 9877 12676 9911
rect 12624 9868 12676 9877
rect 12808 9868 12860 9920
rect 17868 9936 17920 9988
rect 19892 9868 19944 9920
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 2688 9664 2740 9716
rect 3700 9707 3752 9716
rect 1216 9596 1268 9648
rect 1492 9596 1544 9648
rect 2504 9596 2556 9648
rect 3700 9673 3709 9707
rect 3709 9673 3743 9707
rect 3743 9673 3752 9707
rect 3700 9664 3752 9673
rect 4068 9664 4120 9716
rect 9128 9707 9180 9716
rect 3976 9596 4028 9648
rect 9128 9673 9137 9707
rect 9137 9673 9171 9707
rect 9171 9673 9180 9707
rect 9128 9664 9180 9673
rect 12808 9664 12860 9716
rect 12900 9664 12952 9716
rect 16488 9664 16540 9716
rect 16580 9664 16632 9716
rect 11520 9596 11572 9648
rect 6644 9528 6696 9580
rect 7564 9528 7616 9580
rect 10416 9528 10468 9580
rect 1492 9503 1544 9512
rect 1492 9469 1501 9503
rect 1501 9469 1535 9503
rect 1535 9469 1544 9503
rect 1492 9460 1544 9469
rect 3240 9460 3292 9512
rect 5172 9460 5224 9512
rect 7748 9503 7800 9512
rect 7748 9469 7757 9503
rect 7757 9469 7791 9503
rect 7791 9469 7800 9503
rect 7748 9460 7800 9469
rect 12808 9460 12860 9512
rect 13452 9460 13504 9512
rect 14464 9460 14516 9512
rect 19984 9664 20036 9716
rect 20444 9664 20496 9716
rect 20720 9664 20772 9716
rect 21088 9664 21140 9716
rect 21180 9664 21232 9716
rect 21364 9664 21416 9716
rect 15936 9528 15988 9580
rect 18052 9571 18104 9580
rect 18052 9537 18061 9571
rect 18061 9537 18095 9571
rect 18095 9537 18104 9571
rect 18052 9528 18104 9537
rect 15292 9460 15344 9512
rect 20260 9503 20312 9512
rect 20260 9469 20269 9503
rect 20269 9469 20303 9503
rect 20303 9469 20312 9503
rect 20260 9460 20312 9469
rect 2688 9392 2740 9444
rect 5908 9392 5960 9444
rect 3240 9324 3292 9376
rect 7288 9324 7340 9376
rect 7564 9392 7616 9444
rect 10692 9392 10744 9444
rect 11060 9392 11112 9444
rect 10416 9324 10468 9376
rect 11888 9324 11940 9376
rect 15200 9392 15252 9444
rect 15844 9392 15896 9444
rect 17684 9392 17736 9444
rect 19984 9392 20036 9444
rect 15384 9324 15436 9376
rect 16120 9367 16172 9376
rect 16120 9333 16129 9367
rect 16129 9333 16163 9367
rect 16163 9333 16172 9367
rect 16120 9324 16172 9333
rect 16764 9324 16816 9376
rect 17316 9324 17368 9376
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 1492 9120 1544 9172
rect 2872 9120 2924 9172
rect 4252 9163 4304 9172
rect 4252 9129 4261 9163
rect 4261 9129 4295 9163
rect 4295 9129 4304 9163
rect 4252 9120 4304 9129
rect 2504 8984 2556 9036
rect 3976 8984 4028 9036
rect 5908 9120 5960 9172
rect 6552 9163 6604 9172
rect 6552 9129 6561 9163
rect 6561 9129 6595 9163
rect 6595 9129 6604 9163
rect 6552 9120 6604 9129
rect 8300 9120 8352 9172
rect 8392 9120 8444 9172
rect 9036 9120 9088 9172
rect 9128 9120 9180 9172
rect 9496 9120 9548 9172
rect 10048 9120 10100 9172
rect 10692 9120 10744 9172
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 11888 9163 11940 9172
rect 11888 9129 11897 9163
rect 11897 9129 11931 9163
rect 11931 9129 11940 9163
rect 11888 9120 11940 9129
rect 15660 9120 15712 9172
rect 17316 9120 17368 9172
rect 17592 9120 17644 9172
rect 19156 9120 19208 9172
rect 19616 9163 19668 9172
rect 19616 9129 19625 9163
rect 19625 9129 19659 9163
rect 19659 9129 19668 9163
rect 19616 9120 19668 9129
rect 4988 9052 5040 9104
rect 5172 9052 5224 9104
rect 5540 9052 5592 9104
rect 2780 8916 2832 8968
rect 2964 8916 3016 8968
rect 4252 8916 4304 8968
rect 4804 8916 4856 8968
rect 5724 8984 5776 9036
rect 8576 9052 8628 9104
rect 8392 9027 8444 9036
rect 8392 8993 8401 9027
rect 8401 8993 8435 9027
rect 8435 8993 8444 9027
rect 8392 8984 8444 8993
rect 12072 9052 12124 9104
rect 12624 9052 12676 9104
rect 12716 9052 12768 9104
rect 9312 8984 9364 9036
rect 11612 8984 11664 9036
rect 15936 9052 15988 9104
rect 16488 9052 16540 9104
rect 18236 9052 18288 9104
rect 19708 9052 19760 9104
rect 15292 9027 15344 9036
rect 15292 8993 15301 9027
rect 15301 8993 15335 9027
rect 15335 8993 15344 9027
rect 15292 8984 15344 8993
rect 17592 8984 17644 9036
rect 2964 8780 3016 8832
rect 7380 8916 7432 8968
rect 8576 8916 8628 8968
rect 9588 8916 9640 8968
rect 10876 8916 10928 8968
rect 9036 8848 9088 8900
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 7748 8780 7800 8789
rect 8760 8780 8812 8832
rect 15844 8916 15896 8968
rect 19708 8959 19760 8968
rect 19708 8925 19717 8959
rect 19717 8925 19751 8959
rect 19751 8925 19760 8959
rect 19708 8916 19760 8925
rect 18236 8848 18288 8900
rect 19616 8848 19668 8900
rect 12716 8780 12768 8832
rect 13728 8780 13780 8832
rect 14280 8780 14332 8832
rect 15660 8780 15712 8832
rect 17684 8780 17736 8832
rect 20076 8916 20128 8968
rect 20076 8780 20128 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 2964 8576 3016 8628
rect 3516 8576 3568 8628
rect 2964 8440 3016 8492
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 5540 8576 5592 8628
rect 6736 8576 6788 8628
rect 7564 8508 7616 8560
rect 5632 8483 5684 8492
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 5632 8440 5684 8449
rect 6828 8440 6880 8492
rect 7104 8372 7156 8424
rect 10324 8576 10376 8628
rect 10876 8576 10928 8628
rect 12256 8508 12308 8560
rect 12624 8508 12676 8560
rect 12900 8508 12952 8560
rect 8760 8440 8812 8492
rect 8576 8372 8628 8424
rect 9036 8372 9088 8424
rect 9312 8372 9364 8424
rect 15292 8576 15344 8628
rect 15660 8576 15712 8628
rect 18880 8576 18932 8628
rect 15568 8508 15620 8560
rect 16120 8440 16172 8492
rect 18052 8508 18104 8560
rect 19156 8483 19208 8492
rect 19156 8449 19165 8483
rect 19165 8449 19199 8483
rect 19199 8449 19208 8483
rect 19156 8440 19208 8449
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 12440 8372 12492 8381
rect 2872 8304 2924 8356
rect 4068 8304 4120 8356
rect 8760 8304 8812 8356
rect 9588 8304 9640 8356
rect 11336 8304 11388 8356
rect 13452 8372 13504 8424
rect 14464 8372 14516 8424
rect 12900 8304 12952 8356
rect 13176 8304 13228 8356
rect 15292 8304 15344 8356
rect 8484 8236 8536 8288
rect 9036 8236 9088 8288
rect 12348 8236 12400 8288
rect 13268 8236 13320 8288
rect 13452 8236 13504 8288
rect 14280 8236 14332 8288
rect 17224 8372 17276 8424
rect 20168 8372 20220 8424
rect 20536 8372 20588 8424
rect 20904 8372 20956 8424
rect 17132 8236 17184 8288
rect 17776 8236 17828 8288
rect 20168 8236 20220 8288
rect 20352 8236 20404 8288
rect 20536 8279 20588 8288
rect 20536 8245 20545 8279
rect 20545 8245 20579 8279
rect 20579 8245 20588 8279
rect 20536 8236 20588 8245
rect 20628 8236 20680 8288
rect 21456 8236 21508 8288
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 10508 8032 10560 8084
rect 10784 8075 10836 8084
rect 10784 8041 10793 8075
rect 10793 8041 10827 8075
rect 10827 8041 10836 8075
rect 10784 8032 10836 8041
rect 10876 8032 10928 8084
rect 14280 8032 14332 8084
rect 1860 7964 1912 8016
rect 2504 7964 2556 8016
rect 2688 7964 2740 8016
rect 3608 7964 3660 8016
rect 4068 7964 4120 8016
rect 2596 7896 2648 7948
rect 4896 7896 4948 7948
rect 6828 7896 6880 7948
rect 1860 7828 1912 7880
rect 6184 7828 6236 7880
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 2136 7760 2188 7812
rect 2412 7760 2464 7812
rect 4068 7760 4120 7812
rect 1768 7692 1820 7744
rect 6552 7760 6604 7812
rect 11060 7964 11112 8016
rect 11704 7964 11756 8016
rect 12072 7964 12124 8016
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 9956 7896 10008 7948
rect 10508 7896 10560 7948
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 11888 7896 11940 7948
rect 12256 7964 12308 8016
rect 15568 8007 15620 8016
rect 15568 7973 15602 8007
rect 15602 7973 15620 8007
rect 15568 7964 15620 7973
rect 17408 8032 17460 8084
rect 17868 8032 17920 8084
rect 18052 8032 18104 8084
rect 19708 8032 19760 8084
rect 20352 7964 20404 8016
rect 10140 7828 10192 7880
rect 11336 7871 11388 7880
rect 11336 7837 11345 7871
rect 11345 7837 11379 7871
rect 11379 7837 11388 7871
rect 13728 7896 13780 7948
rect 15844 7896 15896 7948
rect 16672 7896 16724 7948
rect 17408 7896 17460 7948
rect 17868 7939 17920 7948
rect 17868 7905 17877 7939
rect 17877 7905 17911 7939
rect 17911 7905 17920 7939
rect 17868 7896 17920 7905
rect 18880 7896 18932 7948
rect 20628 7896 20680 7948
rect 12348 7871 12400 7880
rect 11336 7828 11388 7837
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 9864 7760 9916 7812
rect 11704 7760 11756 7812
rect 17776 7828 17828 7880
rect 19892 7871 19944 7880
rect 17500 7760 17552 7812
rect 19892 7837 19901 7871
rect 19901 7837 19935 7871
rect 19935 7837 19944 7871
rect 19892 7828 19944 7837
rect 20444 7760 20496 7812
rect 10876 7692 10928 7744
rect 12256 7692 12308 7744
rect 12624 7692 12676 7744
rect 16764 7692 16816 7744
rect 19892 7692 19944 7744
rect 20812 7692 20864 7744
rect 21272 7692 21324 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 3332 7488 3384 7540
rect 4896 7531 4948 7540
rect 4896 7497 4905 7531
rect 4905 7497 4939 7531
rect 4939 7497 4948 7531
rect 4896 7488 4948 7497
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 6552 7352 6604 7404
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 1768 7327 1820 7336
rect 1768 7293 1777 7327
rect 1777 7293 1811 7327
rect 1811 7293 1820 7327
rect 1768 7284 1820 7293
rect 4896 7284 4948 7336
rect 5264 7284 5316 7336
rect 12624 7488 12676 7540
rect 15292 7488 15344 7540
rect 16856 7488 16908 7540
rect 17224 7488 17276 7540
rect 8484 7420 8536 7472
rect 11244 7420 11296 7472
rect 7840 7352 7892 7404
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 9496 7284 9548 7336
rect 9956 7352 10008 7404
rect 11152 7352 11204 7404
rect 18880 7420 18932 7472
rect 14280 7352 14332 7404
rect 14464 7352 14516 7404
rect 16580 7352 16632 7404
rect 18512 7352 18564 7404
rect 13176 7284 13228 7336
rect 13268 7284 13320 7336
rect 13544 7284 13596 7336
rect 14924 7284 14976 7336
rect 16396 7284 16448 7336
rect 18052 7327 18104 7336
rect 18052 7293 18071 7327
rect 18071 7293 18104 7327
rect 18052 7284 18104 7293
rect 18880 7284 18932 7336
rect 20352 7488 20404 7540
rect 20444 7420 20496 7472
rect 20904 7420 20956 7472
rect 19156 7352 19208 7404
rect 20536 7284 20588 7336
rect 2044 7259 2096 7268
rect 2044 7225 2053 7259
rect 2053 7225 2087 7259
rect 2087 7225 2096 7259
rect 2044 7216 2096 7225
rect 3056 7216 3108 7268
rect 3240 7216 3292 7268
rect 1032 7148 1084 7200
rect 1768 7148 1820 7200
rect 2596 7148 2648 7200
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 3424 7148 3476 7157
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 5356 7191 5408 7200
rect 5356 7157 5365 7191
rect 5365 7157 5399 7191
rect 5399 7157 5408 7191
rect 7196 7191 7248 7200
rect 5356 7148 5408 7157
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 11336 7216 11388 7268
rect 9588 7191 9640 7200
rect 9588 7157 9597 7191
rect 9597 7157 9631 7191
rect 9631 7157 9640 7191
rect 9588 7148 9640 7157
rect 11060 7148 11112 7200
rect 11704 7148 11756 7200
rect 12716 7191 12768 7200
rect 12716 7157 12725 7191
rect 12725 7157 12759 7191
rect 12759 7157 12768 7191
rect 12716 7148 12768 7157
rect 13360 7148 13412 7200
rect 15292 7148 15344 7200
rect 16580 7216 16632 7268
rect 17960 7148 18012 7200
rect 19892 7148 19944 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 5264 6944 5316 6996
rect 7012 6987 7064 6996
rect 7012 6953 7021 6987
rect 7021 6953 7055 6987
rect 7055 6953 7064 6987
rect 7012 6944 7064 6953
rect 5080 6919 5132 6928
rect 5080 6885 5089 6919
rect 5089 6885 5123 6919
rect 5123 6885 5132 6919
rect 5080 6876 5132 6885
rect 6092 6876 6144 6928
rect 8392 6944 8444 6996
rect 9588 6944 9640 6996
rect 11152 6944 11204 6996
rect 12716 6944 12768 6996
rect 16672 6944 16724 6996
rect 17500 6944 17552 6996
rect 1124 6808 1176 6860
rect 1492 6808 1544 6860
rect 2320 6808 2372 6860
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 8208 6876 8260 6928
rect 14280 6876 14332 6928
rect 16764 6876 16816 6928
rect 17224 6876 17276 6928
rect 18880 6876 18932 6928
rect 8392 6808 8444 6860
rect 9036 6808 9088 6860
rect 9772 6808 9824 6860
rect 9956 6851 10008 6860
rect 9956 6817 9990 6851
rect 9990 6817 10008 6851
rect 9956 6808 10008 6817
rect 11244 6808 11296 6860
rect 12348 6808 12400 6860
rect 2780 6740 2832 6792
rect 3424 6740 3476 6792
rect 4712 6740 4764 6792
rect 5632 6740 5684 6792
rect 7380 6672 7432 6724
rect 1216 6604 1268 6656
rect 8208 6604 8260 6656
rect 8760 6740 8812 6792
rect 9312 6740 9364 6792
rect 15844 6808 15896 6860
rect 18512 6808 18564 6860
rect 12716 6672 12768 6724
rect 15200 6672 15252 6724
rect 17592 6715 17644 6724
rect 17592 6681 17601 6715
rect 17601 6681 17635 6715
rect 17635 6681 17644 6715
rect 17592 6672 17644 6681
rect 13544 6604 13596 6656
rect 14280 6604 14332 6656
rect 17868 6672 17920 6724
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 3792 6400 3844 6452
rect 5356 6400 5408 6452
rect 10232 6400 10284 6452
rect 12440 6443 12492 6452
rect 12440 6409 12449 6443
rect 12449 6409 12483 6443
rect 12483 6409 12492 6443
rect 12440 6400 12492 6409
rect 14648 6400 14700 6452
rect 15844 6400 15896 6452
rect 17776 6400 17828 6452
rect 5816 6332 5868 6384
rect 3608 6264 3660 6316
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 1952 6239 2004 6248
rect 1952 6205 1961 6239
rect 1961 6205 1995 6239
rect 1995 6205 2004 6239
rect 1952 6196 2004 6205
rect 2964 6196 3016 6248
rect 4712 6196 4764 6248
rect 8392 6332 8444 6384
rect 9864 6332 9916 6384
rect 7196 6264 7248 6316
rect 7656 6239 7708 6248
rect 7656 6205 7665 6239
rect 7665 6205 7699 6239
rect 7699 6205 7708 6239
rect 7656 6196 7708 6205
rect 8760 6239 8812 6248
rect 8760 6205 8769 6239
rect 8769 6205 8803 6239
rect 8803 6205 8812 6239
rect 8760 6196 8812 6205
rect 12440 6264 12492 6316
rect 12716 6264 12768 6316
rect 15200 6264 15252 6316
rect 17684 6264 17736 6316
rect 18880 6264 18932 6316
rect 10232 6196 10284 6248
rect 10416 6196 10468 6248
rect 10600 6196 10652 6248
rect 11060 6196 11112 6248
rect 5356 6171 5408 6180
rect 5356 6137 5365 6171
rect 5365 6137 5399 6171
rect 5399 6137 5408 6171
rect 5356 6128 5408 6137
rect 5540 6128 5592 6180
rect 5632 6128 5684 6180
rect 9036 6171 9088 6180
rect 3792 6060 3844 6112
rect 8300 6060 8352 6112
rect 8392 6060 8444 6112
rect 8668 6060 8720 6112
rect 9036 6137 9070 6171
rect 9070 6137 9088 6171
rect 9036 6128 9088 6137
rect 9128 6128 9180 6180
rect 13544 6196 13596 6248
rect 15752 6196 15804 6248
rect 16856 6196 16908 6248
rect 18788 6239 18840 6248
rect 18788 6205 18797 6239
rect 18797 6205 18831 6239
rect 18831 6205 18840 6239
rect 18788 6196 18840 6205
rect 19892 6196 19944 6248
rect 20076 6196 20128 6248
rect 20536 6264 20588 6316
rect 15936 6128 15988 6180
rect 17408 6128 17460 6180
rect 17500 6128 17552 6180
rect 18880 6171 18932 6180
rect 18880 6137 18889 6171
rect 18889 6137 18923 6171
rect 18923 6137 18932 6171
rect 18880 6128 18932 6137
rect 9864 6060 9916 6112
rect 9956 6060 10008 6112
rect 10416 6060 10468 6112
rect 11060 6060 11112 6112
rect 13820 6060 13872 6112
rect 16764 6103 16816 6112
rect 16764 6069 16773 6103
rect 16773 6069 16807 6103
rect 16807 6069 16816 6103
rect 16764 6060 16816 6069
rect 16856 6103 16908 6112
rect 16856 6069 16865 6103
rect 16865 6069 16899 6103
rect 16899 6069 16908 6103
rect 16856 6060 16908 6069
rect 18788 6060 18840 6112
rect 19156 6060 19208 6112
rect 20076 6103 20128 6112
rect 20076 6069 20085 6103
rect 20085 6069 20119 6103
rect 20119 6069 20128 6103
rect 20076 6060 20128 6069
rect 20536 6103 20588 6112
rect 20536 6069 20545 6103
rect 20545 6069 20579 6103
rect 20579 6069 20588 6103
rect 20536 6060 20588 6069
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 2872 5856 2924 5908
rect 3516 5856 3568 5908
rect 4344 5856 4396 5908
rect 5172 5856 5224 5908
rect 6460 5899 6512 5908
rect 6460 5865 6469 5899
rect 6469 5865 6503 5899
rect 6503 5865 6512 5899
rect 6460 5856 6512 5865
rect 2044 5720 2096 5772
rect 4712 5720 4764 5772
rect 7196 5788 7248 5840
rect 6368 5720 6420 5772
rect 8668 5856 8720 5908
rect 10692 5856 10744 5908
rect 12716 5899 12768 5908
rect 3700 5652 3752 5704
rect 9312 5788 9364 5840
rect 8484 5763 8536 5772
rect 8484 5729 8493 5763
rect 8493 5729 8527 5763
rect 8527 5729 8536 5763
rect 8484 5720 8536 5729
rect 8668 5720 8720 5772
rect 9128 5720 9180 5772
rect 11152 5788 11204 5840
rect 11520 5788 11572 5840
rect 12716 5865 12725 5899
rect 12725 5865 12759 5899
rect 12759 5865 12768 5899
rect 12716 5856 12768 5865
rect 13544 5899 13596 5908
rect 13544 5865 13553 5899
rect 13553 5865 13587 5899
rect 13587 5865 13596 5899
rect 13544 5856 13596 5865
rect 14648 5856 14700 5908
rect 15292 5899 15344 5908
rect 15292 5865 15301 5899
rect 15301 5865 15335 5899
rect 15335 5865 15344 5899
rect 15292 5856 15344 5865
rect 16764 5856 16816 5908
rect 19248 5856 19300 5908
rect 19156 5788 19208 5840
rect 6092 5584 6144 5636
rect 9312 5652 9364 5704
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10416 5695 10468 5704
rect 10232 5652 10284 5661
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 11336 5695 11388 5704
rect 11336 5661 11345 5695
rect 11345 5661 11379 5695
rect 11379 5661 11388 5695
rect 11336 5652 11388 5661
rect 6644 5516 6696 5568
rect 8024 5516 8076 5568
rect 8668 5559 8720 5568
rect 8668 5525 8677 5559
rect 8677 5525 8711 5559
rect 8711 5525 8720 5559
rect 8668 5516 8720 5525
rect 9128 5516 9180 5568
rect 9864 5516 9916 5568
rect 11152 5584 11204 5636
rect 12624 5720 12676 5772
rect 15660 5763 15712 5772
rect 15660 5729 15669 5763
rect 15669 5729 15703 5763
rect 15703 5729 15712 5763
rect 15660 5720 15712 5729
rect 17776 5720 17828 5772
rect 17960 5720 18012 5772
rect 14372 5652 14424 5704
rect 15200 5652 15252 5704
rect 17592 5652 17644 5704
rect 18880 5652 18932 5704
rect 10784 5516 10836 5568
rect 13544 5516 13596 5568
rect 18972 5516 19024 5568
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 1584 5312 1636 5364
rect 3148 5312 3200 5364
rect 4160 5355 4212 5364
rect 4160 5321 4169 5355
rect 4169 5321 4203 5355
rect 4203 5321 4212 5355
rect 4160 5312 4212 5321
rect 5448 5312 5500 5364
rect 7564 5312 7616 5364
rect 8208 5355 8260 5364
rect 8208 5321 8217 5355
rect 8217 5321 8251 5355
rect 8251 5321 8260 5355
rect 8208 5312 8260 5321
rect 9496 5312 9548 5364
rect 11060 5312 11112 5364
rect 11704 5312 11756 5364
rect 14188 5312 14240 5364
rect 16856 5312 16908 5364
rect 17960 5312 18012 5364
rect 20260 5312 20312 5364
rect 9312 5244 9364 5296
rect 10324 5244 10376 5296
rect 7104 5176 7156 5228
rect 8576 5176 8628 5228
rect 9036 5176 9088 5228
rect 10692 5176 10744 5228
rect 11336 5219 11388 5228
rect 11336 5185 11345 5219
rect 11345 5185 11379 5219
rect 11379 5185 11388 5219
rect 11336 5176 11388 5185
rect 11704 5176 11756 5228
rect 14372 5176 14424 5228
rect 16672 5176 16724 5228
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 4160 5108 4212 5160
rect 4988 5108 5040 5160
rect 8024 5151 8076 5160
rect 8024 5117 8033 5151
rect 8033 5117 8067 5151
rect 8067 5117 8076 5151
rect 8024 5108 8076 5117
rect 12624 5108 12676 5160
rect 13176 5108 13228 5160
rect 14004 5108 14056 5160
rect 17224 5244 17276 5296
rect 17592 5176 17644 5228
rect 18880 5244 18932 5296
rect 20352 5244 20404 5296
rect 20076 5176 20128 5228
rect 9312 5040 9364 5092
rect 9772 5040 9824 5092
rect 8208 4972 8260 5024
rect 12440 5040 12492 5092
rect 11060 4972 11112 5024
rect 12348 4972 12400 5024
rect 14188 4972 14240 5024
rect 14280 4972 14332 5024
rect 16856 5015 16908 5024
rect 16856 4981 16865 5015
rect 16865 4981 16899 5015
rect 16899 4981 16908 5015
rect 16856 4972 16908 4981
rect 17132 4972 17184 5024
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 1676 4768 1728 4820
rect 4804 4768 4856 4820
rect 6000 4768 6052 4820
rect 7748 4768 7800 4820
rect 8392 4768 8444 4820
rect 10324 4768 10376 4820
rect 11060 4811 11112 4820
rect 11060 4777 11069 4811
rect 11069 4777 11103 4811
rect 11103 4777 11112 4811
rect 11060 4768 11112 4777
rect 11520 4811 11572 4820
rect 11520 4777 11529 4811
rect 11529 4777 11563 4811
rect 11563 4777 11572 4811
rect 11520 4768 11572 4777
rect 3976 4700 4028 4752
rect 12348 4768 12400 4820
rect 13452 4768 13504 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 14648 4768 14700 4820
rect 15476 4811 15528 4820
rect 15476 4777 15485 4811
rect 15485 4777 15519 4811
rect 15519 4777 15528 4811
rect 15476 4768 15528 4777
rect 16856 4768 16908 4820
rect 18788 4768 18840 4820
rect 19340 4768 19392 4820
rect 1860 4632 1912 4684
rect 3332 4632 3384 4684
rect 4252 4632 4304 4684
rect 13360 4700 13412 4752
rect 14188 4700 14240 4752
rect 16672 4700 16724 4752
rect 3976 4564 4028 4616
rect 9404 4632 9456 4684
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 11060 4632 11112 4684
rect 11520 4564 11572 4616
rect 11704 4607 11756 4616
rect 11704 4573 11713 4607
rect 11713 4573 11747 4607
rect 11747 4573 11756 4607
rect 11704 4564 11756 4573
rect 20 4496 72 4548
rect 14556 4564 14608 4616
rect 15384 4632 15436 4684
rect 16396 4632 16448 4684
rect 17684 4700 17736 4752
rect 18144 4700 18196 4752
rect 16856 4675 16908 4684
rect 16856 4641 16865 4675
rect 16865 4641 16899 4675
rect 16899 4641 16908 4675
rect 16856 4632 16908 4641
rect 17500 4632 17552 4684
rect 17592 4632 17644 4684
rect 17224 4564 17276 4616
rect 19524 4700 19576 4752
rect 20260 4700 20312 4752
rect 19432 4632 19484 4684
rect 19524 4564 19576 4616
rect 20720 4564 20772 4616
rect 12440 4496 12492 4548
rect 18788 4496 18840 4548
rect 3792 4428 3844 4480
rect 9036 4428 9088 4480
rect 9588 4428 9640 4480
rect 14280 4428 14332 4480
rect 17132 4428 17184 4480
rect 19616 4428 19668 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 1492 4088 1544 4140
rect 4804 4088 4856 4140
rect 5080 4131 5132 4140
rect 5080 4097 5089 4131
rect 5089 4097 5123 4131
rect 5123 4097 5132 4131
rect 5080 4088 5132 4097
rect 10048 4224 10100 4276
rect 10324 4267 10376 4276
rect 10324 4233 10333 4267
rect 10333 4233 10367 4267
rect 10367 4233 10376 4267
rect 10324 4224 10376 4233
rect 12348 4224 12400 4276
rect 15200 4224 15252 4276
rect 16856 4224 16908 4276
rect 17132 4224 17184 4276
rect 17500 4224 17552 4276
rect 21364 4224 21416 4276
rect 9864 4156 9916 4208
rect 14280 4156 14332 4208
rect 14556 4156 14608 4208
rect 2780 4020 2832 4072
rect 3884 4020 3936 4072
rect 12348 4088 12400 4140
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 13728 4088 13780 4140
rect 16304 4156 16356 4208
rect 17040 4156 17092 4208
rect 17408 4088 17460 4140
rect 18788 4088 18840 4140
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 10784 4020 10836 4072
rect 12256 4020 12308 4072
rect 14740 4020 14792 4072
rect 16120 4020 16172 4072
rect 16304 4020 16356 4072
rect 19340 4020 19392 4072
rect 20444 4020 20496 4072
rect 10048 3952 10100 4004
rect 1400 3884 1452 3936
rect 3056 3927 3108 3936
rect 3056 3893 3065 3927
rect 3065 3893 3099 3927
rect 3099 3893 3108 3927
rect 3056 3884 3108 3893
rect 4160 3927 4212 3936
rect 4160 3893 4169 3927
rect 4169 3893 4203 3927
rect 4203 3893 4212 3927
rect 4160 3884 4212 3893
rect 8208 3884 8260 3936
rect 8944 3884 8996 3936
rect 9680 3884 9732 3936
rect 10508 3952 10560 4004
rect 17500 3952 17552 4004
rect 17868 3952 17920 4004
rect 12440 3884 12492 3936
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 12900 3884 12952 3893
rect 13912 3884 13964 3936
rect 15568 3884 15620 3936
rect 16028 3884 16080 3936
rect 16396 3884 16448 3936
rect 16764 3884 16816 3936
rect 19064 3884 19116 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 2136 3680 2188 3732
rect 4896 3680 4948 3732
rect 5908 3680 5960 3732
rect 9680 3680 9732 3732
rect 10048 3723 10100 3732
rect 10048 3689 10057 3723
rect 10057 3689 10091 3723
rect 10091 3689 10100 3723
rect 10048 3680 10100 3689
rect 11980 3680 12032 3732
rect 12164 3680 12216 3732
rect 12440 3723 12492 3732
rect 12440 3689 12449 3723
rect 12449 3689 12483 3723
rect 12483 3689 12492 3723
rect 12440 3680 12492 3689
rect 12900 3680 12952 3732
rect 14004 3723 14056 3732
rect 14004 3689 14013 3723
rect 14013 3689 14047 3723
rect 14047 3689 14056 3723
rect 14004 3680 14056 3689
rect 16764 3680 16816 3732
rect 16856 3680 16908 3732
rect 17776 3680 17828 3732
rect 18144 3680 18196 3732
rect 19616 3723 19668 3732
rect 19616 3689 19625 3723
rect 19625 3689 19659 3723
rect 19659 3689 19668 3723
rect 19616 3680 19668 3689
rect 8668 3612 8720 3664
rect 2228 3544 2280 3596
rect 4068 3587 4120 3596
rect 4068 3553 4077 3587
rect 4077 3553 4111 3587
rect 4111 3553 4120 3587
rect 4068 3544 4120 3553
rect 10876 3612 10928 3664
rect 12624 3612 12676 3664
rect 13820 3612 13872 3664
rect 14372 3612 14424 3664
rect 16120 3612 16172 3664
rect 9864 3587 9916 3596
rect 9864 3553 9873 3587
rect 9873 3553 9907 3587
rect 9907 3553 9916 3587
rect 9864 3544 9916 3553
rect 10692 3544 10744 3596
rect 13728 3544 13780 3596
rect 14648 3544 14700 3596
rect 17316 3612 17368 3664
rect 10600 3476 10652 3528
rect 12808 3476 12860 3528
rect 14188 3519 14240 3528
rect 14188 3485 14197 3519
rect 14197 3485 14231 3519
rect 14231 3485 14240 3519
rect 16488 3519 16540 3528
rect 14188 3476 14240 3485
rect 16488 3485 16497 3519
rect 16497 3485 16531 3519
rect 16531 3485 16540 3519
rect 16488 3476 16540 3485
rect 18052 3544 18104 3596
rect 19156 3612 19208 3664
rect 18328 3544 18380 3596
rect 19984 3544 20036 3596
rect 18880 3476 18932 3528
rect 19340 3476 19392 3528
rect 20260 3476 20312 3528
rect 4252 3451 4304 3460
rect 4252 3417 4261 3451
rect 4261 3417 4295 3451
rect 4295 3417 4304 3451
rect 4252 3408 4304 3417
rect 3976 3340 4028 3392
rect 5632 3408 5684 3460
rect 5816 3408 5868 3460
rect 17500 3408 17552 3460
rect 4804 3340 4856 3392
rect 11980 3340 12032 3392
rect 12440 3340 12492 3392
rect 20720 3408 20772 3460
rect 19156 3383 19208 3392
rect 19156 3349 19165 3383
rect 19165 3349 19199 3383
rect 19199 3349 19208 3383
rect 19156 3340 19208 3349
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 1308 3136 1360 3188
rect 2504 3136 2556 3188
rect 5816 3136 5868 3188
rect 8576 3111 8628 3120
rect 8576 3077 8585 3111
rect 8585 3077 8619 3111
rect 8619 3077 8628 3111
rect 8576 3068 8628 3077
rect 10968 3136 11020 3188
rect 11796 3136 11848 3188
rect 11980 3136 12032 3188
rect 16304 3136 16356 3188
rect 16488 3136 16540 3188
rect 16672 3136 16724 3188
rect 20168 3136 20220 3188
rect 12440 3068 12492 3120
rect 12624 3068 12676 3120
rect 9312 3000 9364 3052
rect 14556 3043 14608 3052
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 14648 3043 14700 3052
rect 14648 3009 14657 3043
rect 14657 3009 14691 3043
rect 14691 3009 14700 3043
rect 17040 3043 17092 3052
rect 14648 3000 14700 3009
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 2872 2975 2924 2984
rect 2872 2941 2881 2975
rect 2881 2941 2915 2975
rect 2915 2941 2924 2975
rect 2872 2932 2924 2941
rect 8760 2932 8812 2984
rect 10140 2975 10192 2984
rect 10140 2941 10149 2975
rect 10149 2941 10183 2975
rect 10183 2941 10192 2975
rect 10140 2932 10192 2941
rect 11244 2975 11296 2984
rect 11244 2941 11253 2975
rect 11253 2941 11287 2975
rect 11287 2941 11296 2975
rect 11244 2932 11296 2941
rect 12716 2932 12768 2984
rect 14280 2932 14332 2984
rect 15476 2932 15528 2984
rect 16764 2975 16816 2984
rect 16764 2941 16773 2975
rect 16773 2941 16807 2975
rect 16807 2941 16816 2975
rect 16764 2932 16816 2941
rect 19156 2932 19208 2984
rect 19708 2932 19760 2984
rect 7104 2864 7156 2916
rect 7564 2864 7616 2916
rect 10508 2864 10560 2916
rect 10600 2864 10652 2916
rect 14188 2864 14240 2916
rect 16948 2864 17000 2916
rect 19064 2864 19116 2916
rect 3056 2839 3108 2848
rect 3056 2805 3065 2839
rect 3065 2805 3099 2839
rect 3099 2805 3108 2839
rect 3056 2796 3108 2805
rect 7288 2796 7340 2848
rect 11244 2796 11296 2848
rect 16580 2796 16632 2848
rect 19248 2796 19300 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 4068 2592 4120 2644
rect 5356 2592 5408 2644
rect 9128 2592 9180 2644
rect 11060 2592 11112 2644
rect 13268 2592 13320 2644
rect 13820 2635 13872 2644
rect 13820 2601 13829 2635
rect 13829 2601 13863 2635
rect 13863 2601 13872 2635
rect 13820 2592 13872 2601
rect 14188 2635 14240 2644
rect 14188 2601 14197 2635
rect 14197 2601 14231 2635
rect 14231 2601 14240 2635
rect 14188 2592 14240 2601
rect 16396 2592 16448 2644
rect 17132 2592 17184 2644
rect 19800 2592 19852 2644
rect 13544 2524 13596 2576
rect 1860 2499 1912 2508
rect 1860 2465 1869 2499
rect 1869 2465 1903 2499
rect 1903 2465 1912 2499
rect 1860 2456 1912 2465
rect 17868 2524 17920 2576
rect 2780 2388 2832 2440
rect 5448 2388 5500 2440
rect 18052 2456 18104 2508
rect 19432 2499 19484 2508
rect 19432 2465 19441 2499
rect 19441 2465 19475 2499
rect 19475 2465 19484 2499
rect 19432 2456 19484 2465
rect 13728 2320 13780 2372
rect 2044 2295 2096 2304
rect 2044 2261 2053 2295
rect 2053 2261 2087 2295
rect 2087 2261 2096 2295
rect 2044 2252 2096 2261
rect 6920 2252 6972 2304
rect 13452 2252 13504 2304
rect 14280 2431 14332 2440
rect 14280 2397 14289 2431
rect 14289 2397 14323 2431
rect 14323 2397 14332 2431
rect 14280 2388 14332 2397
rect 14648 2388 14700 2440
rect 17316 2388 17368 2440
rect 16212 2320 16264 2372
rect 18696 2252 18748 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 2044 2048 2096 2100
rect 7472 1980 7524 2032
rect 14280 1980 14332 2032
rect 14372 1980 14424 2032
rect 18512 1980 18564 2032
rect 14004 1844 14056 1896
rect 18696 1844 18748 1896
rect 13728 1776 13780 1828
rect 19524 1776 19576 1828
rect 8852 1708 8904 1760
rect 18052 1708 18104 1760
rect 21456 1640 21508 1692
rect 10508 1572 10560 1624
rect 16120 1572 16172 1624
rect 13084 1300 13136 1352
rect 18144 1300 18196 1352
rect 2320 1232 2372 1284
rect 5908 1232 5960 1284
<< metal2 >>
rect 202 22520 258 23000
rect 662 22520 718 23000
rect 1122 22520 1178 23000
rect 1582 22520 1638 23000
rect 2042 22520 2098 23000
rect 2502 22520 2558 23000
rect 2962 22520 3018 23000
rect 3422 22520 3478 23000
rect 3698 22672 3754 22681
rect 3698 22607 3754 22616
rect 18 18864 74 18873
rect 18 18799 74 18808
rect 32 4554 60 18799
rect 216 18086 244 22520
rect 204 18080 256 18086
rect 204 18022 256 18028
rect 676 11937 704 22520
rect 1136 13297 1164 22520
rect 1398 19000 1454 19009
rect 1398 18935 1400 18944
rect 1452 18935 1454 18944
rect 1400 18906 1452 18912
rect 1596 18902 1624 22520
rect 1950 20632 2006 20641
rect 1950 20567 2006 20576
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 1768 19168 1820 19174
rect 1768 19110 1820 19116
rect 1584 18896 1636 18902
rect 1584 18838 1636 18844
rect 1398 18592 1454 18601
rect 1398 18527 1454 18536
rect 1308 18080 1360 18086
rect 1308 18022 1360 18028
rect 1214 16960 1270 16969
rect 1214 16895 1270 16904
rect 1122 13288 1178 13297
rect 1122 13223 1178 13232
rect 662 11928 718 11937
rect 662 11863 718 11872
rect 1228 11665 1256 16895
rect 1214 11656 1270 11665
rect 1214 11591 1270 11600
rect 1124 10804 1176 10810
rect 1124 10746 1176 10752
rect 1030 10704 1086 10713
rect 1030 10639 1086 10648
rect 570 10160 626 10169
rect 570 10095 626 10104
rect 584 9994 612 10095
rect 572 9988 624 9994
rect 572 9930 624 9936
rect 1044 7206 1072 10639
rect 1032 7200 1084 7206
rect 1032 7142 1084 7148
rect 1136 6866 1164 10746
rect 1216 9648 1268 9654
rect 1216 9590 1268 9596
rect 1124 6860 1176 6866
rect 1124 6802 1176 6808
rect 1228 6662 1256 9590
rect 1216 6656 1268 6662
rect 1216 6598 1268 6604
rect 20 4548 72 4554
rect 20 4490 72 4496
rect 1320 3194 1348 18022
rect 1412 3942 1440 18527
rect 1780 18222 1808 19110
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1766 17096 1822 17105
rect 1766 17031 1822 17040
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1504 10810 1532 16594
rect 1674 16144 1730 16153
rect 1674 16079 1730 16088
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1596 10690 1624 15846
rect 1504 10662 1624 10690
rect 1504 9654 1532 10662
rect 1688 10554 1716 16079
rect 1596 10526 1716 10554
rect 1492 9648 1544 9654
rect 1492 9590 1544 9596
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1504 9178 1532 9454
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1504 4146 1532 6802
rect 1596 5370 1624 10526
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10266 1716 10406
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1780 10010 1808 17031
rect 1872 16522 1900 19790
rect 1964 16538 1992 20567
rect 2056 17241 2084 22520
rect 2228 20256 2280 20262
rect 2228 20198 2280 20204
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2042 17232 2098 17241
rect 2042 17167 2098 17176
rect 1860 16516 1912 16522
rect 1964 16510 2084 16538
rect 1860 16458 1912 16464
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1872 12481 1900 12650
rect 1858 12472 1914 12481
rect 1858 12407 1914 12416
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1688 9982 1808 10010
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1688 4826 1716 9982
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1780 8430 1808 9862
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1872 8022 1900 11086
rect 1860 8016 1912 8022
rect 1860 7958 1912 7964
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1780 7342 1808 7686
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1780 4570 1808 7142
rect 1872 4690 1900 7822
rect 1964 6254 1992 15302
rect 2056 7392 2084 16510
rect 2148 7818 2176 19110
rect 2240 18290 2268 20198
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 2516 17762 2544 22520
rect 2976 21298 3004 22520
rect 2976 21270 3188 21298
rect 2962 21176 3018 21185
rect 2962 21111 3018 21120
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2700 19378 2728 20402
rect 2780 20256 2832 20262
rect 2780 20198 2832 20204
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 2332 17734 2544 17762
rect 2332 15910 2360 17734
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2424 17134 2452 17614
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2516 16794 2544 17614
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2320 14816 2372 14822
rect 2320 14758 2372 14764
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2240 12481 2268 13806
rect 2226 12472 2282 12481
rect 2226 12407 2282 12416
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2240 11898 2268 12242
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2226 11792 2282 11801
rect 2226 11727 2282 11736
rect 2240 9489 2268 11727
rect 2226 9480 2282 9489
rect 2226 9415 2282 9424
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 2056 7364 2176 7392
rect 2044 7268 2096 7274
rect 2044 7210 2096 7216
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 2056 5778 2084 7210
rect 2044 5772 2096 5778
rect 2044 5714 2096 5720
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 1780 4542 1900 4570
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 1308 3188 1360 3194
rect 1308 3130 1360 3136
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1780 2825 1808 2926
rect 1766 2816 1822 2825
rect 1766 2751 1822 2760
rect 1872 2514 1900 4542
rect 2148 3738 2176 7364
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 2240 3602 2268 9415
rect 2332 6866 2360 14758
rect 2504 14340 2556 14346
rect 2504 14282 2556 14288
rect 2516 13802 2544 14282
rect 2504 13796 2556 13802
rect 2504 13738 2556 13744
rect 2608 13546 2636 18566
rect 2700 16561 2728 19110
rect 2792 18698 2820 20198
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2884 16810 2912 19654
rect 2792 16782 2912 16810
rect 2686 16552 2742 16561
rect 2686 16487 2742 16496
rect 2792 15722 2820 16782
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 2700 15694 2820 15722
rect 2700 15042 2728 15694
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2792 15162 2820 15506
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 2700 15014 2820 15042
rect 2792 14482 2820 15014
rect 2884 14618 2912 16662
rect 2976 15065 3004 21111
rect 3056 20460 3108 20466
rect 3056 20402 3108 20408
rect 3068 19854 3096 20402
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 3068 19242 3096 19790
rect 3056 19236 3108 19242
rect 3056 19178 3108 19184
rect 3160 19174 3188 21270
rect 3436 19394 3464 22520
rect 3514 22128 3570 22137
rect 3514 22063 3570 22072
rect 3528 21690 3556 22063
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 3514 21584 3570 21593
rect 3514 21519 3570 21528
rect 3528 20806 3556 21519
rect 3712 20874 3740 22607
rect 3882 22520 3938 23000
rect 4342 22520 4398 23000
rect 4802 22520 4858 23000
rect 5262 22520 5318 23000
rect 5722 22520 5778 23000
rect 6182 22520 6238 23000
rect 6642 22520 6698 23000
rect 7102 22520 7158 23000
rect 7562 22520 7618 23000
rect 8022 22520 8078 23000
rect 8482 22520 8538 23000
rect 8942 22520 8998 23000
rect 9402 22520 9458 23000
rect 9862 22520 9918 23000
rect 10322 22520 10378 23000
rect 10782 22520 10838 23000
rect 11242 22520 11298 23000
rect 11702 22520 11758 23000
rect 12162 22520 12218 23000
rect 12622 22520 12678 23000
rect 13082 22520 13138 23000
rect 13542 22520 13598 23000
rect 14002 22520 14058 23000
rect 14462 22520 14518 23000
rect 14922 22520 14978 23000
rect 15382 22520 15438 23000
rect 15842 22520 15898 23000
rect 16302 22520 16358 23000
rect 16762 22520 16818 23000
rect 17222 22520 17278 23000
rect 17682 22520 17738 23000
rect 17866 22672 17922 22681
rect 17866 22607 17922 22616
rect 3700 20868 3752 20874
rect 3700 20810 3752 20816
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3896 20346 3924 22520
rect 3804 20318 3924 20346
rect 3976 20324 4028 20330
rect 3332 19372 3384 19378
rect 3436 19366 3556 19394
rect 3332 19314 3384 19320
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 3344 18290 3372 19314
rect 3528 18329 3556 19366
rect 3700 19236 3752 19242
rect 3700 19178 3752 19184
rect 3514 18320 3570 18329
rect 3332 18284 3384 18290
rect 3514 18255 3570 18264
rect 3332 18226 3384 18232
rect 3146 18184 3202 18193
rect 3056 18148 3108 18154
rect 3146 18119 3202 18128
rect 3056 18090 3108 18096
rect 3068 17678 3096 18090
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 3056 17060 3108 17066
rect 3056 17002 3108 17008
rect 3068 16250 3096 17002
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 3068 15502 3096 16186
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2962 15056 3018 15065
rect 2962 14991 3018 15000
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2884 14498 2912 14554
rect 2780 14476 2832 14482
rect 2884 14470 3004 14498
rect 2780 14418 2832 14424
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2516 13518 2636 13546
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2516 12730 2544 13518
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2608 12850 2636 13398
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2424 11150 2452 12718
rect 2516 12702 2636 12730
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2516 11762 2544 12582
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2424 10606 2452 10950
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2516 9654 2544 10610
rect 2504 9648 2556 9654
rect 2504 9590 2556 9596
rect 2516 9042 2544 9590
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2504 8016 2556 8022
rect 2504 7958 2556 7964
rect 2412 7812 2464 7818
rect 2412 7754 2464 7760
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2424 6361 2452 7754
rect 2410 6352 2466 6361
rect 2410 6287 2466 6296
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2516 3194 2544 7958
rect 2608 7954 2636 12702
rect 2700 10742 2728 14350
rect 2688 10736 2740 10742
rect 2688 10678 2740 10684
rect 2792 10198 2820 14418
rect 2872 13796 2924 13802
rect 2872 13738 2924 13744
rect 2884 13190 2912 13738
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2884 12238 2912 13126
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2976 11744 3004 14470
rect 3160 13394 3188 18119
rect 3344 17678 3372 18226
rect 3332 17672 3384 17678
rect 3238 17640 3294 17649
rect 3332 17614 3384 17620
rect 3238 17575 3294 17584
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 3068 12646 3096 13330
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3068 12458 3096 12582
rect 3068 12430 3179 12458
rect 3151 12424 3179 12430
rect 3151 12396 3188 12424
rect 3054 12336 3110 12345
rect 3054 12271 3110 12280
rect 2884 11716 3004 11744
rect 2780 10192 2832 10198
rect 2884 10169 2912 11716
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2780 10134 2832 10140
rect 2870 10160 2926 10169
rect 2870 10095 2926 10104
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2700 9450 2728 9658
rect 2792 9489 2820 9862
rect 2778 9480 2834 9489
rect 2688 9444 2740 9450
rect 2778 9415 2834 9424
rect 2688 9386 2740 9392
rect 2700 8022 2728 9386
rect 2884 9178 2912 9998
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2596 7948 2648 7954
rect 2596 7890 2648 7896
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 2056 2106 2084 2246
rect 2044 2100 2096 2106
rect 2044 2042 2096 2048
rect 2320 1284 2372 1290
rect 2320 1226 2372 1232
rect 2332 480 2360 1226
rect 2608 1193 2636 7142
rect 2792 6882 2820 8910
rect 2884 8362 2912 9114
rect 2976 8974 3004 11562
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2976 8634 3004 8774
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2792 6854 2912 6882
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2792 4078 2820 6734
rect 2884 5914 2912 6854
rect 2976 6254 3004 8434
rect 3068 7274 3096 12271
rect 3160 11762 3188 12396
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10674 3188 11086
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3252 10554 3280 17575
rect 3344 17338 3372 17614
rect 3712 17338 3740 19178
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3344 16046 3372 17274
rect 3606 16688 3662 16697
rect 3606 16623 3662 16632
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3344 15570 3372 15982
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3344 13870 3372 15506
rect 3514 14648 3570 14657
rect 3514 14583 3570 14592
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3436 13870 3464 14350
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3344 13462 3372 13806
rect 3332 13456 3384 13462
rect 3332 13398 3384 13404
rect 3344 12306 3372 13398
rect 3436 12374 3464 13806
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3424 12164 3476 12170
rect 3424 12106 3476 12112
rect 3436 11506 3464 12106
rect 3528 11665 3556 14583
rect 3514 11656 3570 11665
rect 3514 11591 3570 11600
rect 3436 11478 3556 11506
rect 3160 10526 3280 10554
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 3054 5672 3110 5681
rect 3054 5607 3110 5616
rect 2870 5264 2926 5273
rect 2870 5199 2926 5208
rect 2884 5166 2912 5199
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2870 4720 2926 4729
rect 2870 4655 2926 4664
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2884 2990 2912 4655
rect 3068 3942 3096 5607
rect 3160 5370 3188 10526
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3252 9518 3280 10406
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 7426 3280 9318
rect 3344 7546 3372 10542
rect 3424 10192 3476 10198
rect 3424 10134 3476 10140
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3252 7398 3372 7426
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 3054 2952 3110 2961
rect 3054 2887 3110 2896
rect 3068 2854 3096 2887
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2792 2145 2820 2382
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect 2594 1184 2650 1193
rect 2594 1119 2650 1128
rect 2318 0 2374 480
rect 3252 241 3280 7210
rect 3344 4690 3372 7398
rect 3436 7206 3464 10134
rect 3528 8634 3556 11478
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3620 8242 3648 16623
rect 3712 16590 3740 17274
rect 3804 17270 3832 20318
rect 3976 20266 4028 20272
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3896 17814 3924 20198
rect 3988 20097 4016 20266
rect 3974 20088 4030 20097
rect 3974 20023 4030 20032
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4172 18970 4200 19994
rect 4356 19802 4384 22520
rect 4816 20942 4844 22520
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4712 20256 4764 20262
rect 4712 20198 4764 20204
rect 4724 20058 4752 20198
rect 4908 20074 4936 20742
rect 4988 20324 5040 20330
rect 4988 20266 5040 20272
rect 5000 20210 5028 20266
rect 5000 20182 5120 20210
rect 4712 20052 4764 20058
rect 4908 20046 5028 20074
rect 4712 19994 4764 20000
rect 4896 19848 4948 19854
rect 4356 19774 4844 19802
rect 4896 19790 4948 19796
rect 4250 19680 4306 19689
rect 4250 19615 4306 19624
rect 4264 19258 4292 19615
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4264 19230 4384 19258
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 4080 18737 4108 18906
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 4066 18728 4122 18737
rect 4066 18663 4122 18672
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 3884 17808 3936 17814
rect 3884 17750 3936 17756
rect 3792 17264 3844 17270
rect 3792 17206 3844 17212
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3712 14618 3740 14758
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 3804 14482 3832 16458
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3896 15366 3924 15914
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3896 15026 3924 15302
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3700 14340 3752 14346
rect 3700 14282 3752 14288
rect 3712 12345 3740 14282
rect 3988 14113 4016 18158
rect 4172 17882 4200 18770
rect 4264 18154 4292 19110
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4160 17876 4212 17882
rect 4356 17864 4384 19230
rect 4816 18873 4844 19774
rect 4908 19174 4936 19790
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 5000 18986 5028 20046
rect 4908 18958 5028 18986
rect 4802 18864 4858 18873
rect 4802 18799 4858 18808
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4816 18426 4844 18702
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4160 17818 4212 17824
rect 4264 17836 4384 17864
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4080 15978 4108 16594
rect 4068 15972 4120 15978
rect 4068 15914 4120 15920
rect 4066 15600 4122 15609
rect 4172 15586 4200 16730
rect 4122 15558 4200 15586
rect 4066 15535 4122 15544
rect 4066 15192 4122 15201
rect 4066 15127 4122 15136
rect 3974 14104 4030 14113
rect 3974 14039 4030 14048
rect 4080 13870 4108 15127
rect 4264 14056 4292 17836
rect 4816 17814 4844 18362
rect 4804 17808 4856 17814
rect 4804 17750 4856 17756
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4356 17338 4384 17682
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4632 15706 4660 15846
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4172 14028 4292 14056
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 3974 13696 4030 13705
rect 3974 13631 4030 13640
rect 3790 13152 3846 13161
rect 3790 13087 3846 13096
rect 3698 12336 3754 12345
rect 3698 12271 3754 12280
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 3712 11558 3740 12106
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3712 10713 3740 11494
rect 3698 10704 3754 10713
rect 3698 10639 3754 10648
rect 3700 10600 3752 10606
rect 3698 10568 3700 10577
rect 3752 10568 3754 10577
rect 3698 10503 3754 10512
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3712 10305 3740 10406
rect 3698 10296 3754 10305
rect 3698 10231 3754 10240
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3712 9722 3740 10066
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3698 9616 3754 9625
rect 3698 9551 3754 9560
rect 3528 8214 3648 8242
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3436 2689 3464 6734
rect 3528 5914 3556 8214
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3620 7410 3648 7958
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3712 7290 3740 9551
rect 3620 7262 3740 7290
rect 3620 6322 3648 7262
rect 3804 6458 3832 13087
rect 3882 12608 3938 12617
rect 3882 12543 3938 12552
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3422 2680 3478 2689
rect 3422 2615 3478 2624
rect 3620 649 3648 6258
rect 3790 6216 3846 6225
rect 3790 6151 3846 6160
rect 3804 6118 3832 6151
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3712 3233 3740 5646
rect 3790 5128 3846 5137
rect 3790 5063 3846 5072
rect 3804 4486 3832 5063
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3896 4078 3924 12543
rect 3988 11626 4016 13631
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 4080 12442 4108 13126
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3976 11620 4028 11626
rect 3976 11562 4028 11568
rect 4080 11218 4108 12038
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3988 10266 4016 10610
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3988 9654 4016 10202
rect 4080 9722 4108 10678
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 3974 9480 4030 9489
rect 3974 9415 4030 9424
rect 3988 9042 4016 9415
rect 4066 9344 4122 9353
rect 4066 9279 4122 9288
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3974 8664 4030 8673
rect 3974 8599 4030 8608
rect 3988 4758 4016 8599
rect 4080 8362 4108 9279
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 4080 8022 4108 8055
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 4080 7177 4108 7754
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 4066 6624 4122 6633
rect 4066 6559 4122 6568
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3988 4185 4016 4558
rect 3974 4176 4030 4185
rect 3974 4111 4030 4120
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3974 3632 4030 3641
rect 4080 3602 4108 6559
rect 4172 5370 4200 14028
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4264 11762 4292 12718
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4250 11656 4306 11665
rect 4250 11591 4306 11600
rect 4264 9178 4292 11591
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4160 5160 4212 5166
rect 4158 5128 4160 5137
rect 4212 5128 4214 5137
rect 4158 5063 4214 5072
rect 4264 4690 4292 8910
rect 4356 5914 4384 13330
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4816 12832 4844 16934
rect 4908 14521 4936 18958
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 5000 14929 5028 18702
rect 4986 14920 5042 14929
rect 4986 14855 5042 14864
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 4894 14512 4950 14521
rect 4894 14447 4950 14456
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4908 14006 4936 14350
rect 5000 14346 5028 14758
rect 4988 14340 5040 14346
rect 4988 14282 5040 14288
rect 5092 14226 5120 20182
rect 5184 18766 5212 21626
rect 5276 20602 5304 22520
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 5000 14198 5120 14226
rect 4896 14000 4948 14006
rect 4896 13942 4948 13948
rect 4894 13832 4950 13841
rect 4894 13767 4950 13776
rect 4632 12804 4844 12832
rect 4632 12170 4660 12804
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4620 12164 4672 12170
rect 4724 12152 4752 12650
rect 4724 12124 4844 12152
rect 4620 12106 4672 12112
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 4710 11248 4766 11257
rect 4540 11121 4568 11222
rect 4710 11183 4712 11192
rect 4764 11183 4766 11192
rect 4712 11154 4764 11160
rect 4526 11112 4582 11121
rect 4526 11047 4582 11056
rect 4710 11112 4766 11121
rect 4710 11047 4712 11056
rect 4764 11047 4766 11056
rect 4712 11018 4764 11024
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4526 10024 4582 10033
rect 4526 9959 4528 9968
rect 4580 9959 4582 9968
rect 4528 9930 4580 9936
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4816 8974 4844 12124
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4908 8106 4936 13767
rect 5000 9110 5028 14198
rect 5080 14000 5132 14006
rect 5080 13942 5132 13948
rect 5092 12782 5120 13942
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 5078 12608 5134 12617
rect 5078 12543 5134 12552
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 5092 8786 5120 12543
rect 5184 9518 5212 18566
rect 5276 12481 5304 20198
rect 5368 17814 5396 20878
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5460 19718 5488 19994
rect 5736 19922 5764 22520
rect 6196 21026 6224 22520
rect 6196 20998 6500 21026
rect 6276 20868 6328 20874
rect 6276 20810 6328 20816
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5552 18086 5580 19450
rect 5814 19272 5870 19281
rect 5724 19236 5776 19242
rect 5814 19207 5870 19216
rect 5724 19178 5776 19184
rect 5736 18222 5764 19178
rect 5828 19174 5856 19207
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 5632 18216 5684 18222
rect 5632 18158 5684 18164
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5356 17808 5408 17814
rect 5356 17750 5408 17756
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5368 16726 5396 17274
rect 5356 16720 5408 16726
rect 5354 16688 5356 16697
rect 5408 16688 5410 16697
rect 5354 16623 5410 16632
rect 5448 16516 5500 16522
rect 5448 16458 5500 16464
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5368 16046 5396 16390
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5460 15570 5488 16458
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5552 15978 5580 16390
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5460 15026 5488 15506
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5460 14634 5488 14962
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5368 14606 5488 14634
rect 5368 14414 5396 14606
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5354 14240 5410 14249
rect 5354 14175 5410 14184
rect 5262 12472 5318 12481
rect 5262 12407 5318 12416
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 4816 8078 4936 8106
rect 5000 8758 5120 8786
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4710 7440 4766 7449
rect 4710 7375 4766 7384
rect 4724 6798 4752 7375
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4724 5778 4752 6190
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4816 4826 4844 8078
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4908 7546 4936 7890
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4158 4040 4214 4049
rect 4158 3975 4214 3984
rect 4172 3942 4200 3975
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 3974 3567 4030 3576
rect 4068 3596 4120 3602
rect 3988 3398 4016 3567
rect 4068 3538 4120 3544
rect 4250 3496 4306 3505
rect 4250 3431 4252 3440
rect 4304 3431 4306 3440
rect 4252 3402 4304 3408
rect 4816 3398 4844 4082
rect 4908 3738 4936 7278
rect 5000 5166 5028 8758
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5092 4146 5120 6870
rect 5184 5914 5212 9046
rect 5276 7342 5304 11562
rect 5368 7732 5396 14175
rect 5460 12782 5488 14418
rect 5552 14006 5580 14758
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5552 12782 5580 13670
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5460 12481 5488 12718
rect 5446 12472 5502 12481
rect 5446 12407 5502 12416
rect 5552 12050 5580 12718
rect 5460 12022 5580 12050
rect 5460 7834 5488 12022
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5552 11014 5580 11562
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10606 5580 10950
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5552 10198 5580 10542
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5552 8634 5580 9046
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5552 7936 5580 8570
rect 5644 8498 5672 18158
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5736 14929 5764 16526
rect 5722 14920 5778 14929
rect 5722 14855 5778 14864
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5736 12986 5764 13330
rect 5828 13190 5856 18838
rect 6288 17814 6316 20810
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 6276 17808 6328 17814
rect 6276 17750 6328 17756
rect 6196 15366 6224 17750
rect 6276 16720 6328 16726
rect 6276 16662 6328 16668
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6104 14482 6132 15098
rect 6092 14476 6144 14482
rect 6144 14436 6224 14464
rect 6092 14418 6144 14424
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5920 12322 5948 13806
rect 6012 13462 6040 14214
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 6104 13530 6132 14010
rect 6196 13938 6224 14436
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6000 13456 6052 13462
rect 6288 13410 6316 16662
rect 6000 13398 6052 13404
rect 6104 13382 6316 13410
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5828 12294 5948 12322
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5736 10713 5764 10950
rect 5722 10704 5778 10713
rect 5722 10639 5724 10648
rect 5776 10639 5778 10648
rect 5724 10610 5776 10616
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5736 9042 5764 10134
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5552 7908 5672 7936
rect 5460 7806 5580 7834
rect 5368 7704 5488 7732
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5276 7002 5304 7142
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5368 6458 5396 7142
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 3698 3224 3754 3233
rect 4421 3216 4717 3236
rect 3698 3159 3754 3168
rect 5368 2650 5396 6122
rect 5460 5370 5488 7704
rect 5552 6186 5580 7806
rect 5644 6798 5672 7908
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5644 6322 5672 6734
rect 5828 6390 5856 12294
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5920 9178 5948 9386
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5446 5264 5502 5273
rect 5446 5199 5502 5208
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 4080 1737 4108 2586
rect 5460 2446 5488 5199
rect 5644 3466 5672 6122
rect 6012 4826 6040 13262
rect 6104 6934 6132 13382
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6288 12850 6316 13262
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6288 12442 6316 12786
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6380 11937 6408 19790
rect 6472 18714 6500 20998
rect 6656 19258 6684 22520
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6840 19922 6868 20334
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6920 19304 6972 19310
rect 6656 19230 6776 19258
rect 6920 19246 6972 19252
rect 6472 18698 6684 18714
rect 6472 18692 6696 18698
rect 6472 18686 6644 18692
rect 6644 18634 6696 18640
rect 6642 18592 6698 18601
rect 6642 18527 6698 18536
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6564 17678 6592 18226
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6564 15162 6592 17614
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6564 14618 6592 14894
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6458 12472 6514 12481
rect 6458 12407 6514 12416
rect 6366 11928 6422 11937
rect 6366 11863 6422 11872
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6196 9926 6224 11154
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6196 7886 6224 9862
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6104 5642 6132 6870
rect 6380 5778 6408 11863
rect 6472 5914 6500 12407
rect 6564 12374 6592 14010
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6564 11354 6592 12310
rect 6656 11762 6684 18527
rect 6748 18193 6776 19230
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 18902 6868 19110
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6734 18184 6790 18193
rect 6734 18119 6790 18128
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6748 13818 6776 17750
rect 6840 17542 6868 18702
rect 6932 18222 6960 19246
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 7116 17592 7144 22520
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7300 19854 7328 20402
rect 7288 19848 7340 19854
rect 7340 19808 7420 19836
rect 7288 19790 7340 19796
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7300 19310 7328 19654
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7208 19009 7236 19110
rect 7194 19000 7250 19009
rect 7194 18935 7250 18944
rect 7392 18816 7420 19808
rect 7208 18788 7420 18816
rect 7208 18154 7236 18788
rect 7380 18692 7432 18698
rect 7380 18634 7432 18640
rect 7196 18148 7248 18154
rect 7196 18090 7248 18096
rect 7208 17882 7236 18090
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7116 17564 7328 17592
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6918 17504 6974 17513
rect 6840 15638 6868 17478
rect 6918 17439 6974 17448
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6748 13790 6868 13818
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6656 10130 6684 11562
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6564 9178 6592 10066
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6564 7818 6592 9114
rect 6656 7857 6684 9522
rect 6748 8634 6776 12650
rect 6840 12481 6868 13790
rect 6826 12472 6882 12481
rect 6826 12407 6882 12416
rect 6932 12102 6960 17439
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6840 8498 6868 11290
rect 6932 11218 6960 11630
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 7024 7970 7052 16934
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 7116 14958 7144 15506
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7116 13530 7144 14894
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7208 12442 7236 16934
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7116 10470 7144 11290
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7208 9194 7236 12242
rect 7300 10554 7328 17564
rect 7392 17202 7420 18634
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7392 16590 7420 17138
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7576 16250 7604 22520
rect 8036 20346 8064 22520
rect 8298 20360 8354 20369
rect 8036 20318 8298 20346
rect 8298 20295 8354 20304
rect 8496 20262 8524 22520
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 8208 20256 8260 20262
rect 8484 20256 8536 20262
rect 8208 20198 8260 20204
rect 8482 20224 8484 20233
rect 8536 20224 8538 20233
rect 7668 19666 7696 20198
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 7668 19638 7788 19666
rect 7760 19446 7788 19638
rect 8220 19530 8248 20198
rect 8482 20159 8538 20168
rect 8482 19952 8538 19961
rect 8482 19887 8538 19896
rect 8390 19816 8446 19825
rect 8390 19751 8446 19760
rect 8404 19666 8432 19751
rect 8036 19502 8248 19530
rect 8312 19638 8432 19666
rect 8312 19514 8340 19638
rect 8300 19508 8352 19514
rect 7748 19440 7800 19446
rect 7748 19382 7800 19388
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7668 18766 7696 19246
rect 7656 18760 7708 18766
rect 7656 18702 7708 18708
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7668 17338 7696 17614
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7392 14278 7420 14962
rect 7484 14550 7512 15370
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7392 13870 7420 14214
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7484 10554 7512 12378
rect 7576 11098 7604 15914
rect 7760 15201 7788 19382
rect 8036 19156 8064 19502
rect 8300 19450 8352 19456
rect 8392 19440 8444 19446
rect 8496 19428 8524 19887
rect 8680 19446 8708 20742
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 8772 20262 8800 20538
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 8850 20224 8906 20233
rect 8444 19400 8524 19428
rect 8668 19440 8720 19446
rect 8392 19382 8444 19388
rect 8668 19382 8720 19388
rect 8208 19304 8260 19310
rect 8206 19272 8208 19281
rect 8576 19304 8628 19310
rect 8260 19272 8262 19281
rect 8206 19207 8262 19216
rect 8482 19272 8538 19281
rect 8576 19246 8628 19252
rect 8482 19207 8484 19216
rect 8536 19207 8538 19216
rect 8484 19178 8536 19184
rect 8036 19128 8248 19156
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 8220 18970 8248 19128
rect 8298 19136 8354 19145
rect 8298 19071 8354 19080
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8208 18692 8260 18698
rect 8208 18634 8260 18640
rect 8220 18086 8248 18634
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8220 17814 8248 18022
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8128 17542 8156 17682
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8312 17218 8340 19071
rect 8484 18692 8536 18698
rect 8484 18634 8536 18640
rect 8496 17610 8524 18634
rect 8588 18601 8616 19246
rect 8772 18902 8800 20198
rect 8850 20159 8906 20168
rect 8760 18896 8812 18902
rect 8760 18838 8812 18844
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8574 18592 8630 18601
rect 8574 18527 8630 18536
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8312 17190 8432 17218
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 8206 16688 8262 16697
rect 8312 16658 8340 17002
rect 8206 16623 8262 16632
rect 8300 16652 8352 16658
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8128 16046 8156 16390
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 7746 15192 7802 15201
rect 7746 15127 7802 15136
rect 7748 15088 7800 15094
rect 7748 15030 7800 15036
rect 7760 14056 7788 15030
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7840 14068 7892 14074
rect 7760 14028 7840 14056
rect 7656 13252 7708 13258
rect 7656 13194 7708 13200
rect 7668 12170 7696 13194
rect 7760 12306 7788 14028
rect 7840 14010 7892 14016
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8220 12424 8248 16623
rect 8300 16594 8352 16600
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8312 15706 8340 15982
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8404 14822 8432 17190
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 8404 14634 8432 14758
rect 8312 14606 8432 14634
rect 8312 13802 8340 14606
rect 8300 13796 8352 13802
rect 8300 13738 8352 13744
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8036 12396 8248 12424
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 8036 11676 8064 12396
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8220 11898 8248 12242
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8036 11648 8248 11676
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7576 11070 7696 11098
rect 7760 11082 7788 11494
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7576 10674 7604 10950
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7300 10526 7420 10554
rect 7484 10526 7604 10554
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7300 9382 7328 10406
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7208 9166 7328 9194
rect 7194 8800 7250 8809
rect 7194 8735 7250 8744
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6932 7942 7052 7970
rect 6642 7848 6698 7857
rect 6552 7812 6604 7818
rect 6642 7783 6698 7792
rect 6552 7754 6604 7760
rect 6564 7410 6592 7754
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6656 5574 6684 7783
rect 6840 7546 6868 7890
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5828 3194 5856 3402
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4066 1728 4122 1737
rect 4066 1663 4122 1672
rect 5920 1290 5948 3674
rect 6932 2310 6960 7942
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7024 7002 7052 7822
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 7116 5234 7144 8366
rect 7208 7313 7236 8735
rect 7194 7304 7250 7313
rect 7194 7239 7250 7248
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7208 6322 7236 7142
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 5846 7236 6258
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 7116 1442 7144 2858
rect 7300 2854 7328 9166
rect 7392 8974 7420 10526
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7392 8242 7420 8910
rect 7484 8412 7512 10406
rect 7576 9586 7604 10526
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7576 8566 7604 9386
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7484 8384 7604 8412
rect 7392 8214 7512 8242
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7392 6730 7420 7346
rect 7484 6866 7512 8214
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7470 6760 7526 6769
rect 7380 6724 7432 6730
rect 7470 6695 7526 6704
rect 7380 6666 7432 6672
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7484 2038 7512 6695
rect 7576 5370 7604 8384
rect 7668 6254 7696 11070
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7760 10198 7788 11018
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7760 8838 7788 9454
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7746 8664 7802 8673
rect 7746 8599 7802 8608
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7760 4826 7788 8599
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7838 7440 7894 7449
rect 7838 7375 7840 7384
rect 7892 7375 7894 7384
rect 7840 7346 7892 7352
rect 8220 7313 8248 11648
rect 8312 10418 8340 13126
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8404 10606 8432 12310
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8496 10810 8524 12174
rect 8588 11354 8616 16186
rect 8680 12374 8708 18702
rect 8864 18698 8892 20159
rect 8956 19990 8984 22520
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 9048 19990 9076 20334
rect 8944 19984 8996 19990
rect 8944 19926 8996 19932
rect 9036 19984 9088 19990
rect 9036 19926 9088 19932
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8758 18184 8814 18193
rect 8758 18119 8814 18128
rect 9218 18184 9274 18193
rect 9218 18119 9220 18128
rect 8772 13734 8800 18119
rect 9272 18119 9274 18128
rect 9220 18090 9272 18096
rect 9128 18080 9180 18086
rect 9324 18034 9352 20538
rect 9128 18022 9180 18028
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8864 15026 8892 15642
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8852 15020 8904 15026
rect 8852 14962 8904 14968
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8772 12782 8800 13262
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8680 11218 8708 12106
rect 8758 11792 8814 11801
rect 8758 11727 8814 11736
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8772 11082 8800 11727
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8588 10742 8616 10950
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8312 10390 8432 10418
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8312 9178 8340 9998
rect 8404 9761 8432 10390
rect 8496 10266 8524 10610
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8390 9752 8446 9761
rect 8390 9687 8446 9696
rect 8482 9616 8538 9625
rect 8482 9551 8538 9560
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8404 9042 8432 9114
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8206 7304 8262 7313
rect 8206 7239 8262 7248
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8404 7002 8432 8978
rect 8496 8294 8524 9551
rect 8588 9110 8616 10678
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8576 8968 8628 8974
rect 8574 8936 8576 8945
rect 8628 8936 8630 8945
rect 8574 8871 8630 8880
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8208 6928 8260 6934
rect 8114 6896 8170 6905
rect 8208 6870 8260 6876
rect 8390 6896 8446 6905
rect 8114 6831 8170 6840
rect 8128 6474 8156 6831
rect 8220 6662 8248 6870
rect 8390 6831 8392 6840
rect 8444 6831 8446 6840
rect 8392 6802 8444 6808
rect 8390 6760 8446 6769
rect 8390 6695 8446 6704
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8128 6446 8248 6474
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8036 5166 8064 5510
rect 8220 5370 8248 6446
rect 8404 6390 8432 6695
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 8036 5012 8064 5102
rect 8208 5024 8260 5030
rect 8036 4984 8208 5012
rect 8208 4966 8260 4972
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 8312 4729 8340 6054
rect 8404 4826 8432 6054
rect 8496 5778 8524 7414
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8588 5386 8616 8366
rect 8680 6118 8708 10202
rect 8772 8838 8800 10542
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 8498 8800 8774
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8758 8392 8814 8401
rect 8758 8327 8760 8336
rect 8812 8327 8814 8336
rect 8760 8298 8812 8304
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8772 6254 8800 6734
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8680 5778 8708 5850
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8666 5672 8722 5681
rect 8666 5607 8722 5616
rect 8680 5574 8708 5607
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8588 5358 8708 5386
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8298 4720 8354 4729
rect 8298 4655 8354 4664
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 8220 3641 8248 3878
rect 8206 3632 8262 3641
rect 8206 3567 8262 3576
rect 8588 3126 8616 5170
rect 8680 3670 8708 5358
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8772 2990 8800 6190
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7576 2825 7604 2858
rect 7562 2816 7618 2825
rect 7562 2751 7618 2760
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 7472 2032 7524 2038
rect 7472 1974 7524 1980
rect 8864 1766 8892 14350
rect 8956 3942 8984 15506
rect 9036 14544 9088 14550
rect 9036 14486 9088 14492
rect 9048 14074 9076 14486
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 13258 9076 13670
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 9140 13138 9168 18022
rect 9232 18006 9352 18034
rect 9232 16776 9260 18006
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9324 16969 9352 17274
rect 9416 17066 9444 22520
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9508 19310 9536 19790
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 9508 18222 9536 19246
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9310 16960 9366 16969
rect 9310 16895 9366 16904
rect 9232 16748 9444 16776
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9048 13110 9168 13138
rect 9048 9178 9076 13110
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9140 11801 9168 12174
rect 9126 11792 9182 11801
rect 9126 11727 9182 11736
rect 9232 11642 9260 16594
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9324 14006 9352 15302
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 9324 11898 9352 13194
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9416 11744 9444 16748
rect 9508 15706 9536 18158
rect 9600 17338 9628 18566
rect 9692 17882 9720 18770
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9600 16658 9628 17274
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9588 16176 9640 16182
rect 9588 16118 9640 16124
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9508 14482 9536 15642
rect 9600 14958 9628 16118
rect 9678 15736 9734 15745
rect 9678 15671 9680 15680
rect 9732 15671 9734 15680
rect 9680 15642 9732 15648
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9508 13376 9536 14282
rect 9586 13832 9642 13841
rect 9586 13767 9642 13776
rect 9600 13734 9628 13767
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9508 13348 9628 13376
rect 9494 13288 9550 13297
rect 9494 13223 9550 13232
rect 9508 12374 9536 13223
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9140 11614 9260 11642
rect 9324 11716 9444 11744
rect 9140 10810 9168 11614
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9324 11506 9352 11716
rect 9600 11665 9628 13348
rect 9692 12714 9720 14418
rect 9876 13734 9904 22520
rect 10336 18086 10364 22520
rect 10796 20346 10824 22520
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 10416 20324 10468 20330
rect 10416 20266 10468 20272
rect 10612 20318 10824 20346
rect 10428 20058 10456 20266
rect 10416 20052 10468 20058
rect 10416 19994 10468 20000
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 10428 18358 10456 18906
rect 10612 18766 10640 20318
rect 10692 20256 10744 20262
rect 10968 20256 11020 20262
rect 10692 20198 10744 20204
rect 10966 20224 10968 20233
rect 11020 20224 11022 20233
rect 10704 18970 10732 20198
rect 10966 20159 11022 20168
rect 11072 19854 11100 20402
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 11072 19718 11100 19790
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10796 18766 10824 19110
rect 10600 18760 10652 18766
rect 10506 18728 10562 18737
rect 10600 18702 10652 18708
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 10506 18663 10562 18672
rect 10416 18352 10468 18358
rect 10416 18294 10468 18300
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10428 17898 10456 18294
rect 10244 17882 10456 17898
rect 10232 17876 10456 17882
rect 10284 17870 10456 17876
rect 10232 17818 10284 17824
rect 10416 17808 10468 17814
rect 10336 17768 10416 17796
rect 10336 17762 10364 17768
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 10152 17734 10364 17762
rect 10416 17750 10468 17756
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9876 13394 9904 13670
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9692 12306 9720 12650
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9784 11880 9812 12650
rect 9968 12458 9996 17682
rect 10152 17678 10180 17734
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10244 17270 10272 17478
rect 10140 17264 10192 17270
rect 10140 17206 10192 17212
rect 10232 17264 10284 17270
rect 10232 17206 10284 17212
rect 10152 15502 10180 17206
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10244 15994 10272 16118
rect 10336 16114 10364 16934
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10244 15966 10364 15994
rect 10336 15502 10364 15966
rect 10416 15972 10468 15978
rect 10416 15914 10468 15920
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10428 14226 10456 15914
rect 9959 12430 9996 12458
rect 10152 14198 10456 14226
rect 9959 12424 9987 12430
rect 9692 11852 9812 11880
rect 9876 12396 9987 12424
rect 9586 11656 9642 11665
rect 9586 11591 9642 11600
rect 9692 11540 9720 11852
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9600 11512 9720 11540
rect 9600 11506 9628 11512
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9140 9722 9168 10474
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 9048 8430 9076 8842
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 6866 9076 8230
rect 9140 7342 9168 9114
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9036 6180 9088 6186
rect 9036 6122 9088 6128
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 9048 5234 9076 6122
rect 9140 5778 9168 6122
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9128 5568 9180 5574
rect 9126 5536 9128 5545
rect 9180 5536 9182 5545
rect 9126 5471 9182 5480
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 9048 4078 9076 4422
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 9232 3210 9260 11494
rect 9324 11478 9444 11506
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 10470 9352 10950
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9324 8430 9352 8978
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9324 6798 9352 8366
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9310 6352 9366 6361
rect 9310 6287 9366 6296
rect 9324 5846 9352 6287
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9324 5302 9352 5646
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9140 3182 9260 3210
rect 9140 2650 9168 3182
rect 9324 3058 9352 5034
rect 9416 4690 9444 11478
rect 9508 11478 9628 11506
rect 9508 11150 9536 11478
rect 9586 11384 9642 11393
rect 9784 11354 9812 11698
rect 9876 11642 9904 12396
rect 10048 12368 10100 12374
rect 9968 12328 10048 12356
rect 9968 11762 9996 12328
rect 10048 12310 10100 12316
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10060 11762 10088 12038
rect 10152 11778 10180 14198
rect 10414 13968 10470 13977
rect 10414 13903 10470 13912
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10244 12986 10272 13262
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 10244 12374 10272 12922
rect 10428 12918 10456 13903
rect 10520 13802 10548 18663
rect 10600 18624 10652 18630
rect 10600 18566 10652 18572
rect 10508 13796 10560 13802
rect 10508 13738 10560 13744
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10232 12368 10284 12374
rect 10232 12310 10284 12316
rect 10414 11792 10470 11801
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 10048 11756 10100 11762
rect 10152 11750 10364 11778
rect 10048 11698 10100 11704
rect 10232 11688 10284 11694
rect 9876 11614 10088 11642
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9586 11319 9642 11328
rect 9772 11348 9824 11354
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9508 9178 9536 10746
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9600 9058 9628 11319
rect 9772 11290 9824 11296
rect 9770 11248 9826 11257
rect 9770 11183 9826 11192
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9508 9030 9628 9058
rect 9508 8242 9536 9030
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9600 8362 9628 8910
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9508 8214 9628 8242
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9600 7290 9628 8214
rect 9692 7954 9720 10474
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9678 7304 9734 7313
rect 9508 5370 9536 7278
rect 9600 7262 9678 7290
rect 9678 7239 9734 7248
rect 9588 7200 9640 7206
rect 9784 7177 9812 11183
rect 9876 7818 9904 11494
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9968 7954 9996 11154
rect 10060 9178 10088 11614
rect 10152 11636 10232 11642
rect 10152 11630 10284 11636
rect 10152 11614 10272 11630
rect 10152 10606 10180 11614
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10244 11121 10272 11222
rect 10230 11112 10286 11121
rect 10230 11047 10286 11056
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10336 8786 10364 11750
rect 10414 11727 10470 11736
rect 10428 11694 10456 11727
rect 10416 11688 10468 11694
rect 10520 11665 10548 12582
rect 10416 11630 10468 11636
rect 10506 11656 10562 11665
rect 10428 10810 10456 11630
rect 10506 11591 10562 11600
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10428 9586 10456 9862
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10060 8758 10364 8786
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9588 7142 9640 7148
rect 9770 7168 9826 7177
rect 9600 7041 9628 7142
rect 9770 7103 9826 7112
rect 9586 7032 9642 7041
rect 9586 6967 9588 6976
rect 9640 6967 9642 6976
rect 9588 6938 9640 6944
rect 9600 6907 9628 6938
rect 9968 6866 9996 7346
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9586 6080 9642 6089
rect 9586 6015 9642 6024
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9600 4486 9628 6015
rect 9784 5098 9812 6802
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9876 6118 9904 6326
rect 9968 6118 9996 6802
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9954 5944 10010 5953
rect 9954 5879 10010 5888
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9784 4865 9812 5034
rect 9770 4856 9826 4865
rect 9770 4791 9826 4800
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9678 4312 9734 4321
rect 9600 4270 9678 4298
rect 9600 3097 9628 4270
rect 9678 4247 9734 4256
rect 9876 4214 9904 5510
rect 9968 4690 9996 5879
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 10060 4282 10088 8758
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10230 8528 10286 8537
rect 10230 8463 10286 8472
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 10046 4176 10102 4185
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3738 9720 3878
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9876 3602 9904 4150
rect 10046 4111 10102 4120
rect 10060 4010 10088 4111
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10046 3768 10102 3777
rect 10046 3703 10048 3712
rect 10100 3703 10102 3712
rect 10048 3674 10100 3680
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9586 3088 9642 3097
rect 9312 3052 9364 3058
rect 9586 3023 9642 3032
rect 9312 2994 9364 3000
rect 10152 2990 10180 7822
rect 10244 6458 10272 8463
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10244 5710 10272 6190
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10244 5273 10272 5646
rect 10336 5302 10364 8570
rect 10428 6254 10456 9318
rect 10520 8090 10548 9862
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10428 5710 10456 6054
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10324 5296 10376 5302
rect 10230 5264 10286 5273
rect 10324 5238 10376 5244
rect 10230 5199 10286 5208
rect 10428 5137 10456 5646
rect 10414 5128 10470 5137
rect 10414 5063 10470 5072
rect 10322 4992 10378 5001
rect 10322 4927 10378 4936
rect 10336 4826 10364 4927
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 10322 4584 10378 4593
rect 10322 4519 10378 4528
rect 10336 4282 10364 4519
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10520 4010 10548 7890
rect 10612 6254 10640 18566
rect 10796 18222 10824 18702
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10704 17202 10732 18022
rect 10888 17649 10916 19654
rect 11072 19242 11100 19654
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10980 18358 11008 19110
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 10968 18352 11020 18358
rect 10968 18294 11020 18300
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10874 17640 10930 17649
rect 10874 17575 10930 17584
rect 10980 17513 11008 18158
rect 11072 17678 11100 18702
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 10966 17504 11022 17513
rect 10966 17439 11022 17448
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10704 16046 10732 17138
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10704 15502 10732 15982
rect 10888 15978 10916 16934
rect 10968 16788 11020 16794
rect 11072 16776 11100 17614
rect 11256 17320 11284 22520
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11532 18766 11560 19246
rect 11716 19174 11744 22520
rect 12176 20398 12204 22520
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12348 20256 12400 20262
rect 12346 20224 12348 20233
rect 12400 20224 12402 20233
rect 12346 20159 12402 20168
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11610 19000 11666 19009
rect 11610 18935 11666 18944
rect 11624 18834 11652 18935
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11716 18426 11744 18770
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11518 17912 11574 17921
rect 11716 17882 11744 18362
rect 11518 17847 11574 17856
rect 11704 17876 11756 17882
rect 11532 17610 11560 17847
rect 11704 17818 11756 17824
rect 11520 17604 11572 17610
rect 11520 17546 11572 17552
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11020 16748 11100 16776
rect 11164 17292 11284 17320
rect 10968 16730 11020 16736
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10704 14006 10732 14962
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10690 13560 10746 13569
rect 10690 13495 10692 13504
rect 10744 13495 10746 13504
rect 10692 13466 10744 13472
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10704 12986 10732 13330
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10704 9450 10732 12582
rect 10796 12374 10824 15574
rect 10784 12368 10836 12374
rect 10888 12345 10916 15914
rect 10980 14396 11008 16730
rect 11164 15638 11192 17292
rect 11242 17232 11298 17241
rect 11242 17167 11298 17176
rect 11256 16454 11284 17167
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11518 15600 11574 15609
rect 11518 15535 11520 15544
rect 11572 15535 11574 15544
rect 11520 15506 11572 15512
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11072 14890 11100 15302
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11610 15056 11666 15065
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 11164 14482 11192 15030
rect 11610 14991 11666 15000
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11060 14408 11112 14414
rect 10980 14368 11060 14396
rect 11256 14385 11284 14894
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11348 14657 11376 14758
rect 11334 14648 11390 14657
rect 11334 14583 11390 14592
rect 11624 14414 11652 14991
rect 11612 14408 11664 14414
rect 11060 14350 11112 14356
rect 11242 14376 11298 14385
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10784 12310 10836 12316
rect 10874 12336 10930 12345
rect 10874 12271 10930 12280
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10704 6769 10732 9114
rect 10796 8090 10824 10066
rect 10888 8974 10916 10134
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10888 8634 10916 8910
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10782 7984 10838 7993
rect 10782 7919 10838 7928
rect 10690 6760 10746 6769
rect 10690 6695 10746 6704
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10704 5234 10732 5850
rect 10796 5574 10824 7919
rect 10888 7750 10916 8026
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10874 6216 10930 6225
rect 10874 6151 10930 6160
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10782 4992 10838 5001
rect 10782 4927 10838 4936
rect 10796 4078 10824 4927
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10690 3904 10746 3913
rect 10690 3839 10746 3848
rect 10704 3602 10732 3839
rect 10888 3670 10916 6151
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10612 2922 10640 3470
rect 10980 3194 11008 13466
rect 11072 13326 11100 14350
rect 11612 14350 11664 14356
rect 11242 14311 11298 14320
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 11164 12730 11192 13738
rect 11256 12850 11284 14214
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11716 14006 11744 17002
rect 11704 14000 11756 14006
rect 11704 13942 11756 13948
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11348 13462 11376 13874
rect 11336 13456 11388 13462
rect 11520 13456 11572 13462
rect 11336 13398 11388 13404
rect 11518 13424 11520 13433
rect 11572 13424 11574 13433
rect 11518 13359 11574 13368
rect 11808 13161 11836 19110
rect 11900 18902 11928 19654
rect 11980 19236 12032 19242
rect 11980 19178 12032 19184
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 11888 17740 11940 17746
rect 11992 17728 12020 19178
rect 12162 18864 12218 18873
rect 12162 18799 12218 18808
rect 11940 17700 12020 17728
rect 11888 17682 11940 17688
rect 11992 16794 12020 17700
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11992 16266 12020 16594
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 11900 16250 12020 16266
rect 11888 16244 12020 16250
rect 11940 16238 12020 16244
rect 11888 16186 11940 16192
rect 12084 15978 12112 16526
rect 12072 15972 12124 15978
rect 12072 15914 12124 15920
rect 12176 15688 12204 18799
rect 12452 18426 12480 19926
rect 12530 19000 12586 19009
rect 12530 18935 12532 18944
rect 12584 18935 12586 18944
rect 12532 18906 12584 18912
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12348 17740 12400 17746
rect 12636 17728 12664 22520
rect 13096 20618 13124 22520
rect 13096 20590 13492 20618
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12912 17814 12940 18226
rect 12716 17808 12768 17814
rect 12348 17682 12400 17688
rect 12452 17700 12664 17728
rect 12714 17776 12716 17785
rect 12900 17808 12952 17814
rect 12768 17776 12770 17785
rect 12900 17750 12952 17756
rect 12714 17711 12770 17720
rect 12808 17740 12860 17746
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 11992 15660 12204 15688
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 11900 13802 11928 15574
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11794 13152 11850 13161
rect 11352 13084 11648 13104
rect 11794 13087 11850 13096
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11072 12617 11100 12718
rect 11164 12702 11284 12730
rect 11058 12608 11114 12617
rect 11058 12543 11114 12552
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11072 12345 11100 12378
rect 11058 12336 11114 12345
rect 11058 12271 11114 12280
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11058 11928 11114 11937
rect 11058 11863 11060 11872
rect 11112 11863 11114 11872
rect 11060 11834 11112 11840
rect 11164 11370 11192 12106
rect 11072 11342 11192 11370
rect 11072 9926 11100 11342
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11072 9178 11100 9386
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11060 8016 11112 8022
rect 11164 8004 11192 11086
rect 11112 7976 11192 8004
rect 11060 7958 11112 7964
rect 11256 7954 11284 12702
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11348 12170 11376 12378
rect 11440 12345 11468 12650
rect 11704 12368 11756 12374
rect 11426 12336 11482 12345
rect 11704 12310 11756 12316
rect 11426 12271 11482 12280
rect 11336 12164 11388 12170
rect 11336 12106 11388 12112
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11624 11393 11652 11494
rect 11610 11384 11666 11393
rect 11610 11319 11666 11328
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11716 9704 11744 12310
rect 11624 9676 11744 9704
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 11532 9081 11560 9590
rect 11624 9353 11652 9676
rect 11808 9568 11836 12922
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11716 9540 11836 9568
rect 11610 9344 11666 9353
rect 11610 9279 11666 9288
rect 11610 9208 11666 9217
rect 11610 9143 11666 9152
rect 11518 9072 11574 9081
rect 11624 9042 11652 9143
rect 11518 9007 11574 9016
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11348 7886 11376 8298
rect 11716 8022 11744 9540
rect 11900 9466 11928 12854
rect 11808 9438 11928 9466
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11702 7848 11758 7857
rect 11702 7783 11704 7792
rect 11756 7783 11758 7792
rect 11704 7754 11756 7760
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11244 7472 11296 7478
rect 11296 7432 11376 7460
rect 11244 7414 11296 7420
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 6254 11100 7142
rect 11164 7002 11192 7346
rect 11348 7274 11376 7432
rect 11336 7268 11388 7274
rect 11336 7210 11388 7216
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 5370 11100 6054
rect 11164 5953 11192 6938
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11256 6440 11284 6802
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11256 6412 11376 6440
rect 11150 5944 11206 5953
rect 11150 5879 11206 5888
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11164 5642 11192 5782
rect 11348 5710 11376 6412
rect 11518 5944 11574 5953
rect 11518 5879 11574 5888
rect 11532 5846 11560 5879
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11152 5636 11204 5642
rect 11152 5578 11204 5584
rect 11532 5556 11560 5782
rect 11256 5528 11560 5556
rect 11256 5522 11284 5528
rect 11164 5494 11284 5522
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11164 5114 11192 5494
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11716 5370 11744 7142
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11348 5114 11376 5170
rect 11716 5137 11744 5170
rect 11164 5086 11376 5114
rect 11702 5128 11758 5137
rect 11702 5063 11758 5072
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11072 4826 11100 4966
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11242 4720 11298 4729
rect 11060 4684 11112 4690
rect 11242 4655 11298 4664
rect 11060 4626 11112 4632
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10508 2916 10560 2922
rect 10508 2858 10560 2864
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 8852 1760 8904 1766
rect 8852 1702 8904 1708
rect 10520 1630 10548 2858
rect 11072 2650 11100 4626
rect 11256 2990 11284 4655
rect 11532 4622 11560 4762
rect 11716 4622 11744 5063
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11808 3194 11836 9438
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 9178 11928 9318
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11256 1986 11284 2790
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11256 1958 11560 1986
rect 10508 1624 10560 1630
rect 10508 1566 10560 1572
rect 6932 1414 7144 1442
rect 5908 1284 5960 1290
rect 5908 1226 5960 1232
rect 3606 640 3662 649
rect 3606 575 3662 584
rect 6932 480 6960 1414
rect 11532 480 11560 1958
rect 3238 232 3294 241
rect 3238 167 3294 176
rect 6918 0 6974 480
rect 11518 0 11574 480
rect 11900 241 11928 7890
rect 11992 3738 12020 15660
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12084 12986 12112 15506
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12176 14090 12204 15438
rect 12268 15094 12296 16458
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12176 14062 12296 14090
rect 12164 14000 12216 14006
rect 12162 13968 12164 13977
rect 12216 13968 12218 13977
rect 12162 13903 12218 13912
rect 12268 13705 12296 14062
rect 12254 13696 12310 13705
rect 12254 13631 12310 13640
rect 12360 13546 12388 17682
rect 12452 16454 12480 17700
rect 12808 17682 12860 17688
rect 12622 17640 12678 17649
rect 12622 17575 12624 17584
rect 12676 17575 12678 17584
rect 12624 17546 12676 17552
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 17338 12572 17478
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 15706 12480 16390
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12438 15056 12494 15065
rect 12438 14991 12440 15000
rect 12492 14991 12494 15000
rect 12440 14962 12492 14968
rect 12438 14920 12494 14929
rect 12438 14855 12494 14864
rect 12452 14822 12480 14855
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12176 13518 12388 13546
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12070 12880 12126 12889
rect 12070 12815 12126 12824
rect 12084 12442 12112 12815
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12070 12336 12126 12345
rect 12070 12271 12126 12280
rect 12084 10169 12112 12271
rect 12070 10160 12126 10169
rect 12070 10095 12126 10104
rect 12070 9208 12126 9217
rect 12070 9143 12126 9152
rect 12084 9110 12112 9143
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11992 3194 12020 3334
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12084 1193 12112 7958
rect 12176 3738 12204 13518
rect 12452 13190 12480 14418
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12440 12640 12492 12646
rect 12346 12608 12402 12617
rect 12440 12582 12492 12588
rect 12346 12543 12402 12552
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12268 11354 12296 12174
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12360 11098 12388 12543
rect 12452 11218 12480 12582
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12256 11076 12308 11082
rect 12360 11070 12480 11098
rect 12256 11018 12308 11024
rect 12268 10985 12296 11018
rect 12254 10976 12310 10985
rect 12254 10911 12310 10920
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12360 10266 12388 10474
rect 12452 10470 12480 11070
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10266 12480 10406
rect 12348 10260 12400 10266
rect 12268 10220 12348 10248
rect 12268 8566 12296 10220
rect 12348 10202 12400 10208
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12438 10160 12494 10169
rect 12438 10095 12494 10104
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12360 8412 12388 9998
rect 12452 8945 12480 10095
rect 12438 8936 12494 8945
rect 12438 8871 12494 8880
rect 12268 8384 12388 8412
rect 12440 8424 12492 8430
rect 12268 8022 12296 8384
rect 12440 8366 12492 8372
rect 12348 8288 12400 8294
rect 12348 8230 12400 8236
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 12360 7886 12388 8230
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12268 6610 12296 7686
rect 12360 6866 12388 7822
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12268 6582 12388 6610
rect 12360 5692 12388 6582
rect 12452 6458 12480 8366
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12268 5664 12388 5692
rect 12268 4078 12296 5664
rect 12452 5409 12480 6258
rect 12438 5400 12494 5409
rect 12438 5335 12494 5344
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12360 4826 12388 4966
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12452 4554 12480 5034
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12360 4146 12388 4218
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12544 3890 12572 16934
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12636 15065 12664 15982
rect 12622 15056 12678 15065
rect 12622 14991 12678 15000
rect 12728 14550 12756 17002
rect 12820 16794 12848 17682
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 12716 14544 12768 14550
rect 12716 14486 12768 14492
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12728 13802 12756 13874
rect 12900 13864 12952 13870
rect 12898 13832 12900 13841
rect 12952 13832 12954 13841
rect 12716 13796 12768 13802
rect 12898 13767 12954 13776
rect 12716 13738 12768 13744
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 13004 13569 13032 13670
rect 12990 13560 13046 13569
rect 12990 13495 13046 13504
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12636 12850 12664 13330
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12622 12744 12678 12753
rect 12622 12679 12678 12688
rect 12636 12170 12664 12679
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12636 10130 12664 12106
rect 12728 11626 12756 12786
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 12820 10810 12848 12582
rect 12898 12336 12954 12345
rect 12898 12271 12954 12280
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12728 9994 12756 10678
rect 12912 10198 12940 12271
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12636 9110 12664 9862
rect 12820 9722 12848 9862
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12728 8838 12756 9046
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12636 7750 12664 8502
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12636 5778 12664 7482
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12728 7002 12756 7142
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12728 6322 12756 6666
rect 12820 6633 12848 9454
rect 12912 8566 12940 9658
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12806 6624 12862 6633
rect 12806 6559 12862 6568
rect 12806 6352 12862 6361
rect 12716 6316 12768 6322
rect 12806 6287 12862 6296
rect 12716 6258 12768 6264
rect 12728 5914 12756 6258
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12636 4593 12664 5102
rect 12622 4584 12678 4593
rect 12622 4519 12678 4528
rect 12714 4312 12770 4321
rect 12714 4247 12770 4256
rect 12452 3738 12480 3878
rect 12544 3862 12664 3890
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12636 3670 12664 3862
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12452 3126 12480 3334
rect 12440 3120 12492 3126
rect 12624 3120 12676 3126
rect 12440 3062 12492 3068
rect 12622 3088 12624 3097
rect 12676 3088 12678 3097
rect 12622 3023 12678 3032
rect 12728 2990 12756 4247
rect 12820 4185 12848 6287
rect 12806 4176 12862 4185
rect 12806 4111 12862 4120
rect 12912 4026 12940 8298
rect 13004 4146 13032 12582
rect 13096 12345 13124 15506
rect 13188 15042 13216 20198
rect 13280 19786 13308 20402
rect 13268 19780 13320 19786
rect 13268 19722 13320 19728
rect 13280 18698 13308 19722
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 13280 18290 13308 18634
rect 13372 18329 13400 20402
rect 13358 18320 13414 18329
rect 13268 18284 13320 18290
rect 13358 18255 13414 18264
rect 13268 18226 13320 18232
rect 13266 17912 13322 17921
rect 13266 17847 13268 17856
rect 13320 17847 13322 17856
rect 13268 17818 13320 17824
rect 13372 17377 13400 18255
rect 13358 17368 13414 17377
rect 13358 17303 13414 17312
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13188 15014 13308 15042
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13188 14657 13216 14826
rect 13174 14648 13230 14657
rect 13174 14583 13230 14592
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13188 13938 13216 14214
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13082 12336 13138 12345
rect 13082 12271 13138 12280
rect 13188 12209 13216 13126
rect 13280 12714 13308 15014
rect 13372 14482 13400 17138
rect 13464 14906 13492 20590
rect 13556 18426 13584 22520
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 13924 19990 13952 20538
rect 13912 19984 13964 19990
rect 13912 19926 13964 19932
rect 14016 19174 14044 22520
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14384 19922 14412 20334
rect 14372 19916 14424 19922
rect 14372 19858 14424 19864
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14108 18834 14136 19722
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 14108 18737 14136 18770
rect 14094 18728 14150 18737
rect 14094 18663 14150 18672
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13544 18148 13596 18154
rect 13544 18090 13596 18096
rect 13636 18148 13688 18154
rect 13636 18090 13688 18096
rect 13832 18142 14320 18170
rect 13556 17377 13584 18090
rect 13542 17368 13598 17377
rect 13542 17303 13598 17312
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13556 15745 13584 16662
rect 13542 15736 13598 15745
rect 13542 15671 13598 15680
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13556 15026 13584 15438
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13464 14878 13584 14906
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13464 14346 13492 14758
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 13174 12200 13230 12209
rect 13174 12135 13230 12144
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13096 11694 13124 12038
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13096 10674 13124 11494
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12820 3998 12940 4026
rect 12820 3534 12848 3998
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12912 3738 12940 3878
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 13096 1358 13124 10406
rect 13188 8362 13216 12038
rect 13280 10470 13308 12650
rect 13372 12617 13400 14214
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13464 13274 13492 13942
rect 13556 13394 13584 14878
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13464 13246 13584 13274
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13464 12782 13492 13126
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13358 12608 13414 12617
rect 13358 12543 13414 12552
rect 13358 12472 13414 12481
rect 13358 12407 13414 12416
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 13280 8294 13308 10134
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13372 7936 13400 12407
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13464 9518 13492 11630
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13464 8430 13492 9454
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13188 7908 13400 7936
rect 13188 7342 13216 7908
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13188 5166 13216 7278
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13280 2650 13308 7278
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 7041 13400 7142
rect 13358 7032 13414 7041
rect 13358 6967 13414 6976
rect 13372 4758 13400 6967
rect 13464 4826 13492 8230
rect 13556 7342 13584 13246
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13556 6254 13584 6598
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13542 5944 13598 5953
rect 13542 5879 13544 5888
rect 13596 5879 13598 5888
rect 13544 5850 13596 5856
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13360 4752 13412 4758
rect 13360 4694 13412 4700
rect 13556 4264 13584 5510
rect 13648 4826 13676 18090
rect 13832 18086 13860 18142
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13740 16794 13768 17070
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13832 16658 13860 17206
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13740 12102 13768 14282
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 12753 13860 13806
rect 13818 12744 13874 12753
rect 13818 12679 13874 12688
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13832 11898 13860 12242
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13740 10713 13768 11562
rect 13832 11150 13860 11834
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13726 10704 13782 10713
rect 13726 10639 13782 10648
rect 13726 10296 13782 10305
rect 13726 10231 13782 10240
rect 13820 10260 13872 10266
rect 13740 8922 13768 10231
rect 13820 10202 13872 10208
rect 13832 9081 13860 10202
rect 13818 9072 13874 9081
rect 13818 9007 13874 9016
rect 13740 8894 13860 8922
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13740 7954 13768 8774
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13832 7800 13860 8894
rect 13740 7772 13860 7800
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13464 4236 13584 4264
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13464 2310 13492 4236
rect 13542 4176 13598 4185
rect 13740 4146 13768 7772
rect 13820 6112 13872 6118
rect 13818 6080 13820 6089
rect 13872 6080 13874 6089
rect 13818 6015 13874 6024
rect 13818 5944 13874 5953
rect 13818 5879 13874 5888
rect 13542 4111 13598 4120
rect 13728 4140 13780 4146
rect 13556 2582 13584 4111
rect 13728 4082 13780 4088
rect 13740 3602 13768 4082
rect 13832 3670 13860 5879
rect 13924 3942 13952 18022
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14016 15978 14044 17070
rect 14108 16046 14136 17070
rect 14188 17060 14240 17066
rect 14188 17002 14240 17008
rect 14200 16726 14228 17002
rect 14188 16720 14240 16726
rect 14188 16662 14240 16668
rect 14186 16552 14242 16561
rect 14186 16487 14242 16496
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 14016 15706 14044 15914
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 14108 15094 14136 15982
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14016 14074 14044 14554
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14108 14385 14136 14418
rect 14094 14376 14150 14385
rect 14094 14311 14150 14320
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 14016 12442 14044 13262
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14108 12646 14136 12922
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14004 11280 14056 11286
rect 14004 11222 14056 11228
rect 14016 10470 14044 11222
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14016 5166 14044 10066
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 14016 3738 14044 5102
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13818 3224 13874 3233
rect 13818 3159 13874 3168
rect 13832 2650 13860 3159
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13544 2576 13596 2582
rect 13544 2518 13596 2524
rect 13728 2372 13780 2378
rect 13728 2314 13780 2320
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 13740 1834 13768 2314
rect 14016 1902 14044 3674
rect 14108 3516 14136 12038
rect 14200 5370 14228 16487
rect 14292 11626 14320 18142
rect 14384 17746 14412 19858
rect 14476 18834 14504 22520
rect 14936 20346 14964 22520
rect 15200 21208 15252 21214
rect 15200 21150 15252 21156
rect 15212 20602 15240 21150
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 14752 20318 14964 20346
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 14556 19236 14608 19242
rect 14556 19178 14608 19184
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14462 18184 14518 18193
rect 14568 18170 14596 19178
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14660 18290 14688 19110
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14568 18142 14688 18170
rect 14462 18119 14518 18128
rect 14476 18068 14504 18119
rect 14556 18080 14608 18086
rect 14476 18040 14556 18068
rect 14556 18022 14608 18028
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14384 17105 14412 17682
rect 14370 17096 14426 17105
rect 14370 17031 14426 17040
rect 14660 16998 14688 18142
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14462 16552 14518 16561
rect 14462 16487 14518 16496
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14384 15502 14412 15642
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14372 15088 14424 15094
rect 14372 15030 14424 15036
rect 14384 14618 14412 15030
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14292 8838 14320 10610
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14292 8090 14320 8230
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14292 6934 14320 7346
rect 14280 6928 14332 6934
rect 14280 6870 14332 6876
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14292 5030 14320 6598
rect 14384 5710 14412 14350
rect 14476 12918 14504 16487
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14568 14414 14596 15846
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 14554 13424 14610 13433
rect 14554 13359 14610 13368
rect 14464 12912 14516 12918
rect 14464 12854 14516 12860
rect 14568 12850 14596 13359
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14568 12102 14596 12786
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14476 10674 14504 11494
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14462 10568 14518 10577
rect 14462 10503 14464 10512
rect 14516 10503 14518 10512
rect 14464 10474 14516 10480
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14476 8430 14504 9454
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14476 7410 14504 8366
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14568 7256 14596 11562
rect 14476 7228 14596 7256
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14384 5234 14412 5646
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14200 4758 14228 4966
rect 14188 4752 14240 4758
rect 14292 4729 14320 4966
rect 14188 4694 14240 4700
rect 14278 4720 14334 4729
rect 14278 4655 14334 4664
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14292 4214 14320 4422
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14188 3528 14240 3534
rect 14108 3488 14188 3516
rect 14188 3470 14240 3476
rect 14292 2990 14320 4150
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 14200 2650 14228 2858
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 14292 2038 14320 2382
rect 14384 2038 14412 3606
rect 14476 3040 14504 7228
rect 14660 7154 14688 16934
rect 14752 16776 14780 20318
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 15212 19394 15240 20334
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 15304 19825 15332 19858
rect 15290 19816 15346 19825
rect 15290 19751 15346 19760
rect 15212 19366 15332 19394
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 15212 17814 15240 18906
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15028 17202 15056 17614
rect 15212 17542 15240 17614
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 14752 16748 14872 16776
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14568 7126 14688 7154
rect 14568 4622 14596 7126
rect 14646 7032 14702 7041
rect 14646 6967 14702 6976
rect 14660 6458 14688 6967
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14646 5944 14702 5953
rect 14646 5879 14648 5888
rect 14700 5879 14702 5888
rect 14648 5850 14700 5856
rect 14646 5400 14702 5409
rect 14646 5335 14702 5344
rect 14660 4826 14688 5335
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14568 4214 14596 4558
rect 14556 4208 14608 4214
rect 14556 4150 14608 4156
rect 14752 4078 14780 16594
rect 14844 16522 14872 16748
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 15212 15910 15240 17478
rect 15304 16590 15332 19366
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15304 15706 15332 16526
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14844 12102 14872 12242
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14844 11937 14872 12038
rect 14830 11928 14886 11937
rect 14830 11863 14886 11872
rect 15014 11928 15070 11937
rect 15014 11863 15070 11872
rect 15028 11694 15056 11863
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15212 11218 15240 13126
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15304 11234 15332 12650
rect 15396 11393 15424 22520
rect 15476 19236 15528 19242
rect 15528 19196 15608 19224
rect 15476 19178 15528 19184
rect 15580 18834 15608 19196
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15382 11384 15438 11393
rect 15382 11319 15438 11328
rect 15200 11212 15252 11218
rect 15304 11206 15424 11234
rect 15200 11154 15252 11160
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 14830 10704 14886 10713
rect 14830 10639 14832 10648
rect 14884 10639 14886 10648
rect 14832 10610 14884 10616
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15106 10024 15162 10033
rect 15106 9959 15162 9968
rect 15120 9489 15148 9959
rect 15304 9518 15332 11018
rect 15396 11014 15424 11206
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 15382 10840 15438 10849
rect 15382 10775 15438 10784
rect 15292 9512 15344 9518
rect 15106 9480 15162 9489
rect 15396 9489 15424 10775
rect 15292 9454 15344 9460
rect 15382 9480 15438 9489
rect 15106 9415 15162 9424
rect 15200 9444 15252 9450
rect 15382 9415 15438 9424
rect 15200 9386 15252 9392
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 14924 7336 14976 7342
rect 14922 7304 14924 7313
rect 14976 7304 14978 7313
rect 14922 7239 14978 7248
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 15212 6730 15240 9386
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15304 8634 15332 8978
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15304 7546 15332 8298
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 15212 6322 15240 6666
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 15212 5710 15240 6258
rect 15304 5914 15332 7142
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15290 5264 15346 5273
rect 15290 5199 15346 5208
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 15212 3777 15240 4218
rect 15304 4185 15332 5199
rect 15396 4690 15424 9318
rect 15488 4826 15516 18770
rect 15580 16658 15608 18770
rect 15660 18420 15712 18426
rect 15660 18362 15712 18368
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15580 16114 15608 16594
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15580 14550 15608 15506
rect 15568 14544 15620 14550
rect 15568 14486 15620 14492
rect 15580 14074 15608 14486
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15580 10849 15608 13874
rect 15566 10840 15622 10849
rect 15566 10775 15622 10784
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15580 10441 15608 10474
rect 15566 10432 15622 10441
rect 15566 10367 15622 10376
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15580 8922 15608 10134
rect 15672 9178 15700 18362
rect 15750 18184 15806 18193
rect 15750 18119 15806 18128
rect 15764 17105 15792 18119
rect 15856 17490 15884 22520
rect 16316 20890 16344 22520
rect 16040 20862 16344 20890
rect 15936 17808 15988 17814
rect 15934 17776 15936 17785
rect 15988 17776 15990 17785
rect 15934 17711 15990 17720
rect 15856 17462 15976 17490
rect 15750 17096 15806 17105
rect 15750 17031 15806 17040
rect 15948 16998 15976 17462
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15764 14482 15792 16050
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15764 13433 15792 14418
rect 15750 13424 15806 13433
rect 15750 13359 15806 13368
rect 15764 12850 15792 13359
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15856 12374 15884 16458
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 15948 12481 15976 15846
rect 16040 13938 16068 20862
rect 16776 20346 16804 22520
rect 17236 20618 17264 22520
rect 16592 20318 16804 20346
rect 16868 20590 17264 20618
rect 16592 19242 16620 20318
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16684 20058 16712 20198
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16580 19236 16632 19242
rect 16580 19178 16632 19184
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16316 17241 16344 19110
rect 16684 17626 16712 19314
rect 16762 18184 16818 18193
rect 16762 18119 16818 18128
rect 16592 17598 16712 17626
rect 16302 17232 16358 17241
rect 16302 17167 16358 17176
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16132 14074 16160 14214
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 15934 12472 15990 12481
rect 15934 12407 15990 12416
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 15752 12232 15804 12238
rect 16132 12209 16160 12242
rect 15752 12174 15804 12180
rect 16118 12200 16174 12209
rect 15764 11132 15792 12174
rect 16118 12135 16174 12144
rect 15844 12096 15896 12102
rect 16120 12096 16172 12102
rect 15896 12056 15976 12084
rect 15844 12038 15896 12044
rect 15844 11144 15896 11150
rect 15764 11104 15844 11132
rect 15844 11086 15896 11092
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15764 10577 15792 10678
rect 15750 10568 15806 10577
rect 15750 10503 15806 10512
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 10198 15792 10406
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15764 9330 15792 9998
rect 15856 9450 15884 11086
rect 15948 9586 15976 12056
rect 16026 12064 16082 12073
rect 16120 12038 16172 12044
rect 16026 11999 16082 12008
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 15764 9302 15884 9330
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15856 8974 15884 9302
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 15844 8968 15896 8974
rect 15580 8894 15792 8922
rect 15844 8910 15896 8916
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15672 8634 15700 8774
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 15580 8022 15608 8502
rect 15658 8392 15714 8401
rect 15658 8327 15714 8336
rect 15568 8016 15620 8022
rect 15568 7958 15620 7964
rect 15672 7834 15700 8327
rect 15580 7806 15700 7834
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15290 4176 15346 4185
rect 15290 4111 15346 4120
rect 15580 3942 15608 7806
rect 15764 6361 15792 8894
rect 15856 7954 15884 8910
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15856 6866 15884 7890
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15842 6624 15898 6633
rect 15842 6559 15898 6568
rect 15856 6458 15884 6559
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15750 6352 15806 6361
rect 15750 6287 15806 6296
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15672 5273 15700 5714
rect 15658 5264 15714 5273
rect 15658 5199 15714 5208
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15198 3768 15254 3777
rect 15198 3703 15254 3712
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 14660 3058 14688 3538
rect 15764 3233 15792 6190
rect 15948 6186 15976 9046
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 16040 3942 16068 11999
rect 16132 10266 16160 12038
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16132 8498 16160 9318
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16118 8392 16174 8401
rect 16118 8327 16174 8336
rect 16132 4078 16160 8327
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 16118 3904 16174 3913
rect 16118 3839 16174 3848
rect 16132 3670 16160 3839
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 15750 3224 15806 3233
rect 15750 3159 15806 3168
rect 14556 3052 14608 3058
rect 14476 3012 14556 3040
rect 14556 2994 14608 3000
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14660 2446 14688 2994
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 15488 2689 15516 2926
rect 15474 2680 15530 2689
rect 15474 2615 15530 2624
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 16224 2378 16252 16934
rect 16316 15162 16344 16934
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 16408 15366 16436 15914
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16408 15042 16436 15302
rect 16316 15014 16436 15042
rect 16316 4214 16344 15014
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16408 13530 16436 13670
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16500 13410 16528 16662
rect 16592 14929 16620 17598
rect 16578 14920 16634 14929
rect 16578 14855 16634 14864
rect 16776 14600 16804 18119
rect 16408 13382 16528 13410
rect 16592 14572 16804 14600
rect 16408 7970 16436 13382
rect 16592 11778 16620 14572
rect 16868 14498 16896 20590
rect 17132 20460 17184 20466
rect 17316 20460 17368 20466
rect 17132 20402 17184 20408
rect 17236 20420 17316 20448
rect 17040 20324 17092 20330
rect 17040 20266 17092 20272
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 16960 18834 16988 19450
rect 17052 18970 17080 20266
rect 17144 19961 17172 20402
rect 17130 19952 17186 19961
rect 17130 19887 17186 19896
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16960 18290 16988 18770
rect 17144 18426 17172 19790
rect 17236 19514 17264 20420
rect 17316 20402 17368 20408
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17328 18970 17356 19790
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 17590 18184 17646 18193
rect 17590 18119 17646 18128
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16960 15065 16988 18022
rect 17604 17814 17632 18119
rect 17696 18057 17724 22520
rect 17880 20602 17908 22607
rect 18142 22522 18198 23000
rect 18142 22520 18276 22522
rect 18602 22520 18658 23000
rect 19062 22520 19118 23000
rect 19522 22520 19578 23000
rect 19982 22520 20038 23000
rect 20442 22520 20498 23000
rect 20902 22520 20958 23000
rect 21362 22520 21418 23000
rect 21822 22520 21878 23000
rect 22282 22520 22338 23000
rect 22742 22520 22798 23000
rect 18156 22494 18276 22520
rect 17958 22128 18014 22137
rect 17958 22063 18014 22072
rect 17972 21214 18000 22063
rect 17960 21208 18012 21214
rect 17960 21150 18012 21156
rect 18050 21176 18106 21185
rect 18050 21111 18106 21120
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17868 20596 17920 20602
rect 17868 20538 17920 20544
rect 17972 19446 18000 20946
rect 18064 20806 18092 21111
rect 18248 21010 18276 22494
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17972 18290 18000 18770
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17776 18148 17828 18154
rect 17776 18090 17828 18096
rect 17682 18048 17738 18057
rect 17682 17983 17738 17992
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17222 17368 17278 17377
rect 17222 17303 17278 17312
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17144 15910 17172 16594
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 16946 15056 17002 15065
rect 16946 14991 17002 15000
rect 16948 14884 17000 14890
rect 16948 14826 17000 14832
rect 16500 11750 16620 11778
rect 16684 14470 16896 14498
rect 16500 11626 16528 11750
rect 16684 11744 16712 14470
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16776 11898 16804 13670
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16684 11716 16804 11744
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16500 11354 16528 11562
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16500 9722 16528 10474
rect 16592 10198 16620 11630
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16684 11286 16712 11494
rect 16672 11280 16724 11286
rect 16672 11222 16724 11228
rect 16670 11112 16726 11121
rect 16670 11047 16726 11056
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16592 9722 16620 10134
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 16500 8537 16528 9046
rect 16486 8528 16542 8537
rect 16486 8463 16542 8472
rect 16408 7942 16528 7970
rect 16394 7440 16450 7449
rect 16394 7375 16450 7384
rect 16408 7342 16436 7375
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16408 5137 16436 7278
rect 16394 5128 16450 5137
rect 16394 5063 16450 5072
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16408 4593 16436 4626
rect 16394 4584 16450 4593
rect 16394 4519 16450 4528
rect 16304 4208 16356 4214
rect 16304 4150 16356 4156
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16316 3194 16344 4014
rect 16396 3936 16448 3942
rect 16500 3913 16528 7942
rect 16592 7410 16620 9658
rect 16684 7954 16712 11047
rect 16776 9625 16804 11716
rect 16762 9616 16818 9625
rect 16762 9551 16818 9560
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16776 7834 16804 9318
rect 16684 7806 16804 7834
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16578 7304 16634 7313
rect 16578 7239 16580 7248
rect 16632 7239 16634 7248
rect 16580 7210 16632 7216
rect 16684 7154 16712 7806
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16592 7126 16712 7154
rect 16396 3878 16448 3884
rect 16486 3904 16542 3913
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16408 2650 16436 3878
rect 16486 3839 16542 3848
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16500 3194 16528 3470
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16592 2854 16620 7126
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16684 5234 16712 6938
rect 16776 6934 16804 7686
rect 16868 7546 16896 13806
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16960 7392 16988 14826
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 17052 12986 17080 14418
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17052 11694 17080 12038
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17052 11393 17080 11494
rect 17038 11384 17094 11393
rect 17038 11319 17094 11328
rect 17144 11200 17172 15846
rect 17236 12374 17264 17303
rect 17696 16726 17724 17478
rect 17684 16720 17736 16726
rect 17684 16662 17736 16668
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17224 12368 17276 12374
rect 17224 12310 17276 12316
rect 16868 7364 16988 7392
rect 17052 11172 17172 11200
rect 16764 6928 16816 6934
rect 16764 6870 16816 6876
rect 16868 6254 16896 7364
rect 16946 7304 17002 7313
rect 16946 7239 17002 7248
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16776 5914 16804 6054
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16868 5370 16896 6054
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16868 4826 16896 4966
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16854 4720 16910 4729
rect 16684 4434 16712 4694
rect 16854 4655 16856 4664
rect 16908 4655 16910 4664
rect 16856 4626 16908 4632
rect 16684 4406 16804 4434
rect 16776 4162 16804 4406
rect 16868 4282 16896 4626
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16776 4134 16896 4162
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16776 3738 16804 3878
rect 16868 3738 16896 4134
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 16670 3632 16726 3641
rect 16670 3567 16726 3576
rect 16684 3194 16712 3567
rect 16762 3224 16818 3233
rect 16672 3188 16724 3194
rect 16762 3159 16818 3168
rect 16672 3130 16724 3136
rect 16776 2990 16804 3159
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16960 2922 16988 7239
rect 17052 4214 17080 11172
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17144 10470 17172 11018
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17144 10130 17172 10406
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17236 8430 17264 12310
rect 17328 9382 17356 14758
rect 17696 14346 17724 15506
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17696 14090 17724 14282
rect 17604 14062 17724 14090
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17144 7313 17172 8230
rect 17222 7848 17278 7857
rect 17222 7783 17278 7792
rect 17236 7546 17264 7783
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17130 7304 17186 7313
rect 17130 7239 17186 7248
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 17236 5302 17264 6870
rect 17224 5296 17276 5302
rect 17224 5238 17276 5244
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17144 4486 17172 4966
rect 17236 4622 17264 5238
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 17052 3058 17080 4150
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 17144 2650 17172 4218
rect 17328 3670 17356 9114
rect 17420 8090 17448 13330
rect 17512 11286 17540 13874
rect 17500 11280 17552 11286
rect 17500 11222 17552 11228
rect 17512 10266 17540 11222
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17420 7698 17448 7890
rect 17512 7818 17540 10202
rect 17604 9178 17632 14062
rect 17682 13424 17738 13433
rect 17682 13359 17684 13368
rect 17736 13359 17738 13368
rect 17684 13330 17736 13336
rect 17788 12730 17816 18090
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17972 17338 18000 17682
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 18064 17218 18092 19654
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17972 17190 18092 17218
rect 17696 12702 17816 12730
rect 17696 12617 17724 12702
rect 17682 12608 17738 12617
rect 17682 12543 17738 12552
rect 17682 12336 17738 12345
rect 17682 12271 17738 12280
rect 17696 10810 17724 12271
rect 17880 11778 17908 17138
rect 17972 16998 18000 17190
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 18050 16144 18106 16153
rect 18050 16079 18106 16088
rect 18064 15638 18092 16079
rect 18052 15632 18104 15638
rect 18052 15574 18104 15580
rect 17958 15056 18014 15065
rect 17958 14991 18014 15000
rect 17972 14074 18000 14991
rect 18156 14385 18184 19382
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18616 17864 18644 22520
rect 18786 21584 18842 21593
rect 18786 21519 18842 21528
rect 18694 20632 18750 20641
rect 18694 20567 18750 20576
rect 18708 20534 18736 20567
rect 18696 20528 18748 20534
rect 18696 20470 18748 20476
rect 18694 19680 18750 19689
rect 18694 19615 18750 19624
rect 18708 19378 18736 19615
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18800 18630 18828 21519
rect 19076 20346 19104 22520
rect 18892 20318 19104 20346
rect 18892 18873 18920 20318
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 18984 19378 19012 20198
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18878 18864 18934 18873
rect 18878 18799 18934 18808
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18972 18148 19024 18154
rect 18972 18090 19024 18096
rect 18616 17836 18920 17864
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18616 17202 18644 17682
rect 18788 17604 18840 17610
rect 18788 17546 18840 17552
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18142 14376 18198 14385
rect 18142 14311 18198 14320
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18156 13870 18184 14214
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 18050 13696 18106 13705
rect 18050 13631 18106 13640
rect 18064 13462 18092 13631
rect 18052 13456 18104 13462
rect 18156 13433 18184 13806
rect 18052 13398 18104 13404
rect 18142 13424 18198 13433
rect 17960 13388 18012 13394
rect 18142 13359 18198 13368
rect 17960 13330 18012 13336
rect 17972 13274 18000 13330
rect 17972 13246 18092 13274
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17972 11898 18000 13126
rect 18064 12617 18092 13246
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18328 12912 18380 12918
rect 18234 12880 18290 12889
rect 18616 12866 18644 16934
rect 18328 12854 18380 12860
rect 18234 12815 18290 12824
rect 18248 12714 18276 12815
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 18050 12608 18106 12617
rect 18050 12543 18106 12552
rect 18050 12472 18106 12481
rect 18050 12407 18106 12416
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17958 11792 18014 11801
rect 17880 11750 17958 11778
rect 17958 11727 18014 11736
rect 18064 11642 18092 12407
rect 18142 12336 18198 12345
rect 18142 12271 18198 12280
rect 18340 12288 18368 12854
rect 18432 12838 18644 12866
rect 18432 12481 18460 12838
rect 18708 12782 18736 17070
rect 18800 16046 18828 17546
rect 18892 17218 18920 17836
rect 18984 17338 19012 18090
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18892 17190 19012 17218
rect 18878 17096 18934 17105
rect 18878 17031 18934 17040
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18800 15094 18828 15846
rect 18788 15088 18840 15094
rect 18788 15030 18840 15036
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18800 14278 18828 14894
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18786 14104 18842 14113
rect 18786 14039 18842 14048
rect 18800 14006 18828 14039
rect 18788 14000 18840 14006
rect 18788 13942 18840 13948
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18800 12986 18828 13330
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18892 12866 18920 17031
rect 18800 12838 18920 12866
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18418 12472 18474 12481
rect 18418 12407 18474 12416
rect 18524 12306 18552 12582
rect 18512 12300 18564 12306
rect 17972 11614 18092 11642
rect 17774 11520 17830 11529
rect 17774 11455 17830 11464
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17684 9444 17736 9450
rect 17684 9386 17736 9392
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17420 7670 17540 7698
rect 17512 7002 17540 7670
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17498 6896 17554 6905
rect 17498 6831 17554 6840
rect 17512 6186 17540 6831
rect 17604 6730 17632 8978
rect 17696 8838 17724 9386
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 17500 6180 17552 6186
rect 17500 6122 17552 6128
rect 17420 4146 17448 6122
rect 17604 5710 17632 6666
rect 17696 6322 17724 8774
rect 17788 8294 17816 11455
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17880 10985 17908 11222
rect 17866 10976 17922 10985
rect 17866 10911 17922 10920
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17880 8090 17908 9930
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17788 6458 17816 7822
rect 17880 6730 17908 7890
rect 17972 7324 18000 11614
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 10606 18092 11494
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18064 9586 18092 10066
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18064 8566 18092 9522
rect 18052 8560 18104 8566
rect 18052 8502 18104 8508
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 18064 7449 18092 8026
rect 18050 7440 18106 7449
rect 18050 7375 18106 7384
rect 18052 7336 18104 7342
rect 17972 7296 18052 7324
rect 18052 7278 18104 7284
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 18050 7168 18106 7177
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17972 6202 18000 7142
rect 18050 7103 18106 7112
rect 17696 6174 18000 6202
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17604 5234 17632 5646
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17590 5128 17646 5137
rect 17590 5063 17646 5072
rect 17604 4690 17632 5063
rect 17696 4758 17724 6174
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17684 4752 17736 4758
rect 17788 4729 17816 5714
rect 17972 5370 18000 5714
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17684 4694 17736 4700
rect 17774 4720 17830 4729
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17592 4684 17644 4690
rect 17774 4655 17830 4664
rect 17592 4626 17644 4632
rect 17512 4282 17540 4626
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17500 4004 17552 4010
rect 17500 3946 17552 3952
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17316 3664 17368 3670
rect 17316 3606 17368 3612
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17328 2446 17356 3606
rect 17512 3466 17540 3946
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 17788 3641 17816 3674
rect 17774 3632 17830 3641
rect 17774 3567 17830 3576
rect 17500 3460 17552 3466
rect 17500 3402 17552 3408
rect 17880 2582 17908 3946
rect 18064 3602 18092 7103
rect 18156 4758 18184 12271
rect 18340 12260 18460 12288
rect 18432 12186 18460 12260
rect 18616 12288 18644 12650
rect 18800 12345 18828 12838
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18786 12336 18842 12345
rect 18616 12260 18736 12288
rect 18786 12271 18842 12280
rect 18512 12242 18564 12248
rect 18432 12158 18644 12186
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 18248 10169 18276 10678
rect 18234 10160 18290 10169
rect 18234 10095 18290 10104
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18234 9344 18290 9353
rect 18234 9279 18290 9288
rect 18248 9110 18276 9279
rect 18236 9104 18288 9110
rect 18236 9046 18288 9052
rect 18234 8936 18290 8945
rect 18234 8871 18236 8880
rect 18288 8871 18290 8880
rect 18236 8842 18288 8848
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18524 6866 18552 7346
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18144 4752 18196 4758
rect 18144 4694 18196 4700
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18142 3904 18198 3913
rect 18142 3839 18198 3848
rect 18156 3738 18184 3839
rect 18326 3768 18382 3777
rect 18144 3732 18196 3738
rect 18326 3703 18382 3712
rect 18144 3674 18196 3680
rect 18340 3602 18368 3703
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18616 3058 18644 12158
rect 18708 12050 18736 12260
rect 18708 12022 18828 12050
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18708 11354 18736 11834
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18708 10198 18736 11290
rect 18696 10192 18748 10198
rect 18696 10134 18748 10140
rect 18800 10044 18828 12022
rect 18708 10016 18828 10044
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 16212 2372 16264 2378
rect 16212 2314 16264 2320
rect 14280 2032 14332 2038
rect 14280 1974 14332 1980
rect 14372 2032 14424 2038
rect 14372 1974 14424 1980
rect 14004 1896 14056 1902
rect 14004 1838 14056 1844
rect 13728 1828 13780 1834
rect 13728 1770 13780 1776
rect 18064 1766 18092 2450
rect 18708 2310 18736 10016
rect 18786 8664 18842 8673
rect 18892 8634 18920 12718
rect 18786 8599 18842 8608
rect 18880 8628 18932 8634
rect 18800 6254 18828 8599
rect 18880 8570 18932 8576
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 18892 7478 18920 7890
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 18880 7336 18932 7342
rect 18878 7304 18880 7313
rect 18932 7304 18934 7313
rect 18878 7239 18934 7248
rect 18880 6928 18932 6934
rect 18880 6870 18932 6876
rect 18892 6322 18920 6870
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 18788 6248 18840 6254
rect 18788 6190 18840 6196
rect 18878 6216 18934 6225
rect 18878 6151 18880 6160
rect 18932 6151 18934 6160
rect 18880 6122 18932 6128
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 18800 4826 18828 6054
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18892 5302 18920 5646
rect 18984 5574 19012 17190
rect 19076 14385 19104 20198
rect 19154 20088 19210 20097
rect 19154 20023 19210 20032
rect 19168 17728 19196 20023
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 19260 19310 19288 19654
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19168 17700 19380 17728
rect 19246 17640 19302 17649
rect 19246 17575 19302 17584
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 19168 16794 19196 17478
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 19156 16584 19208 16590
rect 19156 16526 19208 16532
rect 19168 15910 19196 16526
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 19168 14958 19196 15846
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19062 14376 19118 14385
rect 19260 14362 19288 17575
rect 19352 15978 19380 17700
rect 19536 16114 19564 22520
rect 19996 20618 20024 22520
rect 19628 20590 20024 20618
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19628 15994 19656 20590
rect 19892 20460 19944 20466
rect 19892 20402 19944 20408
rect 19904 19854 19932 20402
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19800 19236 19852 19242
rect 19800 19178 19852 19184
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19444 15966 19656 15994
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19352 14618 19380 15506
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19062 14311 19118 14320
rect 19168 14334 19288 14362
rect 19168 12782 19196 14334
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18878 4584 18934 4593
rect 18788 4548 18840 4554
rect 18878 4519 18934 4528
rect 18788 4490 18840 4496
rect 18800 4146 18828 4490
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18892 3534 18920 4519
rect 19076 4026 19104 12378
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19168 9178 19196 11494
rect 19260 11218 19288 14214
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19352 12918 19380 13126
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19248 10600 19300 10606
rect 19248 10542 19300 10548
rect 19260 10130 19288 10542
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19168 7410 19196 8434
rect 19246 7712 19302 7721
rect 19246 7647 19302 7656
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19260 7290 19288 7647
rect 19168 7262 19288 7290
rect 19168 6769 19196 7262
rect 19154 6760 19210 6769
rect 19154 6695 19210 6704
rect 19168 6118 19196 6695
rect 19246 6624 19302 6633
rect 19246 6559 19302 6568
rect 19156 6112 19208 6118
rect 19156 6054 19208 6060
rect 19260 5914 19288 6559
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19156 5840 19208 5846
rect 19156 5782 19208 5788
rect 19246 5808 19302 5817
rect 19168 5681 19196 5782
rect 19246 5743 19302 5752
rect 19154 5672 19210 5681
rect 19154 5607 19210 5616
rect 19076 3998 19196 4026
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 19076 2922 19104 3878
rect 19168 3670 19196 3998
rect 19156 3664 19208 3670
rect 19156 3606 19208 3612
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19168 2990 19196 3334
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 19064 2916 19116 2922
rect 19064 2858 19116 2864
rect 19260 2854 19288 5743
rect 19352 4826 19380 12310
rect 19444 11354 19472 15966
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19628 14618 19656 15302
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19524 13796 19576 13802
rect 19524 13738 19576 13744
rect 19536 12646 19564 13738
rect 19616 13184 19668 13190
rect 19616 13126 19668 13132
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19628 12458 19656 13126
rect 19536 12430 19656 12458
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19444 4690 19472 11086
rect 19536 4758 19564 12430
rect 19720 11898 19748 14350
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19708 11348 19760 11354
rect 19708 11290 19760 11296
rect 19614 10704 19670 10713
rect 19614 10639 19670 10648
rect 19628 9178 19656 10639
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19720 9110 19748 11290
rect 19708 9104 19760 9110
rect 19708 9046 19760 9052
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19616 8900 19668 8906
rect 19616 8842 19668 8848
rect 19628 5658 19656 8842
rect 19720 8090 19748 8910
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 19628 5630 19748 5658
rect 19524 4752 19576 4758
rect 19524 4694 19576 4700
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19524 4616 19576 4622
rect 19524 4558 19576 4564
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19352 3534 19380 4014
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 19430 2544 19486 2553
rect 19430 2479 19432 2488
rect 19484 2479 19486 2488
rect 19432 2450 19484 2456
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18694 2136 18750 2145
rect 18694 2071 18750 2080
rect 18512 2032 18564 2038
rect 18512 1974 18564 1980
rect 18052 1760 18104 1766
rect 18524 1737 18552 1974
rect 18708 1902 18736 2071
rect 18696 1896 18748 1902
rect 18696 1838 18748 1844
rect 19536 1834 19564 4558
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19628 3738 19656 4422
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 19720 2990 19748 5630
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 19812 2650 19840 19178
rect 19904 18630 19932 19790
rect 20456 19394 20484 22520
rect 20168 19372 20220 19378
rect 20456 19366 20668 19394
rect 20168 19314 20220 19320
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19904 18222 19932 18566
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 20088 14521 20116 19246
rect 20180 18086 20208 19314
rect 20640 19292 20668 19366
rect 20640 19264 20852 19292
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20732 18601 20760 19110
rect 20718 18592 20774 18601
rect 20718 18527 20774 18536
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20180 17134 20208 18022
rect 20824 17678 20852 19264
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20444 17604 20496 17610
rect 20444 17546 20496 17552
rect 20456 17338 20484 17546
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 20548 16266 20576 17614
rect 20812 17536 20864 17542
rect 20812 17478 20864 17484
rect 20456 16238 20576 16266
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20272 14822 20300 15438
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20074 14512 20130 14521
rect 20074 14447 20130 14456
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20180 13734 20208 14350
rect 20272 13870 20300 14758
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19996 12102 20024 12650
rect 20074 12608 20130 12617
rect 20074 12543 20130 12552
rect 20088 12442 20116 12543
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19996 11762 20024 12038
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 20076 11552 20128 11558
rect 19996 11512 20076 11540
rect 19996 11286 20024 11512
rect 20076 11494 20128 11500
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 19892 10532 19944 10538
rect 19892 10474 19944 10480
rect 19904 9926 19932 10474
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19904 7886 19932 9862
rect 19996 9722 20024 11222
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19904 7206 19932 7686
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 19904 4049 19932 6190
rect 19890 4040 19946 4049
rect 19890 3975 19946 3984
rect 19996 3602 20024 9386
rect 20088 8974 20116 10746
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 20088 6254 20116 8774
rect 20180 8430 20208 13670
rect 20272 11762 20300 13806
rect 20350 12200 20406 12209
rect 20350 12135 20406 12144
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20364 11626 20392 12135
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20272 9738 20300 11086
rect 20456 9908 20484 16238
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20548 10033 20576 16050
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20640 10810 20668 12242
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20534 10024 20590 10033
rect 20534 9959 20590 9968
rect 20456 9880 20668 9908
rect 20534 9752 20590 9761
rect 20272 9710 20392 9738
rect 20260 9512 20312 9518
rect 20260 9454 20312 9460
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20168 8288 20220 8294
rect 20168 8230 20220 8236
rect 20076 6248 20128 6254
rect 20076 6190 20128 6196
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 20088 5234 20116 6054
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 20180 3194 20208 8230
rect 20272 5370 20300 9454
rect 20364 8294 20392 9710
rect 20444 9716 20496 9722
rect 20534 9687 20590 9696
rect 20444 9658 20496 9664
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20352 8016 20404 8022
rect 20352 7958 20404 7964
rect 20364 7546 20392 7958
rect 20456 7818 20484 9658
rect 20548 8430 20576 9687
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20640 8294 20668 9880
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20536 8288 20588 8294
rect 20536 8230 20588 8236
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20364 5302 20392 7482
rect 20444 7472 20496 7478
rect 20444 7414 20496 7420
rect 20352 5296 20404 5302
rect 20352 5238 20404 5244
rect 20260 4752 20312 4758
rect 20260 4694 20312 4700
rect 20272 4146 20300 4694
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20272 3534 20300 4082
rect 20456 4078 20484 7414
rect 20548 7342 20576 8230
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 20548 6322 20576 7278
rect 20640 7177 20668 7890
rect 20626 7168 20682 7177
rect 20626 7103 20682 7112
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20548 3233 20576 6054
rect 20732 4622 20760 9658
rect 20824 7750 20852 17478
rect 20916 17338 20944 22520
rect 21376 17490 21404 22520
rect 21836 17542 21864 22520
rect 21008 17462 21404 17490
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20916 8514 20944 17138
rect 21008 8786 21036 17462
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21088 10532 21140 10538
rect 21088 10474 21140 10480
rect 21100 9722 21128 10474
rect 21192 9722 21220 17274
rect 22296 17202 22324 22520
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22756 10538 22784 22520
rect 22744 10532 22796 10538
rect 22744 10474 22796 10480
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21008 8758 21220 8786
rect 20916 8486 21036 8514
rect 20904 8424 20956 8430
rect 20904 8366 20956 8372
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20916 7478 20944 8366
rect 20904 7472 20956 7478
rect 20904 7414 20956 7420
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 21008 3505 21036 8486
rect 20994 3496 21050 3505
rect 20720 3460 20772 3466
rect 20994 3431 21050 3440
rect 20720 3402 20772 3408
rect 20534 3224 20590 3233
rect 20168 3188 20220 3194
rect 20534 3159 20590 3168
rect 20168 3130 20220 3136
rect 19800 2644 19852 2650
rect 19800 2586 19852 2592
rect 19524 1828 19576 1834
rect 19524 1770 19576 1776
rect 18052 1702 18104 1708
rect 18510 1728 18566 1737
rect 18510 1663 18566 1672
rect 16120 1624 16172 1630
rect 16120 1566 16172 1572
rect 13084 1352 13136 1358
rect 13084 1294 13136 1300
rect 12070 1184 12126 1193
rect 12070 1119 12126 1128
rect 16132 480 16160 1566
rect 18144 1352 18196 1358
rect 18144 1294 18196 1300
rect 18156 649 18184 1294
rect 18142 640 18198 649
rect 18142 575 18198 584
rect 20732 480 20760 3402
rect 21192 3097 21220 8758
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21178 3088 21234 3097
rect 21178 3023 21234 3032
rect 21284 2961 21312 7686
rect 21376 4282 21404 9658
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21270 2952 21326 2961
rect 21270 2887 21326 2896
rect 21468 1698 21496 8230
rect 22374 5128 22430 5137
rect 22374 5063 22430 5072
rect 22388 5001 22416 5063
rect 22374 4992 22430 5001
rect 22374 4927 22430 4936
rect 21456 1692 21508 1698
rect 21456 1634 21508 1640
rect 11886 232 11942 241
rect 11886 167 11942 176
rect 16118 0 16174 480
rect 20718 0 20774 480
<< via2 >>
rect 3698 22616 3754 22672
rect 18 18808 74 18864
rect 1398 18964 1454 19000
rect 1398 18944 1400 18964
rect 1400 18944 1452 18964
rect 1452 18944 1454 18964
rect 1950 20576 2006 20632
rect 1398 18536 1454 18592
rect 1214 16904 1270 16960
rect 1122 13232 1178 13288
rect 662 11872 718 11928
rect 1214 11600 1270 11656
rect 1030 10648 1086 10704
rect 570 10104 626 10160
rect 1766 17040 1822 17096
rect 1674 16088 1730 16144
rect 2042 17176 2098 17232
rect 1858 12416 1914 12472
rect 2962 21120 3018 21176
rect 2226 12416 2282 12472
rect 2226 11736 2282 11792
rect 2226 9424 2282 9480
rect 1766 2760 1822 2816
rect 2686 16496 2742 16552
rect 3514 22072 3570 22128
rect 3514 21528 3570 21584
rect 17866 22616 17922 22672
rect 3514 18264 3570 18320
rect 3146 18128 3202 18184
rect 2962 15000 3018 15056
rect 2410 6296 2466 6352
rect 3238 17584 3294 17640
rect 3054 12280 3110 12336
rect 2870 10104 2926 10160
rect 2778 9424 2834 9480
rect 3606 16632 3662 16688
rect 3514 14592 3570 14648
rect 3514 11600 3570 11656
rect 3054 5616 3110 5672
rect 2870 5208 2926 5264
rect 2870 4664 2926 4720
rect 3054 2896 3110 2952
rect 2778 2080 2834 2136
rect 2594 1128 2650 1184
rect 3974 20032 4030 20088
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4250 19624 4306 19680
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4066 18672 4122 18728
rect 4802 18808 4858 18864
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4066 15544 4122 15600
rect 4066 15136 4122 15192
rect 3974 14048 4030 14104
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 3974 13640 4030 13696
rect 3790 13096 3846 13152
rect 3698 12280 3754 12336
rect 3698 10648 3754 10704
rect 3698 10548 3700 10568
rect 3700 10548 3752 10568
rect 3752 10548 3754 10568
rect 3698 10512 3754 10548
rect 3698 10240 3754 10296
rect 3698 9560 3754 9616
rect 3882 12552 3938 12608
rect 3422 2624 3478 2680
rect 3790 6160 3846 6216
rect 3790 5072 3846 5128
rect 3974 9424 4030 9480
rect 4066 9288 4122 9344
rect 3974 8608 4030 8664
rect 4066 8064 4122 8120
rect 4066 7112 4122 7168
rect 4066 6568 4122 6624
rect 3974 4120 4030 4176
rect 3974 3576 4030 3632
rect 4250 11600 4306 11656
rect 4158 5108 4160 5128
rect 4160 5108 4212 5128
rect 4212 5108 4214 5128
rect 4158 5072 4214 5108
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4986 14864 5042 14920
rect 4894 14456 4950 14512
rect 4894 13776 4950 13832
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4710 11212 4766 11248
rect 4710 11192 4712 11212
rect 4712 11192 4764 11212
rect 4764 11192 4766 11212
rect 4526 11056 4582 11112
rect 4710 11076 4766 11112
rect 4710 11056 4712 11076
rect 4712 11056 4764 11076
rect 4764 11056 4766 11076
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4526 9988 4582 10024
rect 4526 9968 4528 9988
rect 4528 9968 4580 9988
rect 4580 9968 4582 9988
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 5078 12552 5134 12608
rect 5814 19216 5870 19272
rect 5354 16668 5356 16688
rect 5356 16668 5408 16688
rect 5408 16668 5410 16688
rect 5354 16632 5410 16668
rect 5354 14184 5410 14240
rect 5262 12416 5318 12472
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4710 7384 4766 7440
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4158 3984 4214 4040
rect 4250 3460 4306 3496
rect 4250 3440 4252 3460
rect 4252 3440 4304 3460
rect 4304 3440 4306 3460
rect 5446 12416 5502 12472
rect 5722 14864 5778 14920
rect 5722 10668 5778 10704
rect 5722 10648 5724 10668
rect 5724 10648 5776 10668
rect 5776 10648 5778 10668
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 3698 3168 3754 3224
rect 5446 5208 5502 5264
rect 6642 18536 6698 18592
rect 6458 12416 6514 12472
rect 6366 11872 6422 11928
rect 6734 18128 6790 18184
rect 7194 18944 7250 19000
rect 6918 17448 6974 17504
rect 6826 12416 6882 12472
rect 8298 20304 8354 20360
rect 8482 20204 8484 20224
rect 8484 20204 8536 20224
rect 8536 20204 8538 20224
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 8482 20168 8538 20204
rect 8482 19896 8538 19952
rect 8390 19760 8446 19816
rect 8206 19252 8208 19272
rect 8208 19252 8260 19272
rect 8260 19252 8262 19272
rect 8206 19216 8262 19252
rect 8482 19236 8538 19272
rect 8482 19216 8484 19236
rect 8484 19216 8536 19236
rect 8536 19216 8538 19236
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 8298 19080 8354 19136
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 8850 20168 8906 20224
rect 8574 18536 8630 18592
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 8206 16632 8262 16688
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7746 15136 7802 15192
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7194 8744 7250 8800
rect 6642 7792 6698 7848
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 4066 1672 4122 1728
rect 7194 7248 7250 7304
rect 7470 6704 7526 6760
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 7746 8608 7802 8664
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7838 7404 7894 7440
rect 7838 7384 7840 7404
rect 7840 7384 7892 7404
rect 7892 7384 7894 7404
rect 8758 18128 8814 18184
rect 9218 18148 9274 18184
rect 9218 18128 9220 18148
rect 9220 18128 9272 18148
rect 9272 18128 9274 18148
rect 8758 11736 8814 11792
rect 8390 9696 8446 9752
rect 8482 9560 8538 9616
rect 8206 7248 8262 7304
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 8574 8916 8576 8936
rect 8576 8916 8628 8936
rect 8628 8916 8630 8936
rect 8574 8880 8630 8916
rect 8114 6840 8170 6896
rect 8390 6860 8446 6896
rect 8390 6840 8392 6860
rect 8392 6840 8444 6860
rect 8444 6840 8446 6860
rect 8390 6704 8446 6760
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 8758 8356 8814 8392
rect 8758 8336 8760 8356
rect 8760 8336 8812 8356
rect 8812 8336 8814 8356
rect 8666 5616 8722 5672
rect 8298 4664 8354 4720
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 8206 3576 8262 3632
rect 7562 2760 7618 2816
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 9310 16904 9366 16960
rect 9126 11736 9182 11792
rect 9678 15700 9734 15736
rect 9678 15680 9680 15700
rect 9680 15680 9732 15700
rect 9732 15680 9734 15700
rect 9586 13776 9642 13832
rect 9494 13232 9550 13288
rect 10966 20204 10968 20224
rect 10968 20204 11020 20224
rect 11020 20204 11022 20224
rect 10966 20168 11022 20204
rect 10506 18672 10562 18728
rect 9586 11600 9642 11656
rect 9126 5516 9128 5536
rect 9128 5516 9180 5536
rect 9180 5516 9182 5536
rect 9126 5480 9182 5516
rect 9310 6296 9366 6352
rect 9586 11328 9642 11384
rect 10414 13912 10470 13968
rect 9770 11192 9826 11248
rect 9678 7248 9734 7304
rect 10230 11056 10286 11112
rect 10414 11736 10470 11792
rect 10506 11600 10562 11656
rect 9770 7112 9826 7168
rect 9586 6996 9642 7032
rect 9586 6976 9588 6996
rect 9588 6976 9640 6996
rect 9640 6976 9642 6996
rect 9586 6024 9642 6080
rect 9954 5888 10010 5944
rect 9770 4800 9826 4856
rect 9678 4256 9734 4312
rect 10230 8472 10286 8528
rect 10046 4120 10102 4176
rect 10046 3732 10102 3768
rect 10046 3712 10048 3732
rect 10048 3712 10100 3732
rect 10100 3712 10102 3732
rect 9586 3032 9642 3088
rect 10230 5208 10286 5264
rect 10414 5072 10470 5128
rect 10322 4936 10378 4992
rect 10322 4528 10378 4584
rect 10874 17584 10930 17640
rect 10966 17448 11022 17504
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 12346 20204 12348 20224
rect 12348 20204 12400 20224
rect 12400 20204 12402 20224
rect 12346 20168 12402 20204
rect 11610 18944 11666 19000
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11518 17856 11574 17912
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 10690 13524 10746 13560
rect 10690 13504 10692 13524
rect 10692 13504 10744 13524
rect 10744 13504 10746 13524
rect 11242 17176 11298 17232
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11518 15564 11574 15600
rect 11518 15544 11520 15564
rect 11520 15544 11572 15564
rect 11572 15544 11574 15564
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11610 15000 11666 15056
rect 11334 14592 11390 14648
rect 10874 12280 10930 12336
rect 10782 7928 10838 7984
rect 10690 6704 10746 6760
rect 10874 6160 10930 6216
rect 10782 4936 10838 4992
rect 10690 3848 10746 3904
rect 11242 14320 11298 14376
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11518 13404 11520 13424
rect 11520 13404 11572 13424
rect 11572 13404 11574 13424
rect 11518 13368 11574 13404
rect 12162 18808 12218 18864
rect 12530 18964 12586 19000
rect 12530 18944 12532 18964
rect 12532 18944 12584 18964
rect 12584 18944 12586 18964
rect 12714 17756 12716 17776
rect 12716 17756 12768 17776
rect 12768 17756 12770 17776
rect 12714 17720 12770 17756
rect 11794 13096 11850 13152
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11058 12552 11114 12608
rect 11058 12280 11114 12336
rect 11058 11892 11114 11928
rect 11058 11872 11060 11892
rect 11060 11872 11112 11892
rect 11112 11872 11114 11892
rect 11426 12280 11482 12336
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11610 11328 11666 11384
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11610 9288 11666 9344
rect 11610 9152 11666 9208
rect 11518 9016 11574 9072
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11702 7812 11758 7848
rect 11702 7792 11704 7812
rect 11704 7792 11756 7812
rect 11756 7792 11758 7812
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11150 5888 11206 5944
rect 11518 5888 11574 5944
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11702 5072 11758 5128
rect 11242 4664 11298 4720
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 3606 584 3662 640
rect 3238 176 3294 232
rect 12162 13948 12164 13968
rect 12164 13948 12216 13968
rect 12216 13948 12218 13968
rect 12162 13912 12218 13948
rect 12254 13640 12310 13696
rect 12622 17604 12678 17640
rect 12622 17584 12624 17604
rect 12624 17584 12676 17604
rect 12676 17584 12678 17604
rect 12438 15020 12494 15056
rect 12438 15000 12440 15020
rect 12440 15000 12492 15020
rect 12492 15000 12494 15020
rect 12438 14864 12494 14920
rect 12070 12824 12126 12880
rect 12070 12280 12126 12336
rect 12070 10104 12126 10160
rect 12070 9152 12126 9208
rect 12346 12552 12402 12608
rect 12254 10920 12310 10976
rect 12438 10104 12494 10160
rect 12438 8880 12494 8936
rect 12438 5344 12494 5400
rect 12622 15000 12678 15056
rect 12898 13812 12900 13832
rect 12900 13812 12952 13832
rect 12952 13812 12954 13832
rect 12898 13776 12954 13812
rect 12990 13504 13046 13560
rect 12622 12688 12678 12744
rect 12898 12280 12954 12336
rect 12806 6568 12862 6624
rect 12806 6296 12862 6352
rect 12622 4528 12678 4584
rect 12714 4256 12770 4312
rect 12622 3068 12624 3088
rect 12624 3068 12676 3088
rect 12676 3068 12678 3088
rect 12622 3032 12678 3068
rect 12806 4120 12862 4176
rect 13358 18264 13414 18320
rect 13266 17876 13322 17912
rect 13266 17856 13268 17876
rect 13268 17856 13320 17876
rect 13320 17856 13322 17876
rect 13358 17312 13414 17368
rect 13174 14592 13230 14648
rect 13082 12280 13138 12336
rect 14094 18672 14150 18728
rect 13542 17312 13598 17368
rect 13542 15680 13598 15736
rect 13174 12144 13230 12200
rect 13358 12552 13414 12608
rect 13358 12416 13414 12472
rect 13358 6976 13414 7032
rect 13542 5908 13598 5944
rect 13542 5888 13544 5908
rect 13544 5888 13596 5908
rect 13596 5888 13598 5908
rect 13818 12688 13874 12744
rect 13726 10648 13782 10704
rect 13726 10240 13782 10296
rect 13818 9016 13874 9072
rect 13542 4120 13598 4176
rect 13818 6060 13820 6080
rect 13820 6060 13872 6080
rect 13872 6060 13874 6080
rect 13818 6024 13874 6060
rect 13818 5888 13874 5944
rect 14186 16496 14242 16552
rect 14094 14320 14150 14376
rect 13818 3168 13874 3224
rect 14462 18128 14518 18184
rect 14370 17040 14426 17096
rect 14462 16496 14518 16552
rect 14554 13368 14610 13424
rect 14462 10532 14518 10568
rect 14462 10512 14464 10532
rect 14464 10512 14516 10532
rect 14516 10512 14518 10532
rect 14278 4664 14334 4720
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 15290 19760 15346 19816
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14646 6976 14702 7032
rect 14646 5908 14702 5944
rect 14646 5888 14648 5908
rect 14648 5888 14700 5908
rect 14700 5888 14702 5908
rect 14646 5344 14702 5400
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14830 11872 14886 11928
rect 15014 11872 15070 11928
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 15382 11328 15438 11384
rect 14830 10668 14886 10704
rect 14830 10648 14832 10668
rect 14832 10648 14884 10668
rect 14884 10648 14886 10668
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 15106 9968 15162 10024
rect 15382 10784 15438 10840
rect 15106 9424 15162 9480
rect 15382 9424 15438 9480
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 14922 7284 14924 7304
rect 14924 7284 14976 7304
rect 14976 7284 14978 7304
rect 14922 7248 14978 7284
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 15290 5208 15346 5264
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 15566 10784 15622 10840
rect 15566 10376 15622 10432
rect 15750 18128 15806 18184
rect 15934 17756 15936 17776
rect 15936 17756 15988 17776
rect 15988 17756 15990 17776
rect 15934 17720 15990 17756
rect 15750 17040 15806 17096
rect 15750 13368 15806 13424
rect 16762 18128 16818 18184
rect 16302 17176 16358 17232
rect 15934 12416 15990 12472
rect 16118 12144 16174 12200
rect 15750 10512 15806 10568
rect 16026 12008 16082 12064
rect 15658 8336 15714 8392
rect 15290 4120 15346 4176
rect 15842 6568 15898 6624
rect 15750 6296 15806 6352
rect 15658 5208 15714 5264
rect 15198 3712 15254 3768
rect 16118 8336 16174 8392
rect 16118 3848 16174 3904
rect 15750 3168 15806 3224
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 15474 2624 15530 2680
rect 16578 14864 16634 14920
rect 17130 19896 17186 19952
rect 17590 18128 17646 18184
rect 17958 22072 18014 22128
rect 18050 21120 18106 21176
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 17682 17992 17738 18048
rect 17222 17312 17278 17368
rect 16946 15000 17002 15056
rect 16670 11056 16726 11112
rect 16486 8472 16542 8528
rect 16394 7384 16450 7440
rect 16394 5072 16450 5128
rect 16394 4528 16450 4584
rect 16762 9560 16818 9616
rect 16578 7268 16634 7304
rect 16578 7248 16580 7268
rect 16580 7248 16632 7268
rect 16632 7248 16634 7268
rect 16486 3848 16542 3904
rect 17038 11328 17094 11384
rect 16946 7248 17002 7304
rect 16854 4684 16910 4720
rect 16854 4664 16856 4684
rect 16856 4664 16908 4684
rect 16908 4664 16910 4684
rect 16670 3576 16726 3632
rect 16762 3168 16818 3224
rect 17222 7792 17278 7848
rect 17130 7248 17186 7304
rect 17682 13388 17738 13424
rect 17682 13368 17684 13388
rect 17684 13368 17736 13388
rect 17736 13368 17738 13388
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 17682 12552 17738 12608
rect 17682 12280 17738 12336
rect 18050 16088 18106 16144
rect 17958 15000 18014 15056
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18786 21528 18842 21584
rect 18694 20576 18750 20632
rect 18694 19624 18750 19680
rect 18878 18808 18934 18864
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18142 14320 18198 14376
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18050 13640 18106 13696
rect 18142 13368 18198 13424
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18234 12824 18290 12880
rect 18050 12552 18106 12608
rect 18050 12416 18106 12472
rect 17958 11736 18014 11792
rect 18142 12280 18198 12336
rect 18878 17040 18934 17096
rect 18786 14048 18842 14104
rect 18418 12416 18474 12472
rect 17774 11464 17830 11520
rect 17498 6840 17554 6896
rect 17866 10920 17922 10976
rect 18050 7384 18106 7440
rect 18050 7112 18106 7168
rect 17590 5072 17646 5128
rect 17774 4664 17830 4720
rect 17774 3576 17830 3632
rect 18786 12280 18842 12336
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18234 10104 18290 10160
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18234 9288 18290 9344
rect 18234 8900 18290 8936
rect 18234 8880 18236 8900
rect 18236 8880 18288 8900
rect 18288 8880 18290 8900
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18142 3848 18198 3904
rect 18326 3712 18382 3768
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18786 8608 18842 8664
rect 18878 7284 18880 7304
rect 18880 7284 18932 7304
rect 18932 7284 18934 7304
rect 18878 7248 18934 7284
rect 18878 6180 18934 6216
rect 18878 6160 18880 6180
rect 18880 6160 18932 6180
rect 18932 6160 18934 6180
rect 19154 20032 19210 20088
rect 19246 17584 19302 17640
rect 19062 14320 19118 14376
rect 18878 4528 18934 4584
rect 19246 7656 19302 7712
rect 19154 6704 19210 6760
rect 19246 6568 19302 6624
rect 19246 5752 19302 5808
rect 19154 5616 19210 5672
rect 19614 10648 19670 10704
rect 19430 2508 19486 2544
rect 19430 2488 19432 2508
rect 19432 2488 19484 2508
rect 19484 2488 19486 2508
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 18694 2080 18750 2136
rect 20718 18536 20774 18592
rect 20074 14456 20130 14512
rect 20074 12552 20130 12608
rect 19890 3984 19946 4040
rect 20350 12144 20406 12200
rect 20534 9968 20590 10024
rect 20534 9696 20590 9752
rect 20626 7112 20682 7168
rect 20994 3440 21050 3496
rect 20534 3168 20590 3224
rect 18510 1672 18566 1728
rect 12070 1128 12126 1184
rect 18142 584 18198 640
rect 21178 3032 21234 3088
rect 21270 2896 21326 2952
rect 22374 5072 22430 5128
rect 22374 4936 22430 4992
rect 11886 176 11942 232
<< metal3 >>
rect 0 22674 480 22704
rect 3693 22674 3759 22677
rect 0 22672 3759 22674
rect 0 22616 3698 22672
rect 3754 22616 3759 22672
rect 0 22614 3759 22616
rect 0 22584 480 22614
rect 3693 22611 3759 22614
rect 17861 22674 17927 22677
rect 22520 22674 23000 22704
rect 17861 22672 23000 22674
rect 17861 22616 17866 22672
rect 17922 22616 23000 22672
rect 17861 22614 23000 22616
rect 17861 22611 17927 22614
rect 22520 22584 23000 22614
rect 0 22130 480 22160
rect 3509 22130 3575 22133
rect 0 22128 3575 22130
rect 0 22072 3514 22128
rect 3570 22072 3575 22128
rect 0 22070 3575 22072
rect 0 22040 480 22070
rect 3509 22067 3575 22070
rect 17953 22130 18019 22133
rect 22520 22130 23000 22160
rect 17953 22128 23000 22130
rect 17953 22072 17958 22128
rect 18014 22072 23000 22128
rect 17953 22070 23000 22072
rect 17953 22067 18019 22070
rect 22520 22040 23000 22070
rect 0 21586 480 21616
rect 3509 21586 3575 21589
rect 0 21584 3575 21586
rect 0 21528 3514 21584
rect 3570 21528 3575 21584
rect 0 21526 3575 21528
rect 0 21496 480 21526
rect 3509 21523 3575 21526
rect 18781 21586 18847 21589
rect 22520 21586 23000 21616
rect 18781 21584 23000 21586
rect 18781 21528 18786 21584
rect 18842 21528 23000 21584
rect 18781 21526 23000 21528
rect 18781 21523 18847 21526
rect 22520 21496 23000 21526
rect 0 21178 480 21208
rect 2957 21178 3023 21181
rect 0 21176 3023 21178
rect 0 21120 2962 21176
rect 3018 21120 3023 21176
rect 0 21118 3023 21120
rect 0 21088 480 21118
rect 2957 21115 3023 21118
rect 18045 21178 18111 21181
rect 22520 21178 23000 21208
rect 18045 21176 23000 21178
rect 18045 21120 18050 21176
rect 18106 21120 23000 21176
rect 18045 21118 23000 21120
rect 18045 21115 18111 21118
rect 22520 21088 23000 21118
rect 4409 20704 4729 20705
rect 0 20634 480 20664
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 1945 20634 2011 20637
rect 0 20632 2011 20634
rect 0 20576 1950 20632
rect 2006 20576 2011 20632
rect 0 20574 2011 20576
rect 0 20544 480 20574
rect 1945 20571 2011 20574
rect 18689 20634 18755 20637
rect 22520 20634 23000 20664
rect 18689 20632 23000 20634
rect 18689 20576 18694 20632
rect 18750 20576 23000 20632
rect 18689 20574 23000 20576
rect 18689 20571 18755 20574
rect 22520 20544 23000 20574
rect 8293 20364 8359 20365
rect 8293 20360 8340 20364
rect 8404 20362 8410 20364
rect 8293 20304 8298 20360
rect 8293 20300 8340 20304
rect 8404 20302 8450 20362
rect 8404 20300 8410 20302
rect 8293 20299 8359 20300
rect 8477 20226 8543 20229
rect 8845 20226 8911 20229
rect 8477 20224 8911 20226
rect 8477 20168 8482 20224
rect 8538 20168 8850 20224
rect 8906 20168 8911 20224
rect 8477 20166 8911 20168
rect 8477 20163 8543 20166
rect 8845 20163 8911 20166
rect 10961 20226 11027 20229
rect 12341 20226 12407 20229
rect 10961 20224 12407 20226
rect 10961 20168 10966 20224
rect 11022 20168 12346 20224
rect 12402 20168 12407 20224
rect 10961 20166 12407 20168
rect 10961 20163 11027 20166
rect 12341 20163 12407 20166
rect 7874 20160 8194 20161
rect 0 20090 480 20120
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 3969 20090 4035 20093
rect 0 20088 4035 20090
rect 0 20032 3974 20088
rect 4030 20032 4035 20088
rect 0 20030 4035 20032
rect 0 20000 480 20030
rect 3969 20027 4035 20030
rect 19149 20090 19215 20093
rect 22520 20090 23000 20120
rect 19149 20088 23000 20090
rect 19149 20032 19154 20088
rect 19210 20032 23000 20088
rect 19149 20030 23000 20032
rect 19149 20027 19215 20030
rect 22520 20000 23000 20030
rect 8477 19954 8543 19957
rect 17125 19954 17191 19957
rect 8477 19952 17191 19954
rect 8477 19896 8482 19952
rect 8538 19896 17130 19952
rect 17186 19896 17191 19952
rect 8477 19894 17191 19896
rect 8477 19891 8543 19894
rect 17125 19891 17191 19894
rect 8385 19818 8451 19821
rect 15285 19818 15351 19821
rect 8385 19816 15351 19818
rect 8385 19760 8390 19816
rect 8446 19760 15290 19816
rect 15346 19760 15351 19816
rect 8385 19758 15351 19760
rect 8385 19755 8451 19758
rect 15285 19755 15351 19758
rect 0 19682 480 19712
rect 4245 19682 4311 19685
rect 0 19680 4311 19682
rect 0 19624 4250 19680
rect 4306 19624 4311 19680
rect 0 19622 4311 19624
rect 0 19592 480 19622
rect 4245 19619 4311 19622
rect 18689 19682 18755 19685
rect 22520 19682 23000 19712
rect 18689 19680 23000 19682
rect 18689 19624 18694 19680
rect 18750 19624 23000 19680
rect 18689 19622 23000 19624
rect 18689 19619 18755 19622
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 22520 19592 23000 19622
rect 18270 19551 18590 19552
rect 5809 19274 5875 19277
rect 8201 19274 8267 19277
rect 5809 19272 8267 19274
rect 5809 19216 5814 19272
rect 5870 19216 8206 19272
rect 8262 19216 8267 19272
rect 5809 19214 8267 19216
rect 5809 19211 5875 19214
rect 8201 19211 8267 19214
rect 8477 19274 8543 19277
rect 8477 19272 15394 19274
rect 8477 19216 8482 19272
rect 8538 19216 15394 19272
rect 8477 19214 15394 19216
rect 8477 19211 8543 19214
rect 0 19138 480 19168
rect 8293 19140 8359 19141
rect 0 19078 674 19138
rect 0 19048 480 19078
rect 13 18866 79 18869
rect 614 18866 674 19078
rect 8293 19136 8340 19140
rect 8404 19138 8410 19140
rect 15334 19138 15394 19214
rect 22520 19138 23000 19168
rect 8293 19080 8298 19136
rect 8293 19076 8340 19080
rect 8404 19078 8450 19138
rect 15334 19078 23000 19138
rect 8404 19076 8410 19078
rect 8293 19075 8359 19076
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 22520 19048 23000 19078
rect 14805 19007 15125 19008
rect 1393 19002 1459 19005
rect 7189 19002 7255 19005
rect 1393 19000 7255 19002
rect 1393 18944 1398 19000
rect 1454 18944 7194 19000
rect 7250 18944 7255 19000
rect 1393 18942 7255 18944
rect 1393 18939 1459 18942
rect 7189 18939 7255 18942
rect 11605 19002 11671 19005
rect 12525 19002 12591 19005
rect 11605 19000 12591 19002
rect 11605 18944 11610 19000
rect 11666 18944 12530 19000
rect 12586 18944 12591 19000
rect 11605 18942 12591 18944
rect 11605 18939 11671 18942
rect 12525 18939 12591 18942
rect 13 18864 674 18866
rect 13 18808 18 18864
rect 74 18808 674 18864
rect 13 18806 674 18808
rect 4797 18866 4863 18869
rect 5574 18866 5580 18868
rect 4797 18864 5580 18866
rect 4797 18808 4802 18864
rect 4858 18808 5580 18864
rect 4797 18806 5580 18808
rect 13 18803 79 18806
rect 4797 18803 4863 18806
rect 5574 18804 5580 18806
rect 5644 18804 5650 18868
rect 12157 18866 12223 18869
rect 18873 18866 18939 18869
rect 12157 18864 18939 18866
rect 12157 18808 12162 18864
rect 12218 18808 18878 18864
rect 18934 18808 18939 18864
rect 12157 18806 18939 18808
rect 12157 18803 12223 18806
rect 18873 18803 18939 18806
rect 4061 18730 4127 18733
rect 10501 18730 10567 18733
rect 4061 18728 10567 18730
rect 4061 18672 4066 18728
rect 4122 18672 10506 18728
rect 10562 18672 10567 18728
rect 4061 18670 10567 18672
rect 4061 18667 4127 18670
rect 10501 18667 10567 18670
rect 14089 18730 14155 18733
rect 14590 18730 14596 18732
rect 14089 18728 14596 18730
rect 14089 18672 14094 18728
rect 14150 18672 14596 18728
rect 14089 18670 14596 18672
rect 14089 18667 14155 18670
rect 14590 18668 14596 18670
rect 14660 18668 14666 18732
rect 0 18594 480 18624
rect 1393 18594 1459 18597
rect 0 18592 1459 18594
rect 0 18536 1398 18592
rect 1454 18536 1459 18592
rect 0 18534 1459 18536
rect 0 18504 480 18534
rect 1393 18531 1459 18534
rect 6637 18594 6703 18597
rect 8569 18594 8635 18597
rect 6637 18592 8635 18594
rect 6637 18536 6642 18592
rect 6698 18536 8574 18592
rect 8630 18536 8635 18592
rect 6637 18534 8635 18536
rect 6637 18531 6703 18534
rect 8569 18531 8635 18534
rect 20713 18594 20779 18597
rect 22520 18594 23000 18624
rect 20713 18592 23000 18594
rect 20713 18536 20718 18592
rect 20774 18536 23000 18592
rect 20713 18534 23000 18536
rect 20713 18531 20779 18534
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 22520 18504 23000 18534
rect 18270 18463 18590 18464
rect 3509 18322 3575 18325
rect 13353 18322 13419 18325
rect 3509 18320 13419 18322
rect 3509 18264 3514 18320
rect 3570 18264 13358 18320
rect 13414 18264 13419 18320
rect 3509 18262 13419 18264
rect 3509 18259 3575 18262
rect 13353 18259 13419 18262
rect 0 18186 480 18216
rect 3141 18186 3207 18189
rect 0 18184 3207 18186
rect 0 18128 3146 18184
rect 3202 18128 3207 18184
rect 0 18126 3207 18128
rect 0 18096 480 18126
rect 3141 18123 3207 18126
rect 6729 18186 6795 18189
rect 8753 18186 8819 18189
rect 6729 18184 8819 18186
rect 6729 18128 6734 18184
rect 6790 18128 8758 18184
rect 8814 18128 8819 18184
rect 6729 18126 8819 18128
rect 6729 18123 6795 18126
rect 8753 18123 8819 18126
rect 9213 18186 9279 18189
rect 14457 18186 14523 18189
rect 9213 18184 14523 18186
rect 9213 18128 9218 18184
rect 9274 18128 14462 18184
rect 14518 18128 14523 18184
rect 9213 18126 14523 18128
rect 9213 18123 9279 18126
rect 14457 18123 14523 18126
rect 15745 18186 15811 18189
rect 16757 18186 16823 18189
rect 17585 18186 17651 18189
rect 15745 18184 17651 18186
rect 15745 18128 15750 18184
rect 15806 18128 16762 18184
rect 16818 18128 17590 18184
rect 17646 18128 17651 18184
rect 15745 18126 17651 18128
rect 15745 18123 15811 18126
rect 16757 18123 16823 18126
rect 17585 18123 17651 18126
rect 17718 18124 17724 18188
rect 17788 18186 17794 18188
rect 22520 18186 23000 18216
rect 17788 18126 23000 18186
rect 17788 18124 17794 18126
rect 22520 18096 23000 18126
rect 16614 17988 16620 18052
rect 16684 18050 16690 18052
rect 17677 18050 17743 18053
rect 16684 18048 17743 18050
rect 16684 17992 17682 18048
rect 17738 17992 17743 18048
rect 16684 17990 17743 17992
rect 16684 17988 16690 17990
rect 17677 17987 17743 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 17919 15125 17920
rect 11513 17914 11579 17917
rect 13261 17914 13327 17917
rect 11513 17912 13327 17914
rect 11513 17856 11518 17912
rect 11574 17856 13266 17912
rect 13322 17856 13327 17912
rect 11513 17854 13327 17856
rect 11513 17851 11579 17854
rect 13261 17851 13327 17854
rect 12709 17778 12775 17781
rect 15929 17778 15995 17781
rect 12709 17776 15995 17778
rect 12709 17720 12714 17776
rect 12770 17720 15934 17776
rect 15990 17720 15995 17776
rect 12709 17718 15995 17720
rect 12709 17715 12775 17718
rect 15929 17715 15995 17718
rect 0 17642 480 17672
rect 3233 17642 3299 17645
rect 0 17640 3299 17642
rect 0 17584 3238 17640
rect 3294 17584 3299 17640
rect 0 17582 3299 17584
rect 0 17552 480 17582
rect 3233 17579 3299 17582
rect 10869 17642 10935 17645
rect 12617 17642 12683 17645
rect 10869 17640 12683 17642
rect 10869 17584 10874 17640
rect 10930 17584 12622 17640
rect 12678 17584 12683 17640
rect 10869 17582 12683 17584
rect 10869 17579 10935 17582
rect 12617 17579 12683 17582
rect 19241 17642 19307 17645
rect 22520 17642 23000 17672
rect 19241 17640 23000 17642
rect 19241 17584 19246 17640
rect 19302 17584 23000 17640
rect 19241 17582 23000 17584
rect 19241 17579 19307 17582
rect 22520 17552 23000 17582
rect 6913 17506 6979 17509
rect 10961 17506 11027 17509
rect 6913 17504 11027 17506
rect 6913 17448 6918 17504
rect 6974 17448 10966 17504
rect 11022 17448 11027 17504
rect 6913 17446 11027 17448
rect 6913 17443 6979 17446
rect 10961 17443 11027 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 13353 17372 13419 17373
rect 13302 17308 13308 17372
rect 13372 17370 13419 17372
rect 13537 17370 13603 17373
rect 17217 17370 17283 17373
rect 13372 17368 13464 17370
rect 13414 17312 13464 17368
rect 13372 17310 13464 17312
rect 13537 17368 17283 17370
rect 13537 17312 13542 17368
rect 13598 17312 17222 17368
rect 17278 17312 17283 17368
rect 13537 17310 17283 17312
rect 13372 17308 13419 17310
rect 13353 17307 13419 17308
rect 13537 17307 13603 17310
rect 17217 17307 17283 17310
rect 2037 17234 2103 17237
rect 8518 17234 8524 17236
rect 2037 17232 8524 17234
rect 2037 17176 2042 17232
rect 2098 17176 8524 17232
rect 2037 17174 8524 17176
rect 2037 17171 2103 17174
rect 8518 17172 8524 17174
rect 8588 17172 8594 17236
rect 11237 17234 11303 17237
rect 16297 17234 16363 17237
rect 11237 17232 16363 17234
rect 11237 17176 11242 17232
rect 11298 17176 16302 17232
rect 16358 17176 16363 17232
rect 11237 17174 16363 17176
rect 11237 17171 11303 17174
rect 16297 17171 16363 17174
rect 0 17098 480 17128
rect 1761 17098 1827 17101
rect 14365 17098 14431 17101
rect 15745 17098 15811 17101
rect 0 17096 1827 17098
rect 0 17040 1766 17096
rect 1822 17040 1827 17096
rect 0 17038 1827 17040
rect 0 17008 480 17038
rect 1761 17035 1827 17038
rect 1902 17096 14431 17098
rect 1902 17040 14370 17096
rect 14426 17040 14431 17096
rect 1902 17038 14431 17040
rect 1209 16962 1275 16965
rect 1902 16962 1962 17038
rect 14365 17035 14431 17038
rect 14598 17096 15811 17098
rect 14598 17040 15750 17096
rect 15806 17040 15811 17096
rect 14598 17038 15811 17040
rect 1209 16960 1962 16962
rect 1209 16904 1214 16960
rect 1270 16904 1962 16960
rect 1209 16902 1962 16904
rect 9305 16962 9371 16965
rect 14598 16962 14658 17038
rect 15745 17035 15811 17038
rect 18873 17098 18939 17101
rect 22520 17098 23000 17128
rect 18873 17096 23000 17098
rect 18873 17040 18878 17096
rect 18934 17040 23000 17096
rect 18873 17038 23000 17040
rect 18873 17035 18939 17038
rect 22520 17008 23000 17038
rect 9305 16960 14658 16962
rect 9305 16904 9310 16960
rect 9366 16904 14658 16960
rect 9305 16902 14658 16904
rect 1209 16899 1275 16902
rect 9305 16899 9371 16902
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 0 16690 480 16720
rect 3601 16690 3667 16693
rect 0 16688 3667 16690
rect 0 16632 3606 16688
rect 3662 16632 3667 16688
rect 0 16630 3667 16632
rect 0 16600 480 16630
rect 3601 16627 3667 16630
rect 5206 16628 5212 16692
rect 5276 16690 5282 16692
rect 5349 16690 5415 16693
rect 5276 16688 5415 16690
rect 5276 16632 5354 16688
rect 5410 16632 5415 16688
rect 5276 16630 5415 16632
rect 5276 16628 5282 16630
rect 5349 16627 5415 16630
rect 8201 16690 8267 16693
rect 17718 16690 17724 16692
rect 8201 16688 17724 16690
rect 8201 16632 8206 16688
rect 8262 16632 17724 16688
rect 8201 16630 17724 16632
rect 8201 16627 8267 16630
rect 17718 16628 17724 16630
rect 17788 16628 17794 16692
rect 22520 16690 23000 16720
rect 17864 16630 23000 16690
rect 2681 16554 2747 16557
rect 14181 16554 14247 16557
rect 2681 16552 14247 16554
rect 2681 16496 2686 16552
rect 2742 16496 14186 16552
rect 14242 16496 14247 16552
rect 2681 16494 14247 16496
rect 2681 16491 2747 16494
rect 14181 16491 14247 16494
rect 14457 16554 14523 16557
rect 17864 16554 17924 16630
rect 22520 16600 23000 16630
rect 14457 16552 17924 16554
rect 14457 16496 14462 16552
rect 14518 16496 17924 16552
rect 14457 16494 17924 16496
rect 14457 16491 14523 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16146 480 16176
rect 1669 16146 1735 16149
rect 0 16144 1735 16146
rect 0 16088 1674 16144
rect 1730 16088 1735 16144
rect 0 16086 1735 16088
rect 0 16056 480 16086
rect 1669 16083 1735 16086
rect 18045 16146 18111 16149
rect 22520 16146 23000 16176
rect 18045 16144 23000 16146
rect 18045 16088 18050 16144
rect 18106 16088 23000 16144
rect 18045 16086 23000 16088
rect 18045 16083 18111 16086
rect 22520 16056 23000 16086
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 9673 15738 9739 15741
rect 13537 15738 13603 15741
rect 9673 15736 13603 15738
rect 9673 15680 9678 15736
rect 9734 15680 13542 15736
rect 13598 15680 13603 15736
rect 9673 15678 13603 15680
rect 9673 15675 9739 15678
rect 13537 15675 13603 15678
rect 0 15602 480 15632
rect 4061 15602 4127 15605
rect 0 15600 4127 15602
rect 0 15544 4066 15600
rect 4122 15544 4127 15600
rect 0 15542 4127 15544
rect 0 15512 480 15542
rect 4061 15539 4127 15542
rect 11513 15602 11579 15605
rect 22520 15602 23000 15632
rect 11513 15600 23000 15602
rect 11513 15544 11518 15600
rect 11574 15544 23000 15600
rect 11513 15542 23000 15544
rect 11513 15539 11579 15542
rect 22520 15512 23000 15542
rect 4409 15264 4729 15265
rect 0 15194 480 15224
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 4061 15194 4127 15197
rect 0 15192 4127 15194
rect 0 15136 4066 15192
rect 4122 15136 4127 15192
rect 0 15134 4127 15136
rect 0 15104 480 15134
rect 4061 15131 4127 15134
rect 7230 15132 7236 15196
rect 7300 15194 7306 15196
rect 7741 15194 7807 15197
rect 22520 15194 23000 15224
rect 7300 15192 7807 15194
rect 7300 15136 7746 15192
rect 7802 15136 7807 15192
rect 7300 15134 7807 15136
rect 7300 15132 7306 15134
rect 7741 15131 7807 15134
rect 18830 15134 23000 15194
rect 2957 15058 3023 15061
rect 3366 15058 3372 15060
rect 2957 15056 3372 15058
rect 2957 15000 2962 15056
rect 3018 15000 3372 15056
rect 2957 14998 3372 15000
rect 2957 14995 3023 14998
rect 3366 14996 3372 14998
rect 3436 14996 3442 15060
rect 11605 15058 11671 15061
rect 12433 15058 12499 15061
rect 12617 15058 12683 15061
rect 11605 15056 12683 15058
rect 11605 15000 11610 15056
rect 11666 15000 12438 15056
rect 12494 15000 12622 15056
rect 12678 15000 12683 15056
rect 11605 14998 12683 15000
rect 11605 14995 11671 14998
rect 12433 14995 12499 14998
rect 12617 14995 12683 14998
rect 16941 15060 17007 15061
rect 16941 15056 16988 15060
rect 17052 15058 17058 15060
rect 17953 15058 18019 15061
rect 18830 15058 18890 15134
rect 22520 15104 23000 15134
rect 16941 15000 16946 15056
rect 16941 14996 16988 15000
rect 17052 14998 17098 15058
rect 17953 15056 18890 15058
rect 17953 15000 17958 15056
rect 18014 15000 18890 15056
rect 17953 14998 18890 15000
rect 17052 14996 17058 14998
rect 16941 14995 17007 14996
rect 17953 14995 18019 14998
rect 4981 14922 5047 14925
rect 5717 14922 5783 14925
rect 11830 14922 11836 14924
rect 4981 14920 5274 14922
rect 4981 14864 4986 14920
rect 5042 14864 5274 14920
rect 4981 14862 5274 14864
rect 4981 14859 5047 14862
rect 0 14650 480 14680
rect 3509 14650 3575 14653
rect 0 14648 3575 14650
rect 0 14592 3514 14648
rect 3570 14592 3575 14648
rect 0 14590 3575 14592
rect 0 14560 480 14590
rect 3509 14587 3575 14590
rect 4889 14514 4955 14517
rect 4846 14512 4955 14514
rect 4846 14456 4894 14512
rect 4950 14456 4955 14512
rect 4846 14451 4955 14456
rect 4409 14176 4729 14177
rect 0 14106 480 14136
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 3969 14106 4035 14109
rect 0 14104 4035 14106
rect 0 14048 3974 14104
rect 4030 14048 4035 14104
rect 0 14046 4035 14048
rect 0 14016 480 14046
rect 3969 14043 4035 14046
rect 4846 13837 4906 14451
rect 5214 14242 5274 14862
rect 5717 14920 11836 14922
rect 5717 14864 5722 14920
rect 5778 14864 11836 14920
rect 5717 14862 11836 14864
rect 5717 14859 5783 14862
rect 11830 14860 11836 14862
rect 11900 14860 11906 14924
rect 12433 14922 12499 14925
rect 16573 14922 16639 14925
rect 12433 14920 16639 14922
rect 12433 14864 12438 14920
rect 12494 14864 16578 14920
rect 16634 14864 16639 14920
rect 12433 14862 16639 14864
rect 12433 14859 12499 14862
rect 16573 14859 16639 14862
rect 7874 14720 8194 14721
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 11329 14650 11395 14653
rect 13169 14650 13235 14653
rect 22520 14650 23000 14680
rect 11329 14648 13235 14650
rect 11329 14592 11334 14648
rect 11390 14592 13174 14648
rect 13230 14592 13235 14648
rect 11329 14590 13235 14592
rect 11329 14587 11395 14590
rect 13169 14587 13235 14590
rect 15518 14590 23000 14650
rect 13118 14452 13124 14516
rect 13188 14514 13194 14516
rect 15518 14514 15578 14590
rect 22520 14560 23000 14590
rect 13188 14454 15578 14514
rect 13188 14452 13194 14454
rect 19742 14452 19748 14516
rect 19812 14514 19818 14516
rect 20069 14514 20135 14517
rect 19812 14512 20135 14514
rect 19812 14456 20074 14512
rect 20130 14456 20135 14512
rect 19812 14454 20135 14456
rect 19812 14452 19818 14454
rect 20069 14451 20135 14454
rect 11094 14316 11100 14380
rect 11164 14378 11170 14380
rect 11237 14378 11303 14381
rect 11164 14376 11303 14378
rect 11164 14320 11242 14376
rect 11298 14320 11303 14376
rect 11164 14318 11303 14320
rect 11164 14316 11170 14318
rect 11237 14315 11303 14318
rect 14089 14378 14155 14381
rect 15694 14378 15700 14380
rect 14089 14376 15700 14378
rect 14089 14320 14094 14376
rect 14150 14320 15700 14376
rect 14089 14318 15700 14320
rect 14089 14315 14155 14318
rect 15694 14316 15700 14318
rect 15764 14316 15770 14380
rect 17902 14316 17908 14380
rect 17972 14378 17978 14380
rect 18137 14378 18203 14381
rect 19057 14380 19123 14381
rect 17972 14376 18203 14378
rect 17972 14320 18142 14376
rect 18198 14320 18203 14376
rect 17972 14318 18203 14320
rect 17972 14316 17978 14318
rect 18137 14315 18203 14318
rect 19006 14316 19012 14380
rect 19076 14378 19123 14380
rect 19076 14376 19168 14378
rect 19118 14320 19168 14376
rect 19076 14318 19168 14320
rect 19076 14316 19123 14318
rect 19057 14315 19123 14316
rect 5349 14242 5415 14245
rect 5214 14240 5415 14242
rect 5214 14184 5354 14240
rect 5410 14184 5415 14240
rect 5214 14182 5415 14184
rect 5349 14179 5415 14182
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 18781 14106 18847 14109
rect 22520 14106 23000 14136
rect 18781 14104 23000 14106
rect 18781 14048 18786 14104
rect 18842 14048 23000 14104
rect 18781 14046 23000 14048
rect 18781 14043 18847 14046
rect 22520 14016 23000 14046
rect 10409 13970 10475 13973
rect 12157 13970 12223 13973
rect 10409 13968 12223 13970
rect 10409 13912 10414 13968
rect 10470 13912 12162 13968
rect 12218 13912 12223 13968
rect 10409 13910 12223 13912
rect 10409 13907 10475 13910
rect 12157 13907 12223 13910
rect 4846 13832 4955 13837
rect 4846 13776 4894 13832
rect 4950 13776 4955 13832
rect 4846 13774 4955 13776
rect 4889 13771 4955 13774
rect 9581 13834 9647 13837
rect 12893 13834 12959 13837
rect 9581 13832 12959 13834
rect 9581 13776 9586 13832
rect 9642 13776 12898 13832
rect 12954 13776 12959 13832
rect 9581 13774 12959 13776
rect 9581 13771 9647 13774
rect 12893 13771 12959 13774
rect 0 13698 480 13728
rect 3969 13698 4035 13701
rect 0 13696 4035 13698
rect 0 13640 3974 13696
rect 4030 13640 4035 13696
rect 0 13638 4035 13640
rect 0 13608 480 13638
rect 3969 13635 4035 13638
rect 10174 13636 10180 13700
rect 10244 13698 10250 13700
rect 12249 13698 12315 13701
rect 10244 13696 12315 13698
rect 10244 13640 12254 13696
rect 12310 13640 12315 13696
rect 10244 13638 12315 13640
rect 10244 13636 10250 13638
rect 12249 13635 12315 13638
rect 18045 13698 18111 13701
rect 22520 13698 23000 13728
rect 18045 13696 23000 13698
rect 18045 13640 18050 13696
rect 18106 13640 23000 13696
rect 18045 13638 23000 13640
rect 18045 13635 18111 13638
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 22520 13608 23000 13638
rect 14805 13567 15125 13568
rect 10685 13562 10751 13565
rect 12985 13562 13051 13565
rect 10685 13560 13051 13562
rect 10685 13504 10690 13560
rect 10746 13504 12990 13560
rect 13046 13504 13051 13560
rect 10685 13502 13051 13504
rect 10685 13499 10751 13502
rect 12985 13499 13051 13502
rect 11513 13426 11579 13429
rect 14549 13426 14615 13429
rect 11513 13424 14615 13426
rect 11513 13368 11518 13424
rect 11574 13368 14554 13424
rect 14610 13368 14615 13424
rect 11513 13366 14615 13368
rect 11513 13363 11579 13366
rect 14549 13363 14615 13366
rect 15745 13426 15811 13429
rect 17677 13426 17743 13429
rect 18137 13426 18203 13429
rect 15745 13424 18203 13426
rect 15745 13368 15750 13424
rect 15806 13368 17682 13424
rect 17738 13368 18142 13424
rect 18198 13368 18203 13424
rect 15745 13366 18203 13368
rect 15745 13363 15811 13366
rect 17677 13363 17743 13366
rect 18137 13363 18203 13366
rect 1117 13290 1183 13293
rect 9489 13290 9555 13293
rect 1117 13288 9555 13290
rect 1117 13232 1122 13288
rect 1178 13232 9494 13288
rect 9550 13232 9555 13288
rect 1117 13230 9555 13232
rect 1117 13227 1183 13230
rect 9489 13227 9555 13230
rect 0 13154 480 13184
rect 3785 13154 3851 13157
rect 0 13152 3851 13154
rect 0 13096 3790 13152
rect 3846 13096 3851 13152
rect 0 13094 3851 13096
rect 0 13064 480 13094
rect 3785 13091 3851 13094
rect 11789 13154 11855 13157
rect 22520 13154 23000 13184
rect 11789 13152 12082 13154
rect 11789 13096 11794 13152
rect 11850 13096 12082 13152
rect 11789 13094 12082 13096
rect 11789 13091 11855 13094
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 12022 12885 12082 13094
rect 18830 13094 23000 13154
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 12022 12880 12131 12885
rect 12022 12824 12070 12880
rect 12126 12824 12131 12880
rect 12022 12822 12131 12824
rect 12065 12819 12131 12822
rect 18229 12882 18295 12885
rect 18830 12882 18890 13094
rect 22520 13064 23000 13094
rect 18229 12880 18890 12882
rect 18229 12824 18234 12880
rect 18290 12824 18890 12880
rect 18229 12822 18890 12824
rect 18229 12819 18295 12822
rect 12617 12746 12683 12749
rect 13813 12746 13879 12749
rect 12617 12744 13879 12746
rect 12617 12688 12622 12744
rect 12678 12688 13818 12744
rect 13874 12688 13879 12744
rect 12617 12686 13879 12688
rect 12617 12683 12683 12686
rect 13813 12683 13879 12686
rect 0 12610 480 12640
rect 3877 12610 3943 12613
rect 0 12608 3943 12610
rect 0 12552 3882 12608
rect 3938 12552 3943 12608
rect 0 12550 3943 12552
rect 0 12520 480 12550
rect 3877 12547 3943 12550
rect 5073 12610 5139 12613
rect 5206 12610 5212 12612
rect 5073 12608 5212 12610
rect 5073 12552 5078 12608
rect 5134 12552 5212 12608
rect 5073 12550 5212 12552
rect 5073 12547 5139 12550
rect 5206 12548 5212 12550
rect 5276 12548 5282 12612
rect 11053 12610 11119 12613
rect 12341 12610 12407 12613
rect 11053 12608 12407 12610
rect 11053 12552 11058 12608
rect 11114 12552 12346 12608
rect 12402 12552 12407 12608
rect 11053 12550 12407 12552
rect 11053 12547 11119 12550
rect 12341 12547 12407 12550
rect 12934 12548 12940 12612
rect 13004 12610 13010 12612
rect 13353 12610 13419 12613
rect 13004 12608 13419 12610
rect 13004 12552 13358 12608
rect 13414 12552 13419 12608
rect 13004 12550 13419 12552
rect 13004 12548 13010 12550
rect 13353 12547 13419 12550
rect 17677 12610 17743 12613
rect 18045 12612 18111 12613
rect 17677 12608 17786 12610
rect 17677 12552 17682 12608
rect 17738 12552 17786 12608
rect 17677 12547 17786 12552
rect 18045 12608 18092 12612
rect 18156 12610 18162 12612
rect 20069 12610 20135 12613
rect 22520 12610 23000 12640
rect 18045 12552 18050 12608
rect 18045 12548 18092 12552
rect 18156 12550 18202 12610
rect 20069 12608 23000 12610
rect 20069 12552 20074 12608
rect 20130 12552 23000 12608
rect 20069 12550 23000 12552
rect 18156 12548 18162 12550
rect 18045 12547 18111 12548
rect 20069 12547 20135 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 1853 12476 1919 12477
rect 1853 12472 1900 12476
rect 1964 12474 1970 12476
rect 2221 12474 2287 12477
rect 5257 12476 5323 12477
rect 5441 12476 5507 12477
rect 2446 12474 2452 12476
rect 1853 12416 1858 12472
rect 1853 12412 1900 12416
rect 1964 12414 2010 12474
rect 2221 12472 2452 12474
rect 2221 12416 2226 12472
rect 2282 12416 2452 12472
rect 2221 12414 2452 12416
rect 1964 12412 1970 12414
rect 1853 12411 1919 12412
rect 2221 12411 2287 12414
rect 2446 12412 2452 12414
rect 2516 12412 2522 12476
rect 5206 12474 5212 12476
rect 5166 12414 5212 12474
rect 5276 12472 5323 12476
rect 5318 12416 5323 12472
rect 5206 12412 5212 12414
rect 5276 12412 5323 12416
rect 5390 12412 5396 12476
rect 5460 12474 5507 12476
rect 6453 12474 6519 12477
rect 6821 12474 6887 12477
rect 13353 12476 13419 12477
rect 13302 12474 13308 12476
rect 5460 12472 5552 12474
rect 5502 12416 5552 12472
rect 5460 12414 5552 12416
rect 6453 12472 6887 12474
rect 6453 12416 6458 12472
rect 6514 12416 6826 12472
rect 6882 12416 6887 12472
rect 6453 12414 6887 12416
rect 13262 12414 13308 12474
rect 13372 12472 13419 12476
rect 13414 12416 13419 12472
rect 5460 12412 5507 12414
rect 5257 12411 5323 12412
rect 5441 12411 5507 12412
rect 6453 12411 6519 12414
rect 6821 12411 6887 12414
rect 13302 12412 13308 12414
rect 13372 12412 13419 12416
rect 13353 12411 13419 12412
rect 15929 12474 15995 12477
rect 16062 12474 16068 12476
rect 15929 12472 16068 12474
rect 15929 12416 15934 12472
rect 15990 12416 16068 12472
rect 15929 12414 16068 12416
rect 15929 12411 15995 12414
rect 16062 12412 16068 12414
rect 16132 12412 16138 12476
rect 17726 12341 17786 12547
rect 22520 12520 23000 12550
rect 18045 12474 18111 12477
rect 18413 12474 18479 12477
rect 18045 12472 18479 12474
rect 18045 12416 18050 12472
rect 18106 12416 18418 12472
rect 18474 12416 18479 12472
rect 18045 12414 18479 12416
rect 18045 12411 18111 12414
rect 18413 12411 18479 12414
rect 3049 12338 3115 12341
rect 3693 12338 3759 12341
rect 10869 12338 10935 12341
rect 3049 12336 3759 12338
rect 3049 12280 3054 12336
rect 3110 12280 3698 12336
rect 3754 12280 3759 12336
rect 3049 12278 3759 12280
rect 3049 12275 3115 12278
rect 3693 12275 3759 12278
rect 8342 12336 10935 12338
rect 8342 12280 10874 12336
rect 10930 12280 10935 12336
rect 8342 12278 10935 12280
rect 0 12202 480 12232
rect 8342 12202 8402 12278
rect 10869 12275 10935 12278
rect 11053 12338 11119 12341
rect 11421 12338 11487 12341
rect 11053 12336 11487 12338
rect 11053 12280 11058 12336
rect 11114 12280 11426 12336
rect 11482 12280 11487 12336
rect 11053 12278 11487 12280
rect 11053 12275 11119 12278
rect 11421 12275 11487 12278
rect 11830 12276 11836 12340
rect 11900 12338 11906 12340
rect 12065 12338 12131 12341
rect 12893 12340 12959 12341
rect 12893 12338 12940 12340
rect 11900 12336 12131 12338
rect 11900 12280 12070 12336
rect 12126 12280 12131 12336
rect 11900 12278 12131 12280
rect 12848 12336 12940 12338
rect 12848 12280 12898 12336
rect 12848 12278 12940 12280
rect 11900 12276 11906 12278
rect 12065 12275 12131 12278
rect 12893 12276 12940 12278
rect 13004 12276 13010 12340
rect 13077 12338 13143 12341
rect 15326 12338 15332 12340
rect 13077 12336 15332 12338
rect 13077 12280 13082 12336
rect 13138 12280 15332 12336
rect 13077 12278 15332 12280
rect 12893 12275 12959 12276
rect 13077 12275 13143 12278
rect 15326 12276 15332 12278
rect 15396 12276 15402 12340
rect 17677 12336 17786 12341
rect 18137 12340 18203 12341
rect 18086 12338 18092 12340
rect 17677 12280 17682 12336
rect 17738 12280 17786 12336
rect 17677 12278 17786 12280
rect 18046 12278 18092 12338
rect 18156 12336 18203 12340
rect 18198 12280 18203 12336
rect 17677 12275 17743 12278
rect 18086 12276 18092 12278
rect 18156 12276 18203 12280
rect 18137 12275 18203 12276
rect 18781 12340 18847 12341
rect 18781 12336 18828 12340
rect 18892 12338 18898 12340
rect 18781 12280 18786 12336
rect 18781 12276 18828 12280
rect 18892 12278 18938 12338
rect 18892 12276 18898 12278
rect 18781 12275 18847 12276
rect 0 12142 8402 12202
rect 0 12112 480 12142
rect 8518 12140 8524 12204
rect 8588 12202 8594 12204
rect 13169 12202 13235 12205
rect 13670 12202 13676 12204
rect 8588 12142 12128 12202
rect 8588 12140 8594 12142
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 657 11930 723 11933
rect 6361 11930 6427 11933
rect 11053 11930 11119 11933
rect 657 11928 2698 11930
rect 657 11872 662 11928
rect 718 11872 2698 11928
rect 657 11870 2698 11872
rect 657 11867 723 11870
rect 2221 11794 2287 11797
rect 2446 11794 2452 11796
rect 2221 11792 2452 11794
rect 2221 11736 2226 11792
rect 2282 11736 2452 11792
rect 2221 11734 2452 11736
rect 2221 11731 2287 11734
rect 2446 11732 2452 11734
rect 2516 11732 2522 11796
rect 2638 11794 2698 11870
rect 6361 11928 11119 11930
rect 6361 11872 6366 11928
rect 6422 11872 11058 11928
rect 11114 11872 11119 11928
rect 6361 11870 11119 11872
rect 12068 11930 12128 12142
rect 13169 12200 13676 12202
rect 13169 12144 13174 12200
rect 13230 12144 13676 12200
rect 13169 12142 13676 12144
rect 13169 12139 13235 12142
rect 13670 12140 13676 12142
rect 13740 12140 13746 12204
rect 16113 12202 16179 12205
rect 16430 12202 16436 12204
rect 16113 12200 16436 12202
rect 16113 12144 16118 12200
rect 16174 12144 16436 12200
rect 16113 12142 16436 12144
rect 16113 12139 16179 12142
rect 16430 12140 16436 12142
rect 16500 12140 16506 12204
rect 20345 12202 20411 12205
rect 22520 12202 23000 12232
rect 20345 12200 23000 12202
rect 20345 12144 20350 12200
rect 20406 12144 23000 12200
rect 20345 12142 23000 12144
rect 20345 12139 20411 12142
rect 22520 12112 23000 12142
rect 16021 12068 16087 12069
rect 16021 12066 16068 12068
rect 15976 12064 16068 12066
rect 15976 12008 16026 12064
rect 15976 12006 16068 12008
rect 16021 12004 16068 12006
rect 16132 12004 16138 12068
rect 16021 12003 16087 12004
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 14825 11930 14891 11933
rect 12068 11928 14891 11930
rect 12068 11872 14830 11928
rect 14886 11872 14891 11928
rect 12068 11870 14891 11872
rect 6361 11867 6427 11870
rect 11053 11867 11119 11870
rect 14825 11867 14891 11870
rect 15009 11930 15075 11933
rect 15510 11930 15516 11932
rect 15009 11928 15516 11930
rect 15009 11872 15014 11928
rect 15070 11872 15516 11928
rect 15009 11870 15516 11872
rect 15009 11867 15075 11870
rect 15510 11868 15516 11870
rect 15580 11868 15586 11932
rect 8753 11794 8819 11797
rect 2638 11792 8819 11794
rect 2638 11736 8758 11792
rect 8814 11736 8819 11792
rect 2638 11734 8819 11736
rect 8753 11731 8819 11734
rect 9121 11794 9187 11797
rect 10409 11794 10475 11797
rect 9121 11792 10475 11794
rect 9121 11736 9126 11792
rect 9182 11736 10414 11792
rect 10470 11736 10475 11792
rect 9121 11734 10475 11736
rect 14828 11794 14888 11867
rect 14828 11734 17786 11794
rect 9121 11731 9187 11734
rect 10409 11731 10475 11734
rect 0 11658 480 11688
rect 1209 11658 1275 11661
rect 0 11656 1275 11658
rect 0 11600 1214 11656
rect 1270 11600 1275 11656
rect 0 11598 1275 11600
rect 0 11568 480 11598
rect 1209 11595 1275 11598
rect 3509 11658 3575 11661
rect 4245 11658 4311 11661
rect 3509 11656 4311 11658
rect 3509 11600 3514 11656
rect 3570 11600 4250 11656
rect 4306 11600 4311 11656
rect 3509 11598 4311 11600
rect 3509 11595 3575 11598
rect 4245 11595 4311 11598
rect 9581 11656 9647 11661
rect 9581 11600 9586 11656
rect 9642 11600 9647 11656
rect 9581 11595 9647 11600
rect 10501 11658 10567 11661
rect 10501 11656 16866 11658
rect 10501 11600 10506 11656
rect 10562 11600 16866 11656
rect 10501 11598 16866 11600
rect 10501 11595 10567 11598
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 9584 11389 9644 11595
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 9581 11384 9647 11389
rect 9581 11328 9586 11384
rect 9642 11328 9647 11384
rect 9581 11323 9647 11328
rect 11605 11386 11671 11389
rect 15377 11386 15443 11389
rect 16062 11386 16068 11388
rect 11605 11384 14658 11386
rect 11605 11328 11610 11384
rect 11666 11328 14658 11384
rect 11605 11326 14658 11328
rect 11605 11323 11671 11326
rect 4705 11250 4771 11253
rect 9765 11250 9831 11253
rect 4705 11248 9831 11250
rect 4705 11192 4710 11248
rect 4766 11192 9770 11248
rect 9826 11192 9831 11248
rect 4705 11190 9831 11192
rect 14598 11250 14658 11326
rect 15377 11384 16068 11386
rect 15377 11328 15382 11384
rect 15438 11328 16068 11384
rect 15377 11326 16068 11328
rect 15377 11323 15443 11326
rect 16062 11324 16068 11326
rect 16132 11324 16138 11388
rect 14598 11190 16682 11250
rect 4705 11187 4771 11190
rect 9765 11187 9831 11190
rect 0 11114 480 11144
rect 16622 11117 16682 11190
rect 4521 11114 4587 11117
rect 0 11112 4587 11114
rect 0 11056 4526 11112
rect 4582 11056 4587 11112
rect 0 11054 4587 11056
rect 0 11024 480 11054
rect 4521 11051 4587 11054
rect 4705 11114 4771 11117
rect 5390 11114 5396 11116
rect 4705 11112 5396 11114
rect 4705 11056 4710 11112
rect 4766 11056 5396 11112
rect 4705 11054 5396 11056
rect 4705 11051 4771 11054
rect 5390 11052 5396 11054
rect 5460 11052 5466 11116
rect 10225 11114 10291 11117
rect 14590 11114 14596 11116
rect 10225 11112 14596 11114
rect 10225 11056 10230 11112
rect 10286 11056 14596 11112
rect 10225 11054 14596 11056
rect 10225 11051 10291 11054
rect 14590 11052 14596 11054
rect 14660 11052 14666 11116
rect 16622 11112 16731 11117
rect 16622 11056 16670 11112
rect 16726 11056 16731 11112
rect 16622 11054 16731 11056
rect 16806 11114 16866 11598
rect 17726 11525 17786 11734
rect 17953 11792 18019 11797
rect 17953 11736 17958 11792
rect 18014 11736 18019 11792
rect 17953 11731 18019 11736
rect 17956 11658 18016 11731
rect 22520 11658 23000 11688
rect 17956 11598 23000 11658
rect 22520 11568 23000 11598
rect 17726 11520 17835 11525
rect 17726 11464 17774 11520
rect 17830 11464 17835 11520
rect 17726 11462 17835 11464
rect 17769 11459 17835 11462
rect 17033 11388 17099 11389
rect 16982 11324 16988 11388
rect 17052 11386 17099 11388
rect 17052 11384 17144 11386
rect 17094 11328 17144 11384
rect 17052 11326 17144 11328
rect 17052 11324 17099 11326
rect 17033 11323 17099 11324
rect 19006 11114 19012 11116
rect 16806 11054 19012 11114
rect 16665 11051 16731 11054
rect 19006 11052 19012 11054
rect 19076 11114 19082 11116
rect 22520 11114 23000 11144
rect 19076 11054 23000 11114
rect 19076 11052 19082 11054
rect 22520 11024 23000 11054
rect 12249 10978 12315 10981
rect 17861 10978 17927 10981
rect 12249 10976 17927 10978
rect 12249 10920 12254 10976
rect 12310 10920 17866 10976
rect 17922 10920 17927 10976
rect 12249 10918 17927 10920
rect 12249 10915 12315 10918
rect 17861 10915 17927 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 15377 10842 15443 10845
rect 15561 10842 15627 10845
rect 15377 10840 15627 10842
rect 15377 10784 15382 10840
rect 15438 10784 15566 10840
rect 15622 10784 15627 10840
rect 15377 10782 15627 10784
rect 15377 10779 15443 10782
rect 15561 10779 15627 10782
rect 0 10706 480 10736
rect 1025 10706 1091 10709
rect 0 10704 1091 10706
rect 0 10648 1030 10704
rect 1086 10648 1091 10704
rect 0 10646 1091 10648
rect 0 10616 480 10646
rect 1025 10643 1091 10646
rect 3693 10706 3759 10709
rect 3918 10706 3924 10708
rect 3693 10704 3924 10706
rect 3693 10648 3698 10704
rect 3754 10648 3924 10704
rect 3693 10646 3924 10648
rect 3693 10643 3759 10646
rect 3918 10644 3924 10646
rect 3988 10644 3994 10708
rect 5574 10644 5580 10708
rect 5644 10706 5650 10708
rect 5717 10706 5783 10709
rect 5644 10704 5783 10706
rect 5644 10648 5722 10704
rect 5778 10648 5783 10704
rect 5644 10646 5783 10648
rect 5644 10644 5650 10646
rect 5717 10643 5783 10646
rect 13721 10706 13787 10709
rect 14825 10706 14891 10709
rect 13721 10704 14891 10706
rect 13721 10648 13726 10704
rect 13782 10648 14830 10704
rect 14886 10648 14891 10704
rect 13721 10646 14891 10648
rect 13721 10643 13787 10646
rect 14825 10643 14891 10646
rect 19609 10706 19675 10709
rect 22520 10706 23000 10736
rect 19609 10704 23000 10706
rect 19609 10648 19614 10704
rect 19670 10648 23000 10704
rect 19609 10646 23000 10648
rect 19609 10643 19675 10646
rect 22520 10616 23000 10646
rect 3693 10570 3759 10573
rect 4102 10570 4108 10572
rect 3693 10568 4108 10570
rect 3693 10512 3698 10568
rect 3754 10512 4108 10568
rect 3693 10510 4108 10512
rect 3693 10507 3759 10510
rect 4102 10508 4108 10510
rect 4172 10508 4178 10572
rect 14457 10570 14523 10573
rect 15745 10570 15811 10573
rect 14457 10568 15811 10570
rect 14457 10512 14462 10568
rect 14518 10512 15750 10568
rect 15806 10512 15811 10568
rect 14457 10510 15811 10512
rect 14457 10507 14523 10510
rect 15745 10507 15811 10510
rect 15561 10434 15627 10437
rect 15694 10434 15700 10436
rect 15561 10432 15700 10434
rect 15561 10376 15566 10432
rect 15622 10376 15700 10432
rect 15561 10374 15700 10376
rect 15561 10371 15627 10374
rect 15694 10372 15700 10374
rect 15764 10372 15770 10436
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 3693 10298 3759 10301
rect 13721 10300 13787 10301
rect 3693 10296 3986 10298
rect 3693 10240 3698 10296
rect 3754 10240 3986 10296
rect 3693 10238 3986 10240
rect 3693 10235 3759 10238
rect 0 10162 480 10192
rect 565 10162 631 10165
rect 0 10160 631 10162
rect 0 10104 570 10160
rect 626 10104 631 10160
rect 0 10102 631 10104
rect 0 10072 480 10102
rect 565 10099 631 10102
rect 2865 10162 2931 10165
rect 2865 10160 3618 10162
rect 2865 10104 2870 10160
rect 2926 10104 3618 10160
rect 2865 10102 3618 10104
rect 2865 10099 2931 10102
rect 0 9618 480 9648
rect 3558 9618 3618 10102
rect 3693 9618 3759 9621
rect 0 9558 1410 9618
rect 3558 9616 3759 9618
rect 3558 9560 3698 9616
rect 3754 9560 3759 9616
rect 3558 9558 3759 9560
rect 0 9528 480 9558
rect 1350 9346 1410 9558
rect 3693 9555 3759 9558
rect 3926 9485 3986 10238
rect 13670 10236 13676 10300
rect 13740 10298 13787 10300
rect 13740 10296 13832 10298
rect 13782 10240 13832 10296
rect 13740 10238 13832 10240
rect 13740 10236 13787 10238
rect 13721 10235 13787 10236
rect 12065 10162 12131 10165
rect 12433 10162 12499 10165
rect 12065 10160 12499 10162
rect 12065 10104 12070 10160
rect 12126 10104 12438 10160
rect 12494 10104 12499 10160
rect 12065 10102 12499 10104
rect 12065 10099 12131 10102
rect 12433 10099 12499 10102
rect 18229 10162 18295 10165
rect 22520 10162 23000 10192
rect 18229 10160 23000 10162
rect 18229 10104 18234 10160
rect 18290 10104 23000 10160
rect 18229 10102 23000 10104
rect 18229 10099 18295 10102
rect 22520 10072 23000 10102
rect 4521 10026 4587 10029
rect 7230 10026 7236 10028
rect 4521 10024 7236 10026
rect 4521 9968 4526 10024
rect 4582 9968 7236 10024
rect 4521 9966 7236 9968
rect 4521 9963 4587 9966
rect 7230 9964 7236 9966
rect 7300 9964 7306 10028
rect 7598 9964 7604 10028
rect 7668 10026 7674 10028
rect 13118 10026 13124 10028
rect 7668 9966 13124 10026
rect 7668 9964 7674 9966
rect 13118 9964 13124 9966
rect 13188 9964 13194 10028
rect 15101 10026 15167 10029
rect 15510 10026 15516 10028
rect 15101 10024 15516 10026
rect 15101 9968 15106 10024
rect 15162 9968 15516 10024
rect 15101 9966 15516 9968
rect 15101 9963 15167 9966
rect 15510 9964 15516 9966
rect 15580 9964 15586 10028
rect 20529 10026 20595 10029
rect 20486 10024 20595 10026
rect 20486 9968 20534 10024
rect 20590 9968 20595 10024
rect 20486 9963 20595 9968
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 20486 9757 20546 9963
rect 8385 9754 8451 9757
rect 8342 9752 8451 9754
rect 8342 9696 8390 9752
rect 8446 9696 8451 9752
rect 8342 9691 8451 9696
rect 20486 9752 20595 9757
rect 20486 9696 20534 9752
rect 20590 9696 20595 9752
rect 20486 9694 20595 9696
rect 20529 9691 20595 9694
rect 8342 9618 8402 9691
rect 8477 9618 8543 9621
rect 8342 9616 8543 9618
rect 8342 9560 8482 9616
rect 8538 9560 8543 9616
rect 8342 9558 8543 9560
rect 8477 9555 8543 9558
rect 10542 9556 10548 9620
rect 10612 9618 10618 9620
rect 16757 9618 16823 9621
rect 10612 9616 16823 9618
rect 10612 9560 16762 9616
rect 16818 9560 16823 9616
rect 10612 9558 16823 9560
rect 10612 9556 10618 9558
rect 16757 9555 16823 9558
rect 16982 9556 16988 9620
rect 17052 9618 17058 9620
rect 22520 9618 23000 9648
rect 17052 9558 23000 9618
rect 17052 9556 17058 9558
rect 22520 9528 23000 9558
rect 2221 9482 2287 9485
rect 2773 9482 2839 9485
rect 2221 9480 2839 9482
rect 2221 9424 2226 9480
rect 2282 9424 2778 9480
rect 2834 9424 2839 9480
rect 2221 9422 2839 9424
rect 3926 9480 4035 9485
rect 3926 9424 3974 9480
rect 4030 9424 4035 9480
rect 3926 9422 4035 9424
rect 2221 9419 2287 9422
rect 2773 9419 2839 9422
rect 3969 9419 4035 9422
rect 14038 9420 14044 9484
rect 14108 9482 14114 9484
rect 15101 9482 15167 9485
rect 14108 9480 15167 9482
rect 14108 9424 15106 9480
rect 15162 9424 15167 9480
rect 14108 9422 15167 9424
rect 14108 9420 14114 9422
rect 15101 9419 15167 9422
rect 15377 9482 15443 9485
rect 15510 9482 15516 9484
rect 15377 9480 15516 9482
rect 15377 9424 15382 9480
rect 15438 9424 15516 9480
rect 15377 9422 15516 9424
rect 15377 9419 15443 9422
rect 15510 9420 15516 9422
rect 15580 9420 15586 9484
rect 4061 9346 4127 9349
rect 1350 9344 4127 9346
rect 1350 9288 4066 9344
rect 4122 9288 4127 9344
rect 1350 9286 4127 9288
rect 4061 9283 4127 9286
rect 11605 9346 11671 9349
rect 13302 9346 13308 9348
rect 11605 9344 13308 9346
rect 11605 9288 11610 9344
rect 11666 9288 13308 9344
rect 11605 9286 13308 9288
rect 11605 9283 11671 9286
rect 13302 9284 13308 9286
rect 13372 9284 13378 9348
rect 17902 9284 17908 9348
rect 17972 9346 17978 9348
rect 18229 9346 18295 9349
rect 17972 9344 18295 9346
rect 17972 9288 18234 9344
rect 18290 9288 18295 9344
rect 17972 9286 18295 9288
rect 17972 9284 17978 9286
rect 18229 9283 18295 9286
rect 7874 9280 8194 9281
rect 0 9210 480 9240
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 0 9150 4906 9210
rect 0 9120 480 9150
rect 4846 9074 4906 9150
rect 11094 9148 11100 9212
rect 11164 9210 11170 9212
rect 11605 9210 11671 9213
rect 11164 9208 11671 9210
rect 11164 9152 11610 9208
rect 11666 9152 11671 9208
rect 11164 9150 11671 9152
rect 11164 9148 11170 9150
rect 11102 9074 11162 9148
rect 11605 9147 11671 9150
rect 12065 9210 12131 9213
rect 16798 9210 16804 9212
rect 12065 9208 14704 9210
rect 12065 9152 12070 9208
rect 12126 9152 14704 9208
rect 12065 9150 14704 9152
rect 12065 9147 12131 9150
rect 4846 9014 11162 9074
rect 11513 9074 11579 9077
rect 13813 9076 13879 9077
rect 12566 9074 12572 9076
rect 11513 9072 12572 9074
rect 11513 9016 11518 9072
rect 11574 9016 12572 9072
rect 11513 9014 12572 9016
rect 11513 9011 11579 9014
rect 12566 9012 12572 9014
rect 12636 9012 12642 9076
rect 13813 9072 13860 9076
rect 13924 9074 13930 9076
rect 14644 9074 14704 9150
rect 15334 9150 16804 9210
rect 15334 9074 15394 9150
rect 16798 9148 16804 9150
rect 16868 9210 16874 9212
rect 22520 9210 23000 9240
rect 16868 9150 23000 9210
rect 16868 9148 16874 9150
rect 22520 9120 23000 9150
rect 13813 9016 13818 9072
rect 13813 9012 13860 9016
rect 13924 9014 13970 9074
rect 14644 9014 15394 9074
rect 13924 9012 13930 9014
rect 13813 9011 13879 9012
rect 4102 8876 4108 8940
rect 4172 8938 4178 8940
rect 8569 8938 8635 8941
rect 4172 8936 8635 8938
rect 4172 8880 8574 8936
rect 8630 8880 8635 8936
rect 4172 8878 8635 8880
rect 4172 8876 4178 8878
rect 8569 8875 8635 8878
rect 12433 8938 12499 8941
rect 18229 8938 18295 8941
rect 12433 8936 18295 8938
rect 12433 8880 12438 8936
rect 12494 8880 18234 8936
rect 18290 8880 18295 8936
rect 12433 8878 18295 8880
rect 12433 8875 12499 8878
rect 18229 8875 18295 8878
rect 7189 8804 7255 8805
rect 7189 8802 7236 8804
rect 7144 8800 7236 8802
rect 7144 8744 7194 8800
rect 7144 8742 7236 8744
rect 7189 8740 7236 8742
rect 7300 8740 7306 8804
rect 7189 8739 7255 8740
rect 4409 8736 4729 8737
rect 0 8666 480 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 3969 8666 4035 8669
rect 0 8664 4035 8666
rect 0 8608 3974 8664
rect 4030 8608 4035 8664
rect 0 8606 4035 8608
rect 0 8576 480 8606
rect 3969 8603 4035 8606
rect 7598 8604 7604 8668
rect 7668 8666 7674 8668
rect 7741 8666 7807 8669
rect 7668 8664 7807 8666
rect 7668 8608 7746 8664
rect 7802 8608 7807 8664
rect 7668 8606 7807 8608
rect 7668 8604 7674 8606
rect 7741 8603 7807 8606
rect 18781 8666 18847 8669
rect 22520 8666 23000 8696
rect 18781 8664 23000 8666
rect 18781 8608 18786 8664
rect 18842 8608 23000 8664
rect 18781 8606 23000 8608
rect 18781 8603 18847 8606
rect 22520 8576 23000 8606
rect 10225 8530 10291 8533
rect 16481 8530 16547 8533
rect 10225 8528 16547 8530
rect 10225 8472 10230 8528
rect 10286 8472 16486 8528
rect 16542 8472 16547 8528
rect 10225 8470 16547 8472
rect 10225 8467 10291 8470
rect 16481 8467 16547 8470
rect 8753 8394 8819 8397
rect 15653 8396 15719 8397
rect 16113 8396 16179 8397
rect 15653 8394 15700 8396
rect 8753 8392 15700 8394
rect 15764 8394 15770 8396
rect 8753 8336 8758 8392
rect 8814 8336 15658 8392
rect 8753 8334 15700 8336
rect 8753 8331 8819 8334
rect 15653 8332 15700 8334
rect 15764 8334 15846 8394
rect 15764 8332 15770 8334
rect 16062 8332 16068 8396
rect 16132 8394 16179 8396
rect 16132 8392 16224 8394
rect 16174 8336 16224 8392
rect 16132 8334 16224 8336
rect 16132 8332 16179 8334
rect 15653 8331 15719 8332
rect 16113 8331 16179 8332
rect 7874 8192 8194 8193
rect 0 8122 480 8152
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 4061 8122 4127 8125
rect 0 8120 4127 8122
rect 0 8064 4066 8120
rect 4122 8064 4127 8120
rect 0 8062 4127 8064
rect 0 8032 480 8062
rect 4061 8059 4127 8062
rect 15326 8060 15332 8124
rect 15396 8122 15402 8124
rect 22520 8122 23000 8152
rect 15396 8062 23000 8122
rect 15396 8060 15402 8062
rect 22520 8032 23000 8062
rect 10777 7986 10843 7989
rect 18822 7986 18828 7988
rect 10777 7984 18828 7986
rect 10777 7928 10782 7984
rect 10838 7928 18828 7984
rect 10777 7926 18828 7928
rect 10777 7923 10843 7926
rect 18822 7924 18828 7926
rect 18892 7924 18898 7988
rect 6637 7850 6703 7853
rect 4156 7848 6703 7850
rect 4156 7792 6642 7848
rect 6698 7792 6703 7848
rect 4156 7790 6703 7792
rect 0 7714 480 7744
rect 4156 7714 4216 7790
rect 6637 7787 6703 7790
rect 11697 7850 11763 7853
rect 17217 7850 17283 7853
rect 11697 7848 17283 7850
rect 11697 7792 11702 7848
rect 11758 7792 17222 7848
rect 17278 7792 17283 7848
rect 11697 7790 17283 7792
rect 11697 7787 11763 7790
rect 17217 7787 17283 7790
rect 0 7654 4216 7714
rect 19241 7714 19307 7717
rect 22520 7714 23000 7744
rect 19241 7712 23000 7714
rect 19241 7656 19246 7712
rect 19302 7656 23000 7712
rect 19241 7654 23000 7656
rect 0 7624 480 7654
rect 19241 7651 19307 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 22520 7624 23000 7654
rect 18270 7583 18590 7584
rect 3918 7380 3924 7444
rect 3988 7442 3994 7444
rect 4705 7442 4771 7445
rect 3988 7440 4771 7442
rect 3988 7384 4710 7440
rect 4766 7384 4771 7440
rect 3988 7382 4771 7384
rect 3988 7380 3994 7382
rect 4705 7379 4771 7382
rect 5206 7380 5212 7444
rect 5276 7442 5282 7444
rect 7833 7442 7899 7445
rect 5276 7440 7899 7442
rect 5276 7384 7838 7440
rect 7894 7384 7899 7440
rect 5276 7382 7899 7384
rect 5276 7380 5282 7382
rect 7833 7379 7899 7382
rect 16389 7444 16455 7445
rect 16389 7440 16436 7444
rect 16500 7442 16506 7444
rect 18045 7442 18111 7445
rect 16389 7384 16394 7440
rect 16389 7380 16436 7384
rect 16500 7382 16546 7442
rect 18045 7440 18154 7442
rect 18045 7384 18050 7440
rect 18106 7384 18154 7440
rect 16500 7380 16506 7382
rect 16389 7379 16455 7380
rect 18045 7379 18154 7384
rect 7189 7306 7255 7309
rect 8201 7306 8267 7309
rect 9673 7308 9739 7309
rect 7189 7304 7482 7306
rect 7189 7248 7194 7304
rect 7250 7248 7482 7304
rect 7189 7246 7482 7248
rect 7189 7243 7255 7246
rect 0 7170 480 7200
rect 4061 7170 4127 7173
rect 0 7168 4127 7170
rect 0 7112 4066 7168
rect 4122 7112 4127 7168
rect 0 7110 4127 7112
rect 0 7080 480 7110
rect 4061 7107 4127 7110
rect 7422 6765 7482 7246
rect 7606 7304 8267 7306
rect 7606 7248 8206 7304
rect 8262 7248 8267 7304
rect 7606 7246 8267 7248
rect 7606 6898 7666 7246
rect 8201 7243 8267 7246
rect 9622 7244 9628 7308
rect 9692 7306 9739 7308
rect 14917 7306 14983 7309
rect 9692 7304 9784 7306
rect 9734 7248 9784 7304
rect 9692 7246 9784 7248
rect 14598 7304 14983 7306
rect 14598 7248 14922 7304
rect 14978 7248 14983 7304
rect 14598 7246 14983 7248
rect 9692 7244 9739 7246
rect 9673 7243 9739 7244
rect 9765 7172 9831 7173
rect 9765 7170 9812 7172
rect 9720 7168 9812 7170
rect 9720 7112 9770 7168
rect 9720 7110 9812 7112
rect 9765 7108 9812 7110
rect 9876 7108 9882 7172
rect 9765 7107 9831 7108
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14598 7037 14658 7246
rect 14917 7243 14983 7246
rect 16573 7306 16639 7309
rect 16941 7306 17007 7309
rect 17125 7306 17191 7309
rect 16573 7304 17191 7306
rect 16573 7248 16578 7304
rect 16634 7248 16946 7304
rect 17002 7248 17130 7304
rect 17186 7248 17191 7304
rect 16573 7246 17191 7248
rect 16573 7243 16639 7246
rect 16941 7243 17007 7246
rect 17125 7243 17191 7246
rect 18094 7173 18154 7379
rect 18873 7308 18939 7309
rect 18822 7306 18828 7308
rect 18746 7246 18828 7306
rect 18892 7306 18939 7308
rect 19742 7306 19748 7308
rect 18892 7304 19748 7306
rect 18934 7248 19748 7304
rect 18822 7244 18828 7246
rect 18892 7246 19748 7248
rect 18892 7244 18939 7246
rect 19742 7244 19748 7246
rect 19812 7244 19818 7308
rect 18873 7243 18939 7244
rect 18045 7168 18154 7173
rect 18045 7112 18050 7168
rect 18106 7112 18154 7168
rect 18045 7110 18154 7112
rect 20621 7170 20687 7173
rect 22520 7170 23000 7200
rect 20621 7168 23000 7170
rect 20621 7112 20626 7168
rect 20682 7112 23000 7168
rect 20621 7110 23000 7112
rect 18045 7107 18111 7110
rect 20621 7107 20687 7110
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 22520 7080 23000 7110
rect 14805 7039 15125 7040
rect 9581 7034 9647 7037
rect 13353 7034 13419 7037
rect 9581 7032 13419 7034
rect 9581 6976 9586 7032
rect 9642 6976 13358 7032
rect 13414 6976 13419 7032
rect 9581 6974 13419 6976
rect 14598 7032 14707 7037
rect 14598 6976 14646 7032
rect 14702 6976 14707 7032
rect 14598 6974 14707 6976
rect 9581 6971 9647 6974
rect 13353 6971 13419 6974
rect 14641 6971 14707 6974
rect 8109 6898 8175 6901
rect 7606 6896 8175 6898
rect 7606 6840 8114 6896
rect 8170 6840 8175 6896
rect 7606 6838 8175 6840
rect 8109 6835 8175 6838
rect 8385 6898 8451 6901
rect 17493 6898 17559 6901
rect 8385 6896 17559 6898
rect 8385 6840 8390 6896
rect 8446 6840 17498 6896
rect 17554 6840 17559 6896
rect 8385 6838 17559 6840
rect 8385 6835 8451 6838
rect 17493 6835 17559 6838
rect 7422 6760 7531 6765
rect 7422 6704 7470 6760
rect 7526 6704 7531 6760
rect 7422 6702 7531 6704
rect 7465 6699 7531 6702
rect 8385 6762 8451 6765
rect 10685 6762 10751 6765
rect 19149 6762 19215 6765
rect 8385 6760 19215 6762
rect 8385 6704 8390 6760
rect 8446 6704 10690 6760
rect 10746 6704 19154 6760
rect 19210 6704 19215 6760
rect 8385 6702 19215 6704
rect 8385 6699 8451 6702
rect 10685 6699 10751 6702
rect 19149 6699 19215 6702
rect 0 6626 480 6656
rect 4061 6626 4127 6629
rect 0 6624 4127 6626
rect 0 6568 4066 6624
rect 4122 6568 4127 6624
rect 0 6566 4127 6568
rect 0 6536 480 6566
rect 4061 6563 4127 6566
rect 12801 6626 12867 6629
rect 15837 6626 15903 6629
rect 12801 6624 15903 6626
rect 12801 6568 12806 6624
rect 12862 6568 15842 6624
rect 15898 6568 15903 6624
rect 12801 6566 15903 6568
rect 12801 6563 12867 6566
rect 15837 6563 15903 6566
rect 19241 6626 19307 6629
rect 22520 6626 23000 6656
rect 19241 6624 23000 6626
rect 19241 6568 19246 6624
rect 19302 6568 23000 6624
rect 19241 6566 23000 6568
rect 19241 6563 19307 6566
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 22520 6536 23000 6566
rect 18270 6495 18590 6496
rect 2405 6354 2471 6357
rect 9305 6354 9371 6357
rect 2405 6352 9371 6354
rect 2405 6296 2410 6352
rect 2466 6296 9310 6352
rect 9366 6296 9371 6352
rect 2405 6294 9371 6296
rect 2405 6291 2471 6294
rect 9305 6291 9371 6294
rect 12801 6354 12867 6357
rect 15326 6354 15332 6356
rect 12801 6352 15332 6354
rect 12801 6296 12806 6352
rect 12862 6296 15332 6352
rect 12801 6294 15332 6296
rect 12801 6291 12867 6294
rect 15326 6292 15332 6294
rect 15396 6292 15402 6356
rect 15745 6352 15811 6357
rect 15745 6296 15750 6352
rect 15806 6296 15811 6352
rect 15745 6291 15811 6296
rect 0 6218 480 6248
rect 3785 6218 3851 6221
rect 0 6216 3851 6218
rect 0 6160 3790 6216
rect 3846 6160 3851 6216
rect 0 6158 3851 6160
rect 0 6128 480 6158
rect 3785 6155 3851 6158
rect 10869 6218 10935 6221
rect 15748 6218 15808 6291
rect 10869 6216 15808 6218
rect 10869 6160 10874 6216
rect 10930 6160 15808 6216
rect 10869 6158 15808 6160
rect 18873 6218 18939 6221
rect 22520 6218 23000 6248
rect 18873 6216 23000 6218
rect 18873 6160 18878 6216
rect 18934 6160 23000 6216
rect 18873 6158 23000 6160
rect 10869 6155 10935 6158
rect 18873 6155 18939 6158
rect 22520 6128 23000 6158
rect 9581 6082 9647 6085
rect 13813 6082 13879 6085
rect 14038 6082 14044 6084
rect 9581 6080 14044 6082
rect 9581 6024 9586 6080
rect 9642 6024 13818 6080
rect 13874 6024 14044 6080
rect 9581 6022 14044 6024
rect 9581 6019 9647 6022
rect 13813 6019 13879 6022
rect 14038 6020 14044 6022
rect 14108 6020 14114 6084
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 9806 5884 9812 5948
rect 9876 5946 9882 5948
rect 9949 5946 10015 5949
rect 9876 5944 10015 5946
rect 9876 5888 9954 5944
rect 10010 5888 10015 5944
rect 9876 5886 10015 5888
rect 9876 5884 9882 5886
rect 9949 5883 10015 5886
rect 11145 5946 11211 5949
rect 11513 5946 11579 5949
rect 11145 5944 11579 5946
rect 11145 5888 11150 5944
rect 11206 5888 11518 5944
rect 11574 5888 11579 5944
rect 11145 5886 11579 5888
rect 11145 5883 11211 5886
rect 11513 5883 11579 5886
rect 13302 5884 13308 5948
rect 13372 5946 13378 5948
rect 13537 5946 13603 5949
rect 13813 5948 13879 5949
rect 14641 5948 14707 5949
rect 13813 5946 13860 5948
rect 13372 5944 13603 5946
rect 13372 5888 13542 5944
rect 13598 5888 13603 5944
rect 13372 5886 13603 5888
rect 13768 5944 13860 5946
rect 13768 5888 13818 5944
rect 13768 5886 13860 5888
rect 13372 5884 13378 5886
rect 13537 5883 13603 5886
rect 13813 5884 13860 5886
rect 13924 5884 13930 5948
rect 14590 5946 14596 5948
rect 14550 5886 14596 5946
rect 14660 5944 14707 5948
rect 14702 5888 14707 5944
rect 14590 5884 14596 5886
rect 14660 5884 14707 5888
rect 13813 5883 13879 5884
rect 14641 5883 14707 5884
rect 2868 5750 4906 5810
rect 0 5674 480 5704
rect 2868 5674 2928 5750
rect 0 5614 2928 5674
rect 3049 5674 3115 5677
rect 3366 5674 3372 5676
rect 3049 5672 3372 5674
rect 3049 5616 3054 5672
rect 3110 5616 3372 5672
rect 3049 5614 3372 5616
rect 0 5584 480 5614
rect 3049 5611 3115 5614
rect 3366 5612 3372 5614
rect 3436 5612 3442 5676
rect 4846 5538 4906 5750
rect 15510 5748 15516 5812
rect 15580 5810 15586 5812
rect 19241 5810 19307 5813
rect 15580 5808 19307 5810
rect 15580 5752 19246 5808
rect 19302 5752 19307 5808
rect 15580 5750 19307 5752
rect 15580 5748 15586 5750
rect 19241 5747 19307 5750
rect 8661 5674 8727 5677
rect 16614 5674 16620 5676
rect 8661 5672 16620 5674
rect 8661 5616 8666 5672
rect 8722 5616 16620 5672
rect 8661 5614 16620 5616
rect 8661 5611 8727 5614
rect 16614 5612 16620 5614
rect 16684 5612 16690 5676
rect 19149 5674 19215 5677
rect 22520 5674 23000 5704
rect 19149 5672 23000 5674
rect 19149 5616 19154 5672
rect 19210 5616 23000 5672
rect 19149 5614 23000 5616
rect 19149 5611 19215 5614
rect 22520 5584 23000 5614
rect 9121 5538 9187 5541
rect 4846 5536 9187 5538
rect 4846 5480 9126 5536
rect 9182 5480 9187 5536
rect 4846 5478 9187 5480
rect 9121 5475 9187 5478
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 12433 5402 12499 5405
rect 14641 5402 14707 5405
rect 16982 5402 16988 5404
rect 12433 5400 16988 5402
rect 12433 5344 12438 5400
rect 12494 5344 14646 5400
rect 14702 5344 16988 5400
rect 12433 5342 16988 5344
rect 12433 5339 12499 5342
rect 14641 5339 14707 5342
rect 16982 5340 16988 5342
rect 17052 5340 17058 5404
rect 2865 5266 2931 5269
rect 5441 5268 5507 5269
rect 5206 5266 5212 5268
rect 2865 5264 5212 5266
rect 2865 5208 2870 5264
rect 2926 5208 5212 5264
rect 2865 5206 5212 5208
rect 2865 5203 2931 5206
rect 5206 5204 5212 5206
rect 5276 5204 5282 5268
rect 5390 5266 5396 5268
rect 5350 5206 5396 5266
rect 5460 5264 5507 5268
rect 5502 5208 5507 5264
rect 5390 5204 5396 5206
rect 5460 5204 5507 5208
rect 5441 5203 5507 5204
rect 10225 5266 10291 5269
rect 15285 5266 15351 5269
rect 10225 5264 15351 5266
rect 10225 5208 10230 5264
rect 10286 5208 15290 5264
rect 15346 5208 15351 5264
rect 10225 5206 15351 5208
rect 10225 5203 10291 5206
rect 15285 5203 15351 5206
rect 15653 5266 15719 5269
rect 17902 5266 17908 5268
rect 15653 5264 17908 5266
rect 15653 5208 15658 5264
rect 15714 5208 17908 5264
rect 15653 5206 17908 5208
rect 15653 5203 15719 5206
rect 17902 5204 17908 5206
rect 17972 5204 17978 5268
rect 0 5130 480 5160
rect 3785 5130 3851 5133
rect 4153 5132 4219 5133
rect 4102 5130 4108 5132
rect 0 5128 3851 5130
rect 0 5072 3790 5128
rect 3846 5072 3851 5128
rect 0 5070 3851 5072
rect 4062 5070 4108 5130
rect 4172 5128 4219 5132
rect 4214 5072 4219 5128
rect 0 5040 480 5070
rect 3785 5067 3851 5070
rect 4102 5068 4108 5070
rect 4172 5068 4219 5072
rect 4153 5067 4219 5068
rect 10409 5130 10475 5133
rect 11697 5130 11763 5133
rect 16389 5130 16455 5133
rect 17585 5130 17651 5133
rect 10409 5128 11763 5130
rect 10409 5072 10414 5128
rect 10470 5072 11702 5128
rect 11758 5072 11763 5128
rect 10409 5070 11763 5072
rect 10409 5067 10475 5070
rect 11697 5067 11763 5070
rect 14644 5128 17651 5130
rect 14644 5072 16394 5128
rect 16450 5072 17590 5128
rect 17646 5072 17651 5128
rect 14644 5070 17651 5072
rect 10317 4994 10383 4997
rect 10542 4994 10548 4996
rect 10317 4992 10548 4994
rect 10317 4936 10322 4992
rect 10378 4936 10548 4992
rect 10317 4934 10548 4936
rect 10317 4931 10383 4934
rect 10542 4932 10548 4934
rect 10612 4932 10618 4996
rect 10777 4994 10843 4997
rect 14644 4994 14704 5070
rect 16389 5067 16455 5070
rect 17585 5067 17651 5070
rect 22369 5130 22435 5133
rect 22520 5130 23000 5160
rect 22369 5128 23000 5130
rect 22369 5072 22374 5128
rect 22430 5072 23000 5128
rect 22369 5070 23000 5072
rect 22369 5067 22435 5070
rect 22520 5040 23000 5070
rect 10777 4992 14704 4994
rect 10777 4936 10782 4992
rect 10838 4936 14704 4992
rect 10777 4934 14704 4936
rect 10777 4931 10843 4934
rect 17902 4932 17908 4996
rect 17972 4994 17978 4996
rect 22369 4994 22435 4997
rect 17972 4992 22435 4994
rect 17972 4936 22374 4992
rect 22430 4936 22435 4992
rect 17972 4934 22435 4936
rect 17972 4932 17978 4934
rect 22369 4931 22435 4934
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 9765 4858 9831 4861
rect 9765 4856 14704 4858
rect 9765 4800 9770 4856
rect 9826 4800 14704 4856
rect 9765 4798 14704 4800
rect 9765 4795 9831 4798
rect 0 4722 480 4752
rect 2865 4722 2931 4725
rect 0 4720 2931 4722
rect 0 4664 2870 4720
rect 2926 4664 2931 4720
rect 0 4662 2931 4664
rect 0 4632 480 4662
rect 2865 4659 2931 4662
rect 8293 4722 8359 4725
rect 11237 4722 11303 4725
rect 14273 4722 14339 4725
rect 8293 4720 14339 4722
rect 8293 4664 8298 4720
rect 8354 4664 11242 4720
rect 11298 4664 14278 4720
rect 14334 4664 14339 4720
rect 8293 4662 14339 4664
rect 14644 4722 14704 4798
rect 16849 4722 16915 4725
rect 14644 4720 16915 4722
rect 14644 4664 16854 4720
rect 16910 4664 16915 4720
rect 14644 4662 16915 4664
rect 8293 4659 8359 4662
rect 11237 4659 11303 4662
rect 14273 4659 14339 4662
rect 16849 4659 16915 4662
rect 17769 4722 17835 4725
rect 22520 4722 23000 4752
rect 17769 4720 23000 4722
rect 17769 4664 17774 4720
rect 17830 4664 23000 4720
rect 17769 4662 23000 4664
rect 17769 4659 17835 4662
rect 22520 4632 23000 4662
rect 10317 4586 10383 4589
rect 12617 4586 12683 4589
rect 16389 4586 16455 4589
rect 18873 4586 18939 4589
rect 10317 4584 12450 4586
rect 10317 4528 10322 4584
rect 10378 4528 12450 4584
rect 10317 4526 12450 4528
rect 10317 4523 10383 4526
rect 12390 4450 12450 4526
rect 12617 4584 16455 4586
rect 12617 4528 12622 4584
rect 12678 4528 16394 4584
rect 16450 4528 16455 4584
rect 12617 4526 16455 4528
rect 12617 4523 12683 4526
rect 16389 4523 16455 4526
rect 18140 4584 18939 4586
rect 18140 4528 18878 4584
rect 18934 4528 18939 4584
rect 18140 4526 18939 4528
rect 18140 4450 18200 4526
rect 18873 4523 18939 4526
rect 12390 4390 18200 4450
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 9673 4316 9739 4317
rect 9622 4252 9628 4316
rect 9692 4314 9739 4316
rect 9692 4312 9784 4314
rect 9734 4256 9784 4312
rect 9692 4254 9784 4256
rect 9692 4252 9739 4254
rect 12566 4252 12572 4316
rect 12636 4314 12642 4316
rect 12709 4314 12775 4317
rect 12636 4312 12775 4314
rect 12636 4256 12714 4312
rect 12770 4256 12775 4312
rect 12636 4254 12775 4256
rect 12636 4252 12642 4254
rect 9673 4251 9739 4252
rect 12709 4251 12775 4254
rect 0 4178 480 4208
rect 3969 4178 4035 4181
rect 0 4176 4035 4178
rect 0 4120 3974 4176
rect 4030 4120 4035 4176
rect 0 4118 4035 4120
rect 0 4088 480 4118
rect 3969 4115 4035 4118
rect 10041 4178 10107 4181
rect 12801 4178 12867 4181
rect 13537 4178 13603 4181
rect 10041 4176 13603 4178
rect 10041 4120 10046 4176
rect 10102 4120 12806 4176
rect 12862 4120 13542 4176
rect 13598 4120 13603 4176
rect 10041 4118 13603 4120
rect 10041 4115 10107 4118
rect 12801 4115 12867 4118
rect 13537 4115 13603 4118
rect 15285 4178 15351 4181
rect 22520 4178 23000 4208
rect 15285 4176 23000 4178
rect 15285 4120 15290 4176
rect 15346 4120 23000 4176
rect 15285 4118 23000 4120
rect 15285 4115 15351 4118
rect 22520 4088 23000 4118
rect 4153 4042 4219 4045
rect 19885 4042 19951 4045
rect 4153 4040 19951 4042
rect 4153 3984 4158 4040
rect 4214 3984 19890 4040
rect 19946 3984 19951 4040
rect 4153 3982 19951 3984
rect 4153 3979 4219 3982
rect 19885 3979 19951 3982
rect 10685 3906 10751 3909
rect 16113 3906 16179 3909
rect 16481 3906 16547 3909
rect 10685 3904 14704 3906
rect 10685 3848 10690 3904
rect 10746 3848 14704 3904
rect 10685 3846 14704 3848
rect 10685 3843 10751 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 10041 3770 10107 3773
rect 10174 3770 10180 3772
rect 10041 3768 10180 3770
rect 10041 3712 10046 3768
rect 10102 3712 10180 3768
rect 10041 3710 10180 3712
rect 10041 3707 10107 3710
rect 10174 3708 10180 3710
rect 10244 3708 10250 3772
rect 0 3634 480 3664
rect 3969 3634 4035 3637
rect 0 3632 4035 3634
rect 0 3576 3974 3632
rect 4030 3576 4035 3632
rect 0 3574 4035 3576
rect 0 3544 480 3574
rect 3969 3571 4035 3574
rect 8201 3634 8267 3637
rect 14644 3634 14704 3846
rect 16113 3904 16547 3906
rect 16113 3848 16118 3904
rect 16174 3848 16486 3904
rect 16542 3848 16547 3904
rect 16113 3846 16547 3848
rect 16113 3843 16179 3846
rect 16481 3843 16547 3846
rect 18137 3906 18203 3909
rect 18822 3906 18828 3908
rect 18137 3904 18828 3906
rect 18137 3848 18142 3904
rect 18198 3848 18828 3904
rect 18137 3846 18828 3848
rect 18137 3843 18203 3846
rect 18822 3844 18828 3846
rect 18892 3844 18898 3908
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 3775 15125 3776
rect 15193 3770 15259 3773
rect 18321 3770 18387 3773
rect 15193 3768 18387 3770
rect 15193 3712 15198 3768
rect 15254 3712 18326 3768
rect 18382 3712 18387 3768
rect 15193 3710 18387 3712
rect 15193 3707 15259 3710
rect 18321 3707 18387 3710
rect 16665 3634 16731 3637
rect 8201 3632 12634 3634
rect 8201 3576 8206 3632
rect 8262 3576 12634 3632
rect 8201 3574 12634 3576
rect 14644 3632 16731 3634
rect 14644 3576 16670 3632
rect 16726 3576 16731 3632
rect 14644 3574 16731 3576
rect 8201 3571 8267 3574
rect 4245 3498 4311 3501
rect 12574 3498 12634 3574
rect 16665 3571 16731 3574
rect 17769 3634 17835 3637
rect 22520 3634 23000 3664
rect 17769 3632 23000 3634
rect 17769 3576 17774 3632
rect 17830 3576 23000 3632
rect 17769 3574 23000 3576
rect 17769 3571 17835 3574
rect 22520 3544 23000 3574
rect 20989 3498 21055 3501
rect 4245 3496 12450 3498
rect 4245 3440 4250 3496
rect 4306 3440 12450 3496
rect 4245 3438 12450 3440
rect 12574 3496 21055 3498
rect 12574 3440 20994 3496
rect 21050 3440 21055 3496
rect 12574 3438 21055 3440
rect 4245 3435 4311 3438
rect 12390 3362 12450 3438
rect 20989 3435 21055 3438
rect 12390 3302 12818 3362
rect 4409 3296 4729 3297
rect 0 3226 480 3256
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 3693 3226 3759 3229
rect 0 3224 3759 3226
rect 0 3168 3698 3224
rect 3754 3168 3759 3224
rect 0 3166 3759 3168
rect 0 3136 480 3166
rect 3693 3163 3759 3166
rect 9581 3090 9647 3093
rect 12617 3090 12683 3093
rect 9581 3088 12683 3090
rect 9581 3032 9586 3088
rect 9642 3032 12622 3088
rect 12678 3032 12683 3088
rect 9581 3030 12683 3032
rect 12758 3090 12818 3302
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 13813 3226 13879 3229
rect 15745 3226 15811 3229
rect 16757 3228 16823 3229
rect 16757 3226 16804 3228
rect 13813 3224 15811 3226
rect 13813 3168 13818 3224
rect 13874 3168 15750 3224
rect 15806 3168 15811 3224
rect 13813 3166 15811 3168
rect 16712 3224 16804 3226
rect 16712 3168 16762 3224
rect 16712 3166 16804 3168
rect 13813 3163 13879 3166
rect 15745 3163 15811 3166
rect 16757 3164 16804 3166
rect 16868 3164 16874 3228
rect 20529 3226 20595 3229
rect 22520 3226 23000 3256
rect 20529 3224 23000 3226
rect 20529 3168 20534 3224
rect 20590 3168 23000 3224
rect 20529 3166 23000 3168
rect 16757 3163 16823 3164
rect 20529 3163 20595 3166
rect 22520 3136 23000 3166
rect 21173 3090 21239 3093
rect 12758 3088 21239 3090
rect 12758 3032 21178 3088
rect 21234 3032 21239 3088
rect 12758 3030 21239 3032
rect 9581 3027 9647 3030
rect 12617 3027 12683 3030
rect 21173 3027 21239 3030
rect 3049 2954 3115 2957
rect 21265 2954 21331 2957
rect 3049 2952 21331 2954
rect 3049 2896 3054 2952
rect 3110 2896 21270 2952
rect 21326 2896 21331 2952
rect 3049 2894 21331 2896
rect 3049 2891 3115 2894
rect 21265 2891 21331 2894
rect 1761 2818 1827 2821
rect 7557 2818 7623 2821
rect 1761 2816 7623 2818
rect 1761 2760 1766 2816
rect 1822 2760 7562 2816
rect 7618 2760 7623 2816
rect 1761 2758 7623 2760
rect 1761 2755 1827 2758
rect 7557 2755 7623 2758
rect 7874 2752 8194 2753
rect 0 2682 480 2712
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 3417 2682 3483 2685
rect 0 2680 3483 2682
rect 0 2624 3422 2680
rect 3478 2624 3483 2680
rect 0 2622 3483 2624
rect 0 2592 480 2622
rect 3417 2619 3483 2622
rect 15469 2682 15535 2685
rect 22520 2682 23000 2712
rect 15469 2680 23000 2682
rect 15469 2624 15474 2680
rect 15530 2624 23000 2680
rect 15469 2622 23000 2624
rect 15469 2619 15535 2622
rect 22520 2592 23000 2622
rect 1894 2484 1900 2548
rect 1964 2546 1970 2548
rect 19425 2546 19491 2549
rect 1964 2544 19491 2546
rect 1964 2488 19430 2544
rect 19486 2488 19491 2544
rect 1964 2486 19491 2488
rect 1964 2484 1970 2486
rect 19425 2483 19491 2486
rect 4409 2208 4729 2209
rect 0 2138 480 2168
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 2773 2138 2839 2141
rect 0 2136 2839 2138
rect 0 2080 2778 2136
rect 2834 2080 2839 2136
rect 0 2078 2839 2080
rect 0 2048 480 2078
rect 2773 2075 2839 2078
rect 18689 2138 18755 2141
rect 22520 2138 23000 2168
rect 18689 2136 23000 2138
rect 18689 2080 18694 2136
rect 18750 2080 23000 2136
rect 18689 2078 23000 2080
rect 18689 2075 18755 2078
rect 22520 2048 23000 2078
rect 0 1730 480 1760
rect 4061 1730 4127 1733
rect 0 1728 4127 1730
rect 0 1672 4066 1728
rect 4122 1672 4127 1728
rect 0 1670 4127 1672
rect 0 1640 480 1670
rect 4061 1667 4127 1670
rect 18505 1730 18571 1733
rect 22520 1730 23000 1760
rect 18505 1728 23000 1730
rect 18505 1672 18510 1728
rect 18566 1672 23000 1728
rect 18505 1670 23000 1672
rect 18505 1667 18571 1670
rect 22520 1640 23000 1670
rect 0 1186 480 1216
rect 2589 1186 2655 1189
rect 0 1184 2655 1186
rect 0 1128 2594 1184
rect 2650 1128 2655 1184
rect 0 1126 2655 1128
rect 0 1096 480 1126
rect 2589 1123 2655 1126
rect 12065 1186 12131 1189
rect 22520 1186 23000 1216
rect 12065 1184 23000 1186
rect 12065 1128 12070 1184
rect 12126 1128 23000 1184
rect 12065 1126 23000 1128
rect 12065 1123 12131 1126
rect 22520 1096 23000 1126
rect 0 642 480 672
rect 3601 642 3667 645
rect 0 640 3667 642
rect 0 584 3606 640
rect 3662 584 3667 640
rect 0 582 3667 584
rect 0 552 480 582
rect 3601 579 3667 582
rect 18137 642 18203 645
rect 22520 642 23000 672
rect 18137 640 23000 642
rect 18137 584 18142 640
rect 18198 584 23000 640
rect 18137 582 23000 584
rect 18137 579 18203 582
rect 22520 552 23000 582
rect 0 234 480 264
rect 3233 234 3299 237
rect 0 232 3299 234
rect 0 176 3238 232
rect 3294 176 3299 232
rect 0 174 3299 176
rect 0 144 480 174
rect 3233 171 3299 174
rect 11881 234 11947 237
rect 22520 234 23000 264
rect 11881 232 23000 234
rect 11881 176 11886 232
rect 11942 176 23000 232
rect 11881 174 23000 176
rect 11881 171 11947 174
rect 22520 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 8340 20360 8404 20364
rect 8340 20304 8354 20360
rect 8354 20304 8404 20360
rect 8340 20300 8404 20304
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 8340 19136 8404 19140
rect 8340 19080 8354 19136
rect 8354 19080 8404 19136
rect 8340 19076 8404 19080
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 5580 18804 5644 18868
rect 14596 18668 14660 18732
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 17724 18124 17788 18188
rect 16620 17988 16684 18052
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 13308 17368 13372 17372
rect 13308 17312 13358 17368
rect 13358 17312 13372 17368
rect 13308 17308 13372 17312
rect 8524 17172 8588 17236
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 5212 16628 5276 16692
rect 17724 16628 17788 16692
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7236 15132 7300 15196
rect 3372 14996 3436 15060
rect 16988 15056 17052 15060
rect 16988 15000 17002 15056
rect 17002 15000 17052 15056
rect 16988 14996 17052 15000
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11836 14860 11900 14924
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 13124 14452 13188 14516
rect 19748 14452 19812 14516
rect 11100 14316 11164 14380
rect 15700 14316 15764 14380
rect 17908 14316 17972 14380
rect 19012 14376 19076 14380
rect 19012 14320 19062 14376
rect 19062 14320 19076 14376
rect 19012 14316 19076 14320
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 10180 13636 10244 13700
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 5212 12548 5276 12612
rect 12940 12548 13004 12612
rect 18092 12608 18156 12612
rect 18092 12552 18106 12608
rect 18106 12552 18156 12608
rect 18092 12548 18156 12552
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 1900 12472 1964 12476
rect 1900 12416 1914 12472
rect 1914 12416 1964 12472
rect 1900 12412 1964 12416
rect 2452 12412 2516 12476
rect 5212 12472 5276 12476
rect 5212 12416 5262 12472
rect 5262 12416 5276 12472
rect 5212 12412 5276 12416
rect 5396 12472 5460 12476
rect 5396 12416 5446 12472
rect 5446 12416 5460 12472
rect 5396 12412 5460 12416
rect 13308 12472 13372 12476
rect 13308 12416 13358 12472
rect 13358 12416 13372 12472
rect 13308 12412 13372 12416
rect 16068 12412 16132 12476
rect 11836 12276 11900 12340
rect 12940 12336 13004 12340
rect 12940 12280 12954 12336
rect 12954 12280 13004 12336
rect 12940 12276 13004 12280
rect 15332 12276 15396 12340
rect 18092 12336 18156 12340
rect 18092 12280 18142 12336
rect 18142 12280 18156 12336
rect 18092 12276 18156 12280
rect 18828 12336 18892 12340
rect 18828 12280 18842 12336
rect 18842 12280 18892 12336
rect 18828 12276 18892 12280
rect 8524 12140 8588 12204
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 2452 11732 2516 11796
rect 13676 12140 13740 12204
rect 16436 12140 16500 12204
rect 16068 12064 16132 12068
rect 16068 12008 16082 12064
rect 16082 12008 16132 12064
rect 16068 12004 16132 12008
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 15516 11868 15580 11932
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 16068 11324 16132 11388
rect 5396 11052 5460 11116
rect 14596 11052 14660 11116
rect 16988 11384 17052 11388
rect 16988 11328 17038 11384
rect 17038 11328 17052 11384
rect 16988 11324 17052 11328
rect 19012 11052 19076 11116
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 3924 10644 3988 10708
rect 5580 10644 5644 10708
rect 4108 10508 4172 10572
rect 15700 10372 15764 10436
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 13676 10296 13740 10300
rect 13676 10240 13726 10296
rect 13726 10240 13740 10296
rect 13676 10236 13740 10240
rect 7236 9964 7300 10028
rect 7604 9964 7668 10028
rect 13124 9964 13188 10028
rect 15516 9964 15580 10028
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 10548 9556 10612 9620
rect 16988 9556 17052 9620
rect 14044 9420 14108 9484
rect 15516 9420 15580 9484
rect 13308 9284 13372 9348
rect 17908 9284 17972 9348
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 11100 9148 11164 9212
rect 12572 9012 12636 9076
rect 13860 9072 13924 9076
rect 16804 9148 16868 9212
rect 13860 9016 13874 9072
rect 13874 9016 13924 9072
rect 13860 9012 13924 9016
rect 4108 8876 4172 8940
rect 7236 8800 7300 8804
rect 7236 8744 7250 8800
rect 7250 8744 7300 8800
rect 7236 8740 7300 8744
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7604 8604 7668 8668
rect 15700 8392 15764 8396
rect 15700 8336 15714 8392
rect 15714 8336 15764 8392
rect 15700 8332 15764 8336
rect 16068 8392 16132 8396
rect 16068 8336 16118 8392
rect 16118 8336 16132 8392
rect 16068 8332 16132 8336
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 15332 8060 15396 8124
rect 18828 7924 18892 7988
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 3924 7380 3988 7444
rect 5212 7380 5276 7444
rect 16436 7440 16500 7444
rect 16436 7384 16450 7440
rect 16450 7384 16500 7440
rect 16436 7380 16500 7384
rect 9628 7304 9692 7308
rect 9628 7248 9678 7304
rect 9678 7248 9692 7304
rect 9628 7244 9692 7248
rect 9812 7168 9876 7172
rect 9812 7112 9826 7168
rect 9826 7112 9876 7168
rect 9812 7108 9876 7112
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 18828 7304 18892 7308
rect 18828 7248 18878 7304
rect 18878 7248 18892 7304
rect 18828 7244 18892 7248
rect 19748 7244 19812 7308
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 15332 6292 15396 6356
rect 14044 6020 14108 6084
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 9812 5884 9876 5948
rect 13308 5884 13372 5948
rect 13860 5944 13924 5948
rect 13860 5888 13874 5944
rect 13874 5888 13924 5944
rect 13860 5884 13924 5888
rect 14596 5944 14660 5948
rect 14596 5888 14646 5944
rect 14646 5888 14660 5944
rect 14596 5884 14660 5888
rect 3372 5612 3436 5676
rect 15516 5748 15580 5812
rect 16620 5612 16684 5676
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 16988 5340 17052 5404
rect 5212 5204 5276 5268
rect 5396 5264 5460 5268
rect 5396 5208 5446 5264
rect 5446 5208 5460 5264
rect 5396 5204 5460 5208
rect 17908 5204 17972 5268
rect 4108 5128 4172 5132
rect 4108 5072 4158 5128
rect 4158 5072 4172 5128
rect 4108 5068 4172 5072
rect 10548 4932 10612 4996
rect 17908 4932 17972 4996
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 9628 4312 9692 4316
rect 9628 4256 9678 4312
rect 9678 4256 9692 4312
rect 9628 4252 9692 4256
rect 12572 4252 12636 4316
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 10180 3708 10244 3772
rect 18828 3844 18892 3908
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 16804 3224 16868 3228
rect 16804 3168 16818 3224
rect 16818 3168 16868 3224
rect 16804 3164 16868 3168
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 1900 2484 1964 2548
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 7874 20160 8195 20720
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 8339 20364 8405 20365
rect 8339 20300 8340 20364
rect 8404 20300 8405 20364
rect 8339 20299 8405 20300
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 8342 19141 8402 20299
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 8339 19140 8405 19141
rect 8339 19076 8340 19140
rect 8404 19076 8405 19140
rect 8339 19075 8405 19076
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 5579 18868 5645 18869
rect 5579 18804 5580 18868
rect 5644 18804 5645 18868
rect 5579 18803 5645 18804
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 5211 16692 5277 16693
rect 5211 16628 5212 16692
rect 5276 16628 5277 16692
rect 5211 16627 5277 16628
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 3371 15060 3437 15061
rect 3371 14996 3372 15060
rect 3436 14996 3437 15060
rect 3371 14995 3437 14996
rect 1899 12476 1965 12477
rect 1899 12412 1900 12476
rect 1964 12412 1965 12476
rect 1899 12411 1965 12412
rect 2451 12476 2517 12477
rect 2451 12412 2452 12476
rect 2516 12412 2517 12476
rect 2451 12411 2517 12412
rect 1902 2549 1962 12411
rect 2454 11797 2514 12411
rect 2451 11796 2517 11797
rect 2451 11732 2452 11796
rect 2516 11732 2517 11796
rect 2451 11731 2517 11732
rect 3374 5677 3434 14995
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 5214 12613 5274 16627
rect 5211 12612 5277 12613
rect 5211 12548 5212 12612
rect 5276 12548 5277 12612
rect 5211 12547 5277 12548
rect 5211 12476 5277 12477
rect 5211 12412 5212 12476
rect 5276 12412 5277 12476
rect 5211 12411 5277 12412
rect 5395 12476 5461 12477
rect 5395 12412 5396 12476
rect 5460 12412 5461 12476
rect 5395 12411 5461 12412
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 3923 10708 3989 10709
rect 3923 10644 3924 10708
rect 3988 10644 3989 10708
rect 3923 10643 3989 10644
rect 3926 7445 3986 10643
rect 4107 10572 4173 10573
rect 4107 10508 4108 10572
rect 4172 10508 4173 10572
rect 4107 10507 4173 10508
rect 4110 8941 4170 10507
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4107 8940 4173 8941
rect 4107 8876 4108 8940
rect 4172 8876 4173 8940
rect 4107 8875 4173 8876
rect 3923 7444 3989 7445
rect 3923 7380 3924 7444
rect 3988 7380 3989 7444
rect 3923 7379 3989 7380
rect 3371 5676 3437 5677
rect 3371 5612 3372 5676
rect 3436 5612 3437 5676
rect 3371 5611 3437 5612
rect 4110 5133 4170 8875
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 5214 7445 5274 12411
rect 5398 11117 5458 12411
rect 5395 11116 5461 11117
rect 5395 11052 5396 11116
rect 5460 11052 5461 11116
rect 5395 11051 5461 11052
rect 5211 7444 5277 7445
rect 5211 7380 5212 7444
rect 5276 7380 5277 7444
rect 5211 7379 5277 7380
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4107 5132 4173 5133
rect 4107 5068 4108 5132
rect 4172 5068 4173 5132
rect 4107 5067 4173 5068
rect 4409 4384 4729 5408
rect 5214 5269 5274 7379
rect 5398 5269 5458 11051
rect 5582 10709 5642 18803
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 11340 18528 11660 19552
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14595 18732 14661 18733
rect 14595 18668 14596 18732
rect 14660 18668 14661 18732
rect 14595 18667 14661 18668
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 8523 17236 8589 17237
rect 8523 17172 8524 17236
rect 8588 17172 8589 17236
rect 8523 17171 8589 17172
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7235 15196 7301 15197
rect 7235 15132 7236 15196
rect 7300 15132 7301 15196
rect 7235 15131 7301 15132
rect 5579 10708 5645 10709
rect 5579 10644 5580 10708
rect 5644 10644 5645 10708
rect 5579 10643 5645 10644
rect 7238 10029 7298 15131
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 8526 12205 8586 17171
rect 11340 16352 11660 17376
rect 13307 17372 13373 17373
rect 13307 17308 13308 17372
rect 13372 17308 13373 17372
rect 13307 17307 13373 17308
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11099 14380 11165 14381
rect 11099 14316 11100 14380
rect 11164 14316 11165 14380
rect 11099 14315 11165 14316
rect 10179 13700 10245 13701
rect 10179 13636 10180 13700
rect 10244 13636 10245 13700
rect 10179 13635 10245 13636
rect 8523 12204 8589 12205
rect 8523 12140 8524 12204
rect 8588 12140 8589 12204
rect 8523 12139 8589 12140
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7235 10028 7301 10029
rect 7235 9964 7236 10028
rect 7300 9964 7301 10028
rect 7235 9963 7301 9964
rect 7603 10028 7669 10029
rect 7603 9964 7604 10028
rect 7668 9964 7669 10028
rect 7603 9963 7669 9964
rect 7238 8805 7298 9963
rect 7235 8804 7301 8805
rect 7235 8740 7236 8804
rect 7300 8740 7301 8804
rect 7235 8739 7301 8740
rect 7606 8669 7666 9963
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7603 8668 7669 8669
rect 7603 8604 7604 8668
rect 7668 8604 7669 8668
rect 7603 8603 7669 8604
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 9627 7308 9693 7309
rect 9627 7244 9628 7308
rect 9692 7244 9693 7308
rect 9627 7243 9693 7244
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 5211 5268 5277 5269
rect 5211 5204 5212 5268
rect 5276 5204 5277 5268
rect 5211 5203 5277 5204
rect 5395 5268 5461 5269
rect 5395 5204 5396 5268
rect 5460 5204 5461 5268
rect 5395 5203 5461 5204
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 1899 2548 1965 2549
rect 1899 2484 1900 2548
rect 1964 2484 1965 2548
rect 1899 2483 1965 2484
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 9630 4317 9690 7243
rect 9811 7172 9877 7173
rect 9811 7108 9812 7172
rect 9876 7108 9877 7172
rect 9811 7107 9877 7108
rect 9814 5949 9874 7107
rect 9811 5948 9877 5949
rect 9811 5884 9812 5948
rect 9876 5884 9877 5948
rect 9811 5883 9877 5884
rect 9627 4316 9693 4317
rect 9627 4252 9628 4316
rect 9692 4252 9693 4316
rect 9627 4251 9693 4252
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 10182 3773 10242 13635
rect 10547 9620 10613 9621
rect 10547 9556 10548 9620
rect 10612 9556 10613 9620
rect 10547 9555 10613 9556
rect 10550 4997 10610 9555
rect 11102 9213 11162 14315
rect 11340 14176 11660 15200
rect 11835 14924 11901 14925
rect 11835 14860 11836 14924
rect 11900 14860 11901 14924
rect 11835 14859 11901 14860
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11838 12341 11898 14859
rect 13123 14516 13189 14517
rect 13123 14452 13124 14516
rect 13188 14452 13189 14516
rect 13123 14451 13189 14452
rect 12939 12612 13005 12613
rect 12939 12548 12940 12612
rect 13004 12548 13005 12612
rect 12939 12547 13005 12548
rect 12942 12341 13002 12547
rect 11835 12340 11901 12341
rect 11835 12276 11836 12340
rect 11900 12276 11901 12340
rect 11835 12275 11901 12276
rect 12939 12340 13005 12341
rect 12939 12276 12940 12340
rect 13004 12276 13005 12340
rect 12939 12275 13005 12276
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 13126 10029 13186 14451
rect 13310 12477 13370 17307
rect 13307 12476 13373 12477
rect 13307 12412 13308 12476
rect 13372 12412 13373 12476
rect 13307 12411 13373 12412
rect 13675 12204 13741 12205
rect 13675 12140 13676 12204
rect 13740 12140 13741 12204
rect 13675 12139 13741 12140
rect 13678 10301 13738 12139
rect 14598 11117 14658 18667
rect 14805 17984 15125 19008
rect 18270 20704 18590 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 19616 18590 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 18528 18590 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 17723 18188 17789 18189
rect 17723 18124 17724 18188
rect 17788 18124 17789 18188
rect 17723 18123 17789 18124
rect 16619 18052 16685 18053
rect 16619 17988 16620 18052
rect 16684 17988 16685 18052
rect 16619 17987 16685 17988
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 15699 14380 15765 14381
rect 15699 14316 15700 14380
rect 15764 14316 15765 14380
rect 15699 14315 15765 14316
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 15331 12340 15397 12341
rect 15331 12276 15332 12340
rect 15396 12276 15397 12340
rect 15331 12275 15397 12276
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14595 11116 14661 11117
rect 14595 11052 14596 11116
rect 14660 11052 14661 11116
rect 14595 11051 14661 11052
rect 13675 10300 13741 10301
rect 13675 10236 13676 10300
rect 13740 10236 13741 10300
rect 13675 10235 13741 10236
rect 13123 10028 13189 10029
rect 13123 9964 13124 10028
rect 13188 9964 13189 10028
rect 13123 9963 13189 9964
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11099 9212 11165 9213
rect 11099 9148 11100 9212
rect 11164 9148 11165 9212
rect 11099 9147 11165 9148
rect 11340 8736 11660 9760
rect 14043 9484 14109 9485
rect 14043 9420 14044 9484
rect 14108 9420 14109 9484
rect 14043 9419 14109 9420
rect 13307 9348 13373 9349
rect 13307 9284 13308 9348
rect 13372 9284 13373 9348
rect 13307 9283 13373 9284
rect 12571 9076 12637 9077
rect 12571 9012 12572 9076
rect 12636 9012 12637 9076
rect 12571 9011 12637 9012
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 10547 4996 10613 4997
rect 10547 4932 10548 4996
rect 10612 4932 10613 4996
rect 10547 4931 10613 4932
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 10179 3772 10245 3773
rect 10179 3708 10180 3772
rect 10244 3708 10245 3772
rect 10179 3707 10245 3708
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 3296 11660 4320
rect 12574 4317 12634 9011
rect 13310 5949 13370 9283
rect 13859 9076 13925 9077
rect 13859 9012 13860 9076
rect 13924 9012 13925 9076
rect 13859 9011 13925 9012
rect 13862 5949 13922 9011
rect 14046 6085 14106 9419
rect 14043 6084 14109 6085
rect 14043 6020 14044 6084
rect 14108 6020 14109 6084
rect 14043 6019 14109 6020
rect 14598 5949 14658 11051
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 15334 8125 15394 12275
rect 15515 11932 15581 11933
rect 15515 11868 15516 11932
rect 15580 11868 15581 11932
rect 15515 11867 15581 11868
rect 15518 10029 15578 11867
rect 15702 10437 15762 14315
rect 16067 12476 16133 12477
rect 16067 12412 16068 12476
rect 16132 12412 16133 12476
rect 16067 12411 16133 12412
rect 16070 12069 16130 12411
rect 16435 12204 16501 12205
rect 16435 12140 16436 12204
rect 16500 12140 16501 12204
rect 16435 12139 16501 12140
rect 16067 12068 16133 12069
rect 16067 12004 16068 12068
rect 16132 12004 16133 12068
rect 16067 12003 16133 12004
rect 16067 11388 16133 11389
rect 16067 11324 16068 11388
rect 16132 11324 16133 11388
rect 16067 11323 16133 11324
rect 15699 10436 15765 10437
rect 15699 10372 15700 10436
rect 15764 10372 15765 10436
rect 15699 10371 15765 10372
rect 15515 10028 15581 10029
rect 15515 9964 15516 10028
rect 15580 9964 15581 10028
rect 15515 9963 15581 9964
rect 15515 9484 15581 9485
rect 15515 9420 15516 9484
rect 15580 9420 15581 9484
rect 15515 9419 15581 9420
rect 15331 8124 15397 8125
rect 15331 8060 15332 8124
rect 15396 8060 15397 8124
rect 15331 8059 15397 8060
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 15334 6357 15394 8059
rect 15331 6356 15397 6357
rect 15331 6292 15332 6356
rect 15396 6292 15397 6356
rect 15331 6291 15397 6292
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 13307 5948 13373 5949
rect 13307 5884 13308 5948
rect 13372 5884 13373 5948
rect 13307 5883 13373 5884
rect 13859 5948 13925 5949
rect 13859 5884 13860 5948
rect 13924 5884 13925 5948
rect 13859 5883 13925 5884
rect 14595 5948 14661 5949
rect 14595 5884 14596 5948
rect 14660 5884 14661 5948
rect 14595 5883 14661 5884
rect 14805 4928 15125 5952
rect 15518 5813 15578 9419
rect 15702 8397 15762 10371
rect 16070 8397 16130 11323
rect 15699 8396 15765 8397
rect 15699 8332 15700 8396
rect 15764 8332 15765 8396
rect 15699 8331 15765 8332
rect 16067 8396 16133 8397
rect 16067 8332 16068 8396
rect 16132 8332 16133 8396
rect 16067 8331 16133 8332
rect 16438 7445 16498 12139
rect 16435 7444 16501 7445
rect 16435 7380 16436 7444
rect 16500 7380 16501 7444
rect 16435 7379 16501 7380
rect 15515 5812 15581 5813
rect 15515 5748 15516 5812
rect 15580 5748 15581 5812
rect 15515 5747 15581 5748
rect 16622 5677 16682 17987
rect 17726 16693 17786 18123
rect 18270 17440 18590 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 17723 16692 17789 16693
rect 17723 16628 17724 16692
rect 17788 16628 17789 16692
rect 17723 16627 17789 16628
rect 18270 16352 18590 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 15264 18590 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 16987 15060 17053 15061
rect 16987 14996 16988 15060
rect 17052 14996 17053 15060
rect 16987 14995 17053 14996
rect 16990 11389 17050 14995
rect 17907 14380 17973 14381
rect 17907 14316 17908 14380
rect 17972 14316 17973 14380
rect 17907 14315 17973 14316
rect 16987 11388 17053 11389
rect 16987 11324 16988 11388
rect 17052 11324 17053 11388
rect 16987 11323 17053 11324
rect 16987 9620 17053 9621
rect 16987 9556 16988 9620
rect 17052 9556 17053 9620
rect 16987 9555 17053 9556
rect 16803 9212 16869 9213
rect 16803 9148 16804 9212
rect 16868 9148 16869 9212
rect 16803 9147 16869 9148
rect 16619 5676 16685 5677
rect 16619 5612 16620 5676
rect 16684 5612 16685 5676
rect 16619 5611 16685 5612
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 12571 4316 12637 4317
rect 12571 4252 12572 4316
rect 12636 4252 12637 4316
rect 12571 4251 12637 4252
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 16806 3229 16866 9147
rect 16990 5405 17050 9555
rect 17910 9349 17970 14315
rect 18270 14176 18590 15200
rect 19747 14516 19813 14517
rect 19747 14452 19748 14516
rect 19812 14452 19813 14516
rect 19747 14451 19813 14452
rect 19011 14380 19077 14381
rect 19011 14316 19012 14380
rect 19076 14316 19077 14380
rect 19011 14315 19077 14316
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 13088 18590 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18091 12612 18157 12613
rect 18091 12548 18092 12612
rect 18156 12548 18157 12612
rect 18091 12547 18157 12548
rect 18094 12341 18154 12547
rect 18091 12340 18157 12341
rect 18091 12276 18092 12340
rect 18156 12276 18157 12340
rect 18091 12275 18157 12276
rect 18270 12000 18590 13024
rect 18827 12340 18893 12341
rect 18827 12276 18828 12340
rect 18892 12276 18893 12340
rect 18827 12275 18893 12276
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 10912 18590 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 9824 18590 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 17907 9348 17973 9349
rect 17907 9284 17908 9348
rect 17972 9284 17973 9348
rect 17907 9283 17973 9284
rect 18270 8736 18590 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 7648 18590 8672
rect 18830 7989 18890 12275
rect 19014 11117 19074 14315
rect 19011 11116 19077 11117
rect 19011 11052 19012 11116
rect 19076 11052 19077 11116
rect 19011 11051 19077 11052
rect 18827 7988 18893 7989
rect 18827 7924 18828 7988
rect 18892 7924 18893 7988
rect 18827 7923 18893 7924
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 6560 18590 7584
rect 19750 7309 19810 14451
rect 18827 7308 18893 7309
rect 18827 7244 18828 7308
rect 18892 7244 18893 7308
rect 18827 7243 18893 7244
rect 19747 7308 19813 7309
rect 19747 7244 19748 7308
rect 19812 7244 19813 7308
rect 19747 7243 19813 7244
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 5472 18590 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 16987 5404 17053 5405
rect 16987 5340 16988 5404
rect 17052 5340 17053 5404
rect 16987 5339 17053 5340
rect 17907 5268 17973 5269
rect 17907 5204 17908 5268
rect 17972 5204 17973 5268
rect 17907 5203 17973 5204
rect 17910 4997 17970 5203
rect 17907 4996 17973 4997
rect 17907 4932 17908 4996
rect 17972 4932 17973 4996
rect 17907 4931 17973 4932
rect 18270 4384 18590 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 3296 18590 4320
rect 18830 3909 18890 7243
rect 18827 3908 18893 3909
rect 18827 3844 18828 3908
rect 18892 3844 18893 3908
rect 18827 3843 18893 3844
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 16803 3228 16869 3229
rect 16803 3164 16804 3228
rect 16868 3164 16869 3228
rect 16803 3163 16869 3164
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 2208 18590 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2128 18590 2144
use sky130_fd_sc_hd__decap_4  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _103_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1840 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604681595
transform 1 0 1748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2116 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 2852 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_12 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2208 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3312 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30
timestamp 1604681595
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_23
timestamp 1604681595
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_35
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _057_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_47
timestamp 1604681595
transform 1 0 5428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 7636 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74
timestamp 1604681595
transform 1 0 7912 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1604681595
transform 1 0 8648 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1604681595
transform 1 0 10396 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100
timestamp 1604681595
transform 1 0 10304 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp 1604681595
transform 1 0 10672 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_94
timestamp 1604681595
transform 1 0 9752 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_102
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 12696 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 14076 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130
timestamp 1604681595
transform 1 0 13064 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_133
timestamp 1604681595
transform 1 0 13340 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp 1604681595
transform 1 0 15732 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_150
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_162
timestamp 1604681595
transform 1 0 16008 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_176
timestamp 1604681595
transform 1 0 17296 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_175
timestamp 1604681595
transform 1 0 17204 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_191
timestamp 1604681595
transform 1 0 18676 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_203
timestamp 1604681595
transform 1 0 19780 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_193
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1604681595
transform 1 0 19964 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1604681595
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1604681595
transform 1 0 21068 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604681595
transform 1 0 1840 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_12
timestamp 1604681595
transform 1 0 2208 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_36
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 6532 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_48
timestamp 1604681595
transform 1 0 5520 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_62
timestamp 1604681595
transform 1 0 6808 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 7544 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_73
timestamp 1604681595
transform 1 0 7820 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 9844 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_99
timestamp 1604681595
transform 1 0 10212 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 10948 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12052 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_111
timestamp 1604681595
transform 1 0 11316 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_128
timestamp 1604681595
transform 1 0 12880 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16008 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17572 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_171
timestamp 1604681595
transform 1 0 16836 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19136 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1604681595
transform 1 0 18400 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_205
timestamp 1604681595
transform 1 0 19964 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1604681595
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_11
timestamp 1604681595
transform 1 0 2116 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 3956 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_23
timestamp 1604681595
transform 1 0 3220 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_35
timestamp 1604681595
transform 1 0 4324 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 5060 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_46
timestamp 1604681595
transform 1 0 5336 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1604681595
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 6900 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_66
timestamp 1604681595
transform 1 0 7176 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_78
timestamp 1604681595
transform 1 0 8280 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_90
timestamp 1604681595
transform 1 0 9384 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_102
timestamp 1604681595
transform 1 0 10488 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12512 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 14076 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_133
timestamp 1604681595
transform 1 0 13340 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16100 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_150
timestamp 1604681595
transform 1 0 14904 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_162
timestamp 1604681595
transform 1 0 16008 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_172
timestamp 1604681595
transform 1 0 16928 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_178
timestamp 1604681595
transform 1 0 17480 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_195
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_210
timestamp 1604681595
transform 1 0 20424 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_222
timestamp 1604681595
transform 1 0 21528 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 2852 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_11
timestamp 1604681595
transform 1 0 2116 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_36
timestamp 1604681595
transform 1 0 4416 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 6348 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_48
timestamp 1604681595
transform 1 0 5520 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_60
timestamp 1604681595
transform 1 0 6624 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_72
timestamp 1604681595
transform 1 0 7728 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 9936 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_84
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_100
timestamp 1604681595
transform 1 0 10304 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 12604 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11040 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_128
timestamp 1604681595
transform 1 0 12880 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_158
timestamp 1604681595
transform 1 0 15640 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18124 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16468 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_176
timestamp 1604681595
transform 1 0 17296 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_184
timestamp 1604681595
transform 1 0 18032 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_194
timestamp 1604681595
transform 1 0 18952 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_11
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604681595
transform 1 0 3956 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_23
timestamp 1604681595
transform 1 0 3220 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_35
timestamp 1604681595
transform 1 0 4324 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604681595
transform 1 0 5060 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_47
timestamp 1604681595
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 8004 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 6900 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_67
timestamp 1604681595
transform 1 0 7268 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_79
timestamp 1604681595
transform 1 0 8372 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9108 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_96
timestamp 1604681595
transform 1 0 9936 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_104
timestamp 1604681595
transform 1 0 10672 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13984 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_132
timestamp 1604681595
transform 1 0 13248 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1604681595
transform 1 0 14812 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_161
timestamp 1604681595
transform 1 0 15916 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_165
timestamp 1604681595
transform 1 0 16284 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19964 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1604681595
transform 1 0 18860 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_214
timestamp 1604681595
transform 1 0 20792 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1604681595
transform 1 0 21528 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 2852 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1932 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_11
timestamp 1604681595
transform 1 0 2116 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 3220 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_36
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4968 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_48
timestamp 1604681595
transform 1 0 5520 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_60
timestamp 1604681595
transform 1 0 6624 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 7636 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8740 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_6_72
timestamp 1604681595
transform 1 0 7728 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1604681595
transform 1 0 7544 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_75
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9752 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_84
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_103
timestamp 1604681595
transform 1 0 10580 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_99
timestamp 1604681595
transform 1 0 10212 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 11316 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10948 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1604681595
transform 1 0 11500 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1604681595
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 14352 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1604681595
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_127
timestamp 1604681595
transform 1 0 12788 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_133
timestamp 1604681595
transform 1 0 13340 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_145
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_132
timestamp 1604681595
transform 1 0 13248 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_163
timestamp 1604681595
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_153
timestamp 1604681595
transform 1 0 15180 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_165
timestamp 1604681595
transform 1 0 16284 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_175
timestamp 1604681595
transform 1 0 17204 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_187
timestamp 1604681595
transform 1 0 18308 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20056 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19044 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18400 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_204
timestamp 1604681595
transform 1 0 19872 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_197
timestamp 1604681595
transform 1 0 19228 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_205
timestamp 1604681595
transform 1 0 19964 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1604681595
transform 1 0 20884 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2208 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_11
timestamp 1604681595
transform 1 0 2116 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_18
timestamp 1604681595
transform 1 0 2760 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 4692 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1604681595
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_38
timestamp 1604681595
transform 1 0 4600 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_48
timestamp 1604681595
transform 1 0 5520 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1604681595
transform 1 0 6624 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6992 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_73
timestamp 1604681595
transform 1 0 7820 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1604681595
transform 1 0 11132 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_121
timestamp 1604681595
transform 1 0 12236 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12788 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_8_143
timestamp 1604681595
transform 1 0 14260 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16192 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_162
timestamp 1604681595
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1604681595
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_180
timestamp 1604681595
transform 1 0 17664 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18400 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1604681595
transform 1 0 19228 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1604681595
transform 1 0 20332 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_13
timestamp 1604681595
transform 1 0 2300 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 3036 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4876 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_30
timestamp 1604681595
transform 1 0 3864 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_38
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_50
timestamp 1604681595
transform 1 0 5704 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1604681595
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_71
timestamp 1604681595
transform 1 0 7636 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_83
timestamp 1604681595
transform 1 0 8740 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9200 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_87
timestamp 1604681595
transform 1 0 9108 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_97
timestamp 1604681595
transform 1 0 10028 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14260 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12696 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_152
timestamp 1604681595
transform 1 0 15088 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_164
timestamp 1604681595
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_175
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19320 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_9_190
timestamp 1604681595
transform 1 0 18584 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_214
timestamp 1604681595
transform 1 0 20792 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1604681595
transform 1 0 21528 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_17
timestamp 1604681595
transform 1 0 2668 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_40
timestamp 1604681595
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4968 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1604681595
transform 1 0 5796 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8280 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_76
timestamp 1604681595
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12328 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_114
timestamp 1604681595
transform 1 0 11592 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_138
timestamp 1604681595
transform 1 0 13800 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1604681595
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_170
timestamp 1604681595
transform 1 0 16744 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_187
timestamp 1604681595
transform 1 0 18308 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1604681595
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_206
timestamp 1604681595
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_13
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3128 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_21
timestamp 1604681595
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_38
timestamp 1604681595
transform 1 0 4600 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5336 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_52
timestamp 1604681595
transform 1 0 5888 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1604681595
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_71
timestamp 1604681595
transform 1 0 7636 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_82
timestamp 1604681595
transform 1 0 8648 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9384 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_106
timestamp 1604681595
transform 1 0 10856 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 13800 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_129
timestamp 1604681595
transform 1 0 12972 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_137
timestamp 1604681595
transform 1 0 13708 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_154
timestamp 1604681595
transform 1 0 15272 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1604681595
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_188
timestamp 1604681595
transform 1 0 18400 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_212
timestamp 1604681595
transform 1 0 20608 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_36
timestamp 1604681595
transform 1 0 4416 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_12_60
timestamp 1604681595
transform 1 0 6624 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 7728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_109
timestamp 1604681595
transform 1 0 11132 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13432 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_126
timestamp 1604681595
transform 1 0 12696 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_143
timestamp 1604681595
transform 1 0 14260 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_158
timestamp 1604681595
transform 1 0 15640 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 16468 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_12_183
timestamp 1604681595
transform 1 0 17940 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_195
timestamp 1604681595
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_206
timestamp 1604681595
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1472 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2208 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_20
timestamp 1604681595
transform 1 0 2944 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1604681595
transform 1 0 2116 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4784 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3680 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_37
timestamp 1604681595
transform 1 0 4508 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_21
timestamp 1604681595
transform 1 0 3036 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7084 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7728 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1604681595
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1604681595
transform 1 0 6992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_81
timestamp 1604681595
transform 1 0 8556 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10396 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_88
timestamp 1604681595
transform 1 0 9200 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_100
timestamp 1604681595
transform 1 0 10304 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_89
timestamp 1604681595
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12604 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12604 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 12328 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_112
timestamp 1604681595
transform 1 0 11408 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_110
timestamp 1604681595
transform 1 0 11224 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 14168 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13892 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_13_131
timestamp 1604681595
transform 1 0 13156 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_134
timestamp 1604681595
transform 1 0 13432 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16100 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_155
timestamp 1604681595
transform 1 0 15364 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_162
timestamp 1604681595
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_172
timestamp 1604681595
transform 1 0 16928 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_180
timestamp 1604681595
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_179
timestamp 1604681595
transform 1 0 17572 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_187
timestamp 1604681595
transform 1 0 18308 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_200
timestamp 1604681595
transform 1 0 19504 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_206
timestamp 1604681595
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_214
timestamp 1604681595
transform 1 0 20792 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_222
timestamp 1604681595
transform 1 0 21528 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1656 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3220 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 4876 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_32
timestamp 1604681595
transform 1 0 4048 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_40
timestamp 1604681595
transform 1 0 4784 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7268 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1604681595
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_76
timestamp 1604681595
transform 1 0 8096 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8832 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_100
timestamp 1604681595
transform 1 0 10304 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15548 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_149
timestamp 1604681595
transform 1 0 14812 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_166
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 17112 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_177
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19412 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_190
timestamp 1604681595
transform 1 0 18584 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_198
timestamp 1604681595
transform 1 0 19320 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1604681595
transform 1 0 20884 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_6
timestamp 1604681595
transform 1 0 1656 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_38
timestamp 1604681595
transform 1 0 4600 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5336 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_62
timestamp 1604681595
transform 1 0 6808 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7544 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_79
timestamp 1604681595
transform 1 0 8372 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10488 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 1604681595
transform 1 0 10396 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12328 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 1604681595
transform 1 0 13156 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_163
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 17296 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_175
timestamp 1604681595
transform 1 0 17204 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_192
timestamp 1604681595
transform 1 0 18768 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2208 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_11
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 3772 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_21
timestamp 1604681595
transform 1 0 3036 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_38
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5428 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_46
timestamp 1604681595
transform 1 0 5336 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6992 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_80
timestamp 1604681595
transform 1 0 8464 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9292 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1604681595
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1604681595
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_139
timestamp 1604681595
transform 1 0 13892 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 14628 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_156
timestamp 1604681595
transform 1 0 15456 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_164
timestamp 1604681595
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1604681595
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_193
timestamp 1604681595
transform 1 0 18860 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_210
timestamp 1604681595
transform 1 0 20424 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_222
timestamp 1604681595
transform 1 0 21528 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2208 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp 1604681595
transform 1 0 2116 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_21
timestamp 1604681595
transform 1 0 3036 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_40
timestamp 1604681595
transform 1 0 4784 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_57
timestamp 1604681595
transform 1 0 6348 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 7728 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_69
timestamp 1604681595
transform 1 0 7452 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1604681595
transform 1 0 11132 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_121
timestamp 1604681595
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12788 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_126
timestamp 1604681595
transform 1 0 12696 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_143
timestamp 1604681595
transform 1 0 14260 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_165
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17020 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_182
timestamp 1604681595
transform 1 0 17848 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_206
timestamp 1604681595
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2852 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_11
timestamp 1604681595
transform 1 0 2116 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_35
timestamp 1604681595
transform 1 0 4324 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_41
timestamp 1604681595
transform 1 0 4876 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5612 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5060 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_52
timestamp 1604681595
transform 1 0 5888 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1604681595
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_58
timestamp 1604681595
transform 1 0 6440 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8464 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 7452 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_71
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_79
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_66
timestamp 1604681595
transform 1 0 7176 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_72
timestamp 1604681595
transform 1 0 7728 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_96
timestamp 1604681595
transform 1 0 9936 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 1604681595
transform 1 0 11500 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1604681595
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13984 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_19_132
timestamp 1604681595
transform 1 0 13248 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_126
timestamp 1604681595
transform 1 0 12696 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_143
timestamp 1604681595
transform 1 0 14260 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15732 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16100 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_149
timestamp 1604681595
transform 1 0 14812 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_157
timestamp 1604681595
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_162
timestamp 1604681595
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17664 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_172
timestamp 1604681595
transform 1 0 16928 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19320 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_19_190
timestamp 1604681595
transform 1 0 18584 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_196
timestamp 1604681595
transform 1 0 19136 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_208
timestamp 1604681595
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 1604681595
transform 1 0 20792 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_222
timestamp 1604681595
transform 1 0 21528 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_16
timestamp 1604681595
transform 1 0 2576 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3312 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_40
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 5520 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_52
timestamp 1604681595
transform 1 0 5888 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1604681595
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_78
timestamp 1604681595
transform 1 0 8280 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_95
timestamp 1604681595
transform 1 0 9844 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_103
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13984 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 15548 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1604681595
transform 1 0 14812 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_160
timestamp 1604681595
transform 1 0 15824 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18768 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_6
timestamp 1604681595
transform 1 0 1656 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_3_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1604681595
transform 1 0 4876 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6072 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_53
timestamp 1604681595
transform 1 0 5980 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8280 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_70
timestamp 1604681595
transform 1 0 7544 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_109
timestamp 1604681595
transform 1 0 11132 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_133
timestamp 1604681595
transform 1 0 13340 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16284 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_157
timestamp 1604681595
transform 1 0 15548 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_181
timestamp 1604681595
transform 1 0 17756 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 18492 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1604681595
transform 1 0 18768 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_196
timestamp 1604681595
transform 1 0 19136 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_16
timestamp 1604681595
transform 1 0 2576 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4876 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3312 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_33
timestamp 1604681595
transform 1 0 4140 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_50
timestamp 1604681595
transform 1 0 5704 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_71
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_83
timestamp 1604681595
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 8924 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_101
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12512 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_109
timestamp 1604681595
transform 1 0 11132 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_140
timestamp 1604681595
transform 1 0 13984 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14720 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16284 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_157
timestamp 1604681595
transform 1 0 15548 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_174
timestamp 1604681595
transform 1 0 17112 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1604681595
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18860 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_192
timestamp 1604681595
transform 1 0 18768 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_209
timestamp 1604681595
transform 1 0 20332 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1604681595
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1604681595
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_8
timestamp 1604681595
transform 1 0 1840 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6440 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_48
timestamp 1604681595
transform 1 0 5520 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 8648 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_74
timestamp 1604681595
transform 1 0 7912 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1604681595
transform 1 0 8924 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1604681595
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_119
timestamp 1604681595
transform 1 0 12052 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12788 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 14352 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_136
timestamp 1604681595
transform 1 0 13616 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16192 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_147
timestamp 1604681595
transform 1 0 14628 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_162
timestamp 1604681595
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_180
timestamp 1604681595
transform 1 0 17664 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1604681595
transform 1 0 18768 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_196
timestamp 1604681595
transform 1 0 19136 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1656 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_22
timestamp 1604681595
transform 1 0 3128 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_34
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_47
timestamp 1604681595
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8188 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6900 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_69
timestamp 1604681595
transform 1 0 7452 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10396 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_93
timestamp 1604681595
transform 1 0 9660 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13340 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_131
timestamp 1604681595
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_149
timestamp 1604681595
transform 1 0 14812 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_157
timestamp 1604681595
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18492 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_188
timestamp 1604681595
transform 1 0 18400 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1604681595
transform 1 0 19964 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1604681595
transform 1 0 21068 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2300 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1604681595
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_8
timestamp 1604681595
transform 1 0 1840 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_38
timestamp 1604681595
transform 1 0 4600 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_29
timestamp 1604681595
transform 1 0 3772 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5336 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_55
timestamp 1604681595
transform 1 0 6164 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_46
timestamp 1604681595
transform 1 0 5336 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_58
timestamp 1604681595
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8280 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6992 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_72
timestamp 1604681595
transform 1 0 7728 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_70
timestamp 1604681595
transform 1 0 7544 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10580 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10028 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_84
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1604681595
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_87
timestamp 1604681595
transform 1 0 9108 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_95
timestamp 1604681595
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_119
timestamp 1604681595
transform 1 0 12052 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_106
timestamp 1604681595
transform 1 0 10856 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13984 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_136
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_132
timestamp 1604681595
transform 1 0 13248 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16008 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1604681595
transform 1 0 14720 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1604681595
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_156
timestamp 1604681595
transform 1 0 15456 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_173
timestamp 1604681595
transform 1 0 17020 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_187
timestamp 1604681595
transform 1 0 18308 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19044 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18768 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_201
timestamp 1604681595
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1604681595
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_211
timestamp 1604681595
transform 1 0 20516 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_6
timestamp 1604681595
transform 1 0 1656 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4416 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6624 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_28_52
timestamp 1604681595
transform 1 0 5888 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_76
timestamp 1604681595
transform 1 0 8096 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_88
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_102
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11592 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13800 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_130
timestamp 1604681595
transform 1 0 13064 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_144
timestamp 1604681595
transform 1 0 14352 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1604681595
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_163
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17664 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_175
timestamp 1604681595
transform 1 0 17204 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_179
timestamp 1604681595
transform 1 0 17572 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_189
timestamp 1604681595
transform 1 0 18492 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_206
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_16
timestamp 1604681595
transform 1 0 2576 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 3312 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_40
timestamp 1604681595
transform 1 0 4784 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 5520 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_52
timestamp 1604681595
transform 1 0 5888 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_60
timestamp 1604681595
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_78
timestamp 1604681595
transform 1 0 8280 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9384 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_106
timestamp 1604681595
transform 1 0 10856 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_132
timestamp 1604681595
transform 1 0 13248 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1604681595
transform 1 0 14812 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_161
timestamp 1604681595
transform 1 0 15916 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_165
timestamp 1604681595
transform 1 0 16284 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_175
timestamp 1604681595
transform 1 0 17204 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18768 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_6
timestamp 1604681595
transform 1 0 1656 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1604681595
transform 1 0 4876 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_30_53
timestamp 1604681595
transform 1 0 5980 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_65
timestamp 1604681595
transform 1 0 7084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_82
timestamp 1604681595
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10212 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11776 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_108
timestamp 1604681595
transform 1 0 11040 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_132
timestamp 1604681595
transform 1 0 13248 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_140
timestamp 1604681595
transform 1 0 13984 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_145
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16284 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_157
timestamp 1604681595
transform 1 0 15548 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_181
timestamp 1604681595
transform 1 0 17756 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18492 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_205
timestamp 1604681595
transform 1 0 19964 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1604681595
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_16
timestamp 1604681595
transform 1 0 2576 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3312 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_40
timestamp 1604681595
transform 1 0 4784 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 5612 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_48
timestamp 1604681595
transform 1 0 5520 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_53
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 8372 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_83
timestamp 1604681595
transform 1 0 8740 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9476 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_107
timestamp 1604681595
transform 1 0 10948 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1604681595
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13340 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_131
timestamp 1604681595
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15548 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_149
timestamp 1604681595
transform 1 0 14812 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_173
timestamp 1604681595
transform 1 0 17020 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18860 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_192
timestamp 1604681595
transform 1 0 18768 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_202
timestamp 1604681595
transform 1 0 19688 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_210
timestamp 1604681595
transform 1 0 20424 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_215
timestamp 1604681595
transform 1 0 20884 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_6
timestamp 1604681595
transform 1 0 1656 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4324 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5888 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_61
timestamp 1604681595
transform 1 0 6716 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_73
timestamp 1604681595
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_109
timestamp 1604681595
transform 1 0 11132 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13432 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_126
timestamp 1604681595
transform 1 0 12696 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_143
timestamp 1604681595
transform 1 0 14260 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_160
timestamp 1604681595
transform 1 0 15824 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 18216 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16652 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_168
timestamp 1604681595
transform 1 0 16560 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_189
timestamp 1604681595
transform 1 0 18492 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_6
timestamp 1604681595
transform 1 0 1656 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_23
timestamp 1604681595
transform 1 0 3220 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_35
timestamp 1604681595
transform 1 0 4324 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5060 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_52
timestamp 1604681595
transform 1 0 5888 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_60
timestamp 1604681595
transform 1 0 6624 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 6992 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8096 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_33_63
timestamp 1604681595
transform 1 0 6900 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_68
timestamp 1604681595
transform 1 0 7360 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10672 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_85
timestamp 1604681595
transform 1 0 8924 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_94
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_102
timestamp 1604681595
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12604 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1604681595
transform 1 0 11500 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_121
timestamp 1604681595
transform 1 0 12236 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 14260 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_134
timestamp 1604681595
transform 1 0 13432 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_142
timestamp 1604681595
transform 1 0 14168 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 15548 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_147
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_156
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_161
timestamp 1604681595
transform 1 0 15916 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16652 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_178
timestamp 1604681595
transform 1 0 17480 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_187
timestamp 1604681595
transform 1 0 18308 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18952 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_33_193
timestamp 1604681595
transform 1 0 18860 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_203
timestamp 1604681595
transform 1 0 19780 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1604681595
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 130 592
<< labels >>
rlabel metal2 s 16118 0 16174 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 202 22520 258 23000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 20718 0 20774 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 22742 22520 22798 23000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 ccff_head
port 4 nsew default input
rlabel metal2 s 11518 0 11574 480 6 ccff_tail
port 5 nsew default tristate
rlabel metal3 s 0 3136 480 3256 6 chanx_left_in[0]
port 6 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[10]
port 7 nsew default input
rlabel metal3 s 0 8576 480 8696 6 chanx_left_in[11]
port 8 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[12]
port 9 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[13]
port 10 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[14]
port 11 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[15]
port 12 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[16]
port 13 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_left_in[17]
port 14 nsew default input
rlabel metal3 s 0 12112 480 12232 6 chanx_left_in[18]
port 15 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[19]
port 16 nsew default input
rlabel metal3 s 0 3544 480 3664 6 chanx_left_in[1]
port 17 nsew default input
rlabel metal3 s 0 4088 480 4208 6 chanx_left_in[2]
port 18 nsew default input
rlabel metal3 s 0 4632 480 4752 6 chanx_left_in[3]
port 19 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[4]
port 20 nsew default input
rlabel metal3 s 0 5584 480 5704 6 chanx_left_in[5]
port 21 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[6]
port 22 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[7]
port 23 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[8]
port 24 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[9]
port 25 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_out[0]
port 26 nsew default tristate
rlabel metal3 s 0 18096 480 18216 6 chanx_left_out[10]
port 27 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[11]
port 28 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[12]
port 29 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[13]
port 30 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[14]
port 31 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[15]
port 32 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 33 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[17]
port 34 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 35 nsew default tristate
rlabel metal3 s 0 22584 480 22704 6 chanx_left_out[19]
port 36 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[1]
port 37 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[2]
port 38 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 chanx_left_out[4]
port 40 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[5]
port 41 nsew default tristate
rlabel metal3 s 0 16056 480 16176 6 chanx_left_out[6]
port 42 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[7]
port 43 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chanx_left_out[8]
port 44 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 chanx_left_out[9]
port 45 nsew default tristate
rlabel metal3 s 22520 3136 23000 3256 6 chanx_right_in[0]
port 46 nsew default input
rlabel metal3 s 22520 8032 23000 8152 6 chanx_right_in[10]
port 47 nsew default input
rlabel metal3 s 22520 8576 23000 8696 6 chanx_right_in[11]
port 48 nsew default input
rlabel metal3 s 22520 9120 23000 9240 6 chanx_right_in[12]
port 49 nsew default input
rlabel metal3 s 22520 9528 23000 9648 6 chanx_right_in[13]
port 50 nsew default input
rlabel metal3 s 22520 10072 23000 10192 6 chanx_right_in[14]
port 51 nsew default input
rlabel metal3 s 22520 10616 23000 10736 6 chanx_right_in[15]
port 52 nsew default input
rlabel metal3 s 22520 11024 23000 11144 6 chanx_right_in[16]
port 53 nsew default input
rlabel metal3 s 22520 11568 23000 11688 6 chanx_right_in[17]
port 54 nsew default input
rlabel metal3 s 22520 12112 23000 12232 6 chanx_right_in[18]
port 55 nsew default input
rlabel metal3 s 22520 12520 23000 12640 6 chanx_right_in[19]
port 56 nsew default input
rlabel metal3 s 22520 3544 23000 3664 6 chanx_right_in[1]
port 57 nsew default input
rlabel metal3 s 22520 4088 23000 4208 6 chanx_right_in[2]
port 58 nsew default input
rlabel metal3 s 22520 4632 23000 4752 6 chanx_right_in[3]
port 59 nsew default input
rlabel metal3 s 22520 5040 23000 5160 6 chanx_right_in[4]
port 60 nsew default input
rlabel metal3 s 22520 5584 23000 5704 6 chanx_right_in[5]
port 61 nsew default input
rlabel metal3 s 22520 6128 23000 6248 6 chanx_right_in[6]
port 62 nsew default input
rlabel metal3 s 22520 6536 23000 6656 6 chanx_right_in[7]
port 63 nsew default input
rlabel metal3 s 22520 7080 23000 7200 6 chanx_right_in[8]
port 64 nsew default input
rlabel metal3 s 22520 7624 23000 7744 6 chanx_right_in[9]
port 65 nsew default input
rlabel metal3 s 22520 13064 23000 13184 6 chanx_right_out[0]
port 66 nsew default tristate
rlabel metal3 s 22520 18096 23000 18216 6 chanx_right_out[10]
port 67 nsew default tristate
rlabel metal3 s 22520 18504 23000 18624 6 chanx_right_out[11]
port 68 nsew default tristate
rlabel metal3 s 22520 19048 23000 19168 6 chanx_right_out[12]
port 69 nsew default tristate
rlabel metal3 s 22520 19592 23000 19712 6 chanx_right_out[13]
port 70 nsew default tristate
rlabel metal3 s 22520 20000 23000 20120 6 chanx_right_out[14]
port 71 nsew default tristate
rlabel metal3 s 22520 20544 23000 20664 6 chanx_right_out[15]
port 72 nsew default tristate
rlabel metal3 s 22520 21088 23000 21208 6 chanx_right_out[16]
port 73 nsew default tristate
rlabel metal3 s 22520 21496 23000 21616 6 chanx_right_out[17]
port 74 nsew default tristate
rlabel metal3 s 22520 22040 23000 22160 6 chanx_right_out[18]
port 75 nsew default tristate
rlabel metal3 s 22520 22584 23000 22704 6 chanx_right_out[19]
port 76 nsew default tristate
rlabel metal3 s 22520 13608 23000 13728 6 chanx_right_out[1]
port 77 nsew default tristate
rlabel metal3 s 22520 14016 23000 14136 6 chanx_right_out[2]
port 78 nsew default tristate
rlabel metal3 s 22520 14560 23000 14680 6 chanx_right_out[3]
port 79 nsew default tristate
rlabel metal3 s 22520 15104 23000 15224 6 chanx_right_out[4]
port 80 nsew default tristate
rlabel metal3 s 22520 15512 23000 15632 6 chanx_right_out[5]
port 81 nsew default tristate
rlabel metal3 s 22520 16056 23000 16176 6 chanx_right_out[6]
port 82 nsew default tristate
rlabel metal3 s 22520 16600 23000 16720 6 chanx_right_out[7]
port 83 nsew default tristate
rlabel metal3 s 22520 17008 23000 17128 6 chanx_right_out[8]
port 84 nsew default tristate
rlabel metal3 s 22520 17552 23000 17672 6 chanx_right_out[9]
port 85 nsew default tristate
rlabel metal2 s 4342 22520 4398 23000 6 chany_top_in[0]
port 86 nsew default input
rlabel metal2 s 8942 22520 8998 23000 6 chany_top_in[10]
port 87 nsew default input
rlabel metal2 s 9402 22520 9458 23000 6 chany_top_in[11]
port 88 nsew default input
rlabel metal2 s 9862 22520 9918 23000 6 chany_top_in[12]
port 89 nsew default input
rlabel metal2 s 10322 22520 10378 23000 6 chany_top_in[13]
port 90 nsew default input
rlabel metal2 s 10782 22520 10838 23000 6 chany_top_in[14]
port 91 nsew default input
rlabel metal2 s 11242 22520 11298 23000 6 chany_top_in[15]
port 92 nsew default input
rlabel metal2 s 11702 22520 11758 23000 6 chany_top_in[16]
port 93 nsew default input
rlabel metal2 s 12162 22520 12218 23000 6 chany_top_in[17]
port 94 nsew default input
rlabel metal2 s 12622 22520 12678 23000 6 chany_top_in[18]
port 95 nsew default input
rlabel metal2 s 13082 22520 13138 23000 6 chany_top_in[19]
port 96 nsew default input
rlabel metal2 s 4802 22520 4858 23000 6 chany_top_in[1]
port 97 nsew default input
rlabel metal2 s 5262 22520 5318 23000 6 chany_top_in[2]
port 98 nsew default input
rlabel metal2 s 5722 22520 5778 23000 6 chany_top_in[3]
port 99 nsew default input
rlabel metal2 s 6182 22520 6238 23000 6 chany_top_in[4]
port 100 nsew default input
rlabel metal2 s 6642 22520 6698 23000 6 chany_top_in[5]
port 101 nsew default input
rlabel metal2 s 7102 22520 7158 23000 6 chany_top_in[6]
port 102 nsew default input
rlabel metal2 s 7562 22520 7618 23000 6 chany_top_in[7]
port 103 nsew default input
rlabel metal2 s 8022 22520 8078 23000 6 chany_top_in[8]
port 104 nsew default input
rlabel metal2 s 8482 22520 8538 23000 6 chany_top_in[9]
port 105 nsew default input
rlabel metal2 s 13542 22520 13598 23000 6 chany_top_out[0]
port 106 nsew default tristate
rlabel metal2 s 18142 22520 18198 23000 6 chany_top_out[10]
port 107 nsew default tristate
rlabel metal2 s 18602 22520 18658 23000 6 chany_top_out[11]
port 108 nsew default tristate
rlabel metal2 s 19062 22520 19118 23000 6 chany_top_out[12]
port 109 nsew default tristate
rlabel metal2 s 19522 22520 19578 23000 6 chany_top_out[13]
port 110 nsew default tristate
rlabel metal2 s 19982 22520 20038 23000 6 chany_top_out[14]
port 111 nsew default tristate
rlabel metal2 s 20442 22520 20498 23000 6 chany_top_out[15]
port 112 nsew default tristate
rlabel metal2 s 20902 22520 20958 23000 6 chany_top_out[16]
port 113 nsew default tristate
rlabel metal2 s 21362 22520 21418 23000 6 chany_top_out[17]
port 114 nsew default tristate
rlabel metal2 s 21822 22520 21878 23000 6 chany_top_out[18]
port 115 nsew default tristate
rlabel metal2 s 22282 22520 22338 23000 6 chany_top_out[19]
port 116 nsew default tristate
rlabel metal2 s 14002 22520 14058 23000 6 chany_top_out[1]
port 117 nsew default tristate
rlabel metal2 s 14462 22520 14518 23000 6 chany_top_out[2]
port 118 nsew default tristate
rlabel metal2 s 14922 22520 14978 23000 6 chany_top_out[3]
port 119 nsew default tristate
rlabel metal2 s 15382 22520 15438 23000 6 chany_top_out[4]
port 120 nsew default tristate
rlabel metal2 s 15842 22520 15898 23000 6 chany_top_out[5]
port 121 nsew default tristate
rlabel metal2 s 16302 22520 16358 23000 6 chany_top_out[6]
port 122 nsew default tristate
rlabel metal2 s 16762 22520 16818 23000 6 chany_top_out[7]
port 123 nsew default tristate
rlabel metal2 s 17222 22520 17278 23000 6 chany_top_out[8]
port 124 nsew default tristate
rlabel metal2 s 17682 22520 17738 23000 6 chany_top_out[9]
port 125 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 left_bottom_grid_pin_11_
port 126 nsew default input
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_1_
port 127 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_3_
port 128 nsew default input
rlabel metal3 s 0 1096 480 1216 6 left_bottom_grid_pin_5_
port 129 nsew default input
rlabel metal3 s 0 1640 480 1760 6 left_bottom_grid_pin_7_
port 130 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_9_
port 131 nsew default input
rlabel metal2 s 2318 0 2374 480 6 prog_clk
port 132 nsew default input
rlabel metal3 s 22520 2592 23000 2712 6 right_bottom_grid_pin_11_
port 133 nsew default input
rlabel metal3 s 22520 144 23000 264 6 right_bottom_grid_pin_1_
port 134 nsew default input
rlabel metal3 s 22520 552 23000 672 6 right_bottom_grid_pin_3_
port 135 nsew default input
rlabel metal3 s 22520 1096 23000 1216 6 right_bottom_grid_pin_5_
port 136 nsew default input
rlabel metal3 s 22520 1640 23000 1760 6 right_bottom_grid_pin_7_
port 137 nsew default input
rlabel metal3 s 22520 2048 23000 2168 6 right_bottom_grid_pin_9_
port 138 nsew default input
rlabel metal2 s 662 22520 718 23000 6 top_left_grid_pin_42_
port 139 nsew default input
rlabel metal2 s 1122 22520 1178 23000 6 top_left_grid_pin_43_
port 140 nsew default input
rlabel metal2 s 1582 22520 1638 23000 6 top_left_grid_pin_44_
port 141 nsew default input
rlabel metal2 s 2042 22520 2098 23000 6 top_left_grid_pin_45_
port 142 nsew default input
rlabel metal2 s 2502 22520 2558 23000 6 top_left_grid_pin_46_
port 143 nsew default input
rlabel metal2 s 2962 22520 3018 23000 6 top_left_grid_pin_47_
port 144 nsew default input
rlabel metal2 s 3422 22520 3478 23000 6 top_left_grid_pin_48_
port 145 nsew default input
rlabel metal2 s 3882 22520 3938 23000 6 top_left_grid_pin_49_
port 146 nsew default input
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 147 nsew default input
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 148 nsew default input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
