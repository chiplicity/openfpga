VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_left
  CLASS BLOCK ;
  FOREIGN grid_io_left ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 137.600 14.170 140.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 2.400 43.480 ;
    END
  END address[3]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END enable
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 9.560 140.000 10.160 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 41.490 137.600 41.770 140.000 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 29.280 140.000 29.880 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 49.000 140.000 49.600 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 2.400 61.160 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 2.400 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 2.400 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN right_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 2.400 ;
    END
  END right_width_0_height_0__pin_0_
  PIN right_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 2.400 113.520 ;
    END
  END right_width_0_height_0__pin_10_
  PIN right_width_0_height_0__pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.610 137.600 97.890 140.000 ;
    END
  END right_width_0_height_0__pin_11_
  PIN right_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 129.240 140.000 129.840 ;
    END
  END right_width_0_height_0__pin_12_
  PIN right_width_0_height_0__pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.400 131.200 ;
    END
  END right_width_0_height_0__pin_13_
  PIN right_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 2.400 ;
    END
  END right_width_0_height_0__pin_14_
  PIN right_width_0_height_0__pin_15_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 125.670 137.600 125.950 140.000 ;
    END
  END right_width_0_height_0__pin_15_
  PIN right_width_0_height_0__pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 2.400 ;
    END
  END right_width_0_height_0__pin_1_
  PIN right_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END right_width_0_height_0__pin_2_
  PIN right_width_0_height_0__pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.400 78.840 ;
    END
  END right_width_0_height_0__pin_3_
  PIN right_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END right_width_0_height_0__pin_4_
  PIN right_width_0_height_0__pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END right_width_0_height_0__pin_5_
  PIN right_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 89.120 140.000 89.720 ;
    END
  END right_width_0_height_0__pin_6_
  PIN right_width_0_height_0__pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 2.400 ;
    END
  END right_width_0_height_0__pin_7_
  PIN right_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 2.400 ;
    END
  END right_width_0_height_0__pin_8_
  PIN right_width_0_height_0__pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 109.520 140.000 110.120 ;
    END
  END right_width_0_height_0__pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.530 10.640 134.320 128.080 ;
      LAYER met2 ;
        RECT 0.550 137.320 13.610 137.770 ;
        RECT 14.450 137.320 41.210 137.770 ;
        RECT 42.050 137.320 69.270 137.770 ;
        RECT 70.110 137.320 97.330 137.770 ;
        RECT 98.170 137.320 122.925 137.770 ;
        RECT 0.550 2.680 122.925 137.320 ;
        RECT 0.550 0.270 6.710 2.680 ;
        RECT 7.550 0.270 20.510 2.680 ;
        RECT 21.350 0.270 34.310 2.680 ;
        RECT 35.150 0.270 48.570 2.680 ;
        RECT 49.410 0.270 62.370 2.680 ;
        RECT 63.210 0.270 76.630 2.680 ;
        RECT 77.470 0.270 90.430 2.680 ;
        RECT 91.270 0.270 104.230 2.680 ;
        RECT 105.070 0.270 118.490 2.680 ;
        RECT 119.330 0.270 122.925 2.680 ;
      LAYER met3 ;
        RECT 0.310 113.920 122.985 128.005 ;
        RECT 2.800 112.520 122.985 113.920 ;
        RECT 0.310 96.240 122.985 112.520 ;
        RECT 2.800 94.840 122.985 96.240 ;
        RECT 0.310 79.240 122.985 94.840 ;
        RECT 2.800 77.840 122.985 79.240 ;
        RECT 0.310 61.560 122.985 77.840 ;
        RECT 2.800 60.160 122.985 61.560 ;
        RECT 0.310 43.880 122.985 60.160 ;
        RECT 2.800 42.480 122.985 43.880 ;
        RECT 0.310 26.200 122.985 42.480 ;
        RECT 2.800 24.800 122.985 26.200 ;
        RECT 0.310 10.715 122.985 24.800 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END grid_io_left
END LIBRARY

