magic
tech sky130A
magscale 1 2
timestamp 1605122293
<< locali >>
rect 8953 25143 8987 25313
rect 11805 25211 11839 25381
rect 11897 25279 11931 25449
rect 15393 21471 15427 21641
rect 3709 20791 3743 20961
rect 23121 20927 23155 21097
rect 25329 18683 25363 18921
rect 10241 18207 10275 18309
rect 18613 16643 18647 16745
rect 20545 16575 20579 16745
rect 2697 14807 2731 15113
rect 6837 14875 6871 15113
rect 24961 15011 24995 15113
rect 3249 14263 3283 14569
<< viali >>
rect 2697 25449 2731 25483
rect 8769 25449 8803 25483
rect 10517 25449 10551 25483
rect 11621 25449 11655 25483
rect 11897 25449 11931 25483
rect 24777 25449 24811 25483
rect 8125 25381 8159 25415
rect 11805 25381 11839 25415
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 4077 25313 4111 25347
rect 5733 25313 5767 25347
rect 7481 25313 7515 25347
rect 8585 25313 8619 25347
rect 8953 25313 8987 25347
rect 10333 25313 10367 25347
rect 11462 25313 11496 25347
rect 4261 25177 4295 25211
rect 5917 25177 5951 25211
rect 7665 25177 7699 25211
rect 20085 25381 20119 25415
rect 22753 25381 22787 25415
rect 13001 25313 13035 25347
rect 13093 25313 13127 25347
rect 14289 25313 14323 25347
rect 16037 25313 16071 25347
rect 17233 25313 17267 25347
rect 18889 25313 18923 25347
rect 21189 25313 21223 25347
rect 22477 25313 22511 25347
rect 24593 25313 24627 25347
rect 11897 25245 11931 25279
rect 13185 25245 13219 25279
rect 16129 25245 16163 25279
rect 16313 25245 16347 25279
rect 18981 25245 19015 25279
rect 19165 25245 19199 25279
rect 21465 25245 21499 25279
rect 11805 25177 11839 25211
rect 12633 25177 12667 25211
rect 14473 25177 14507 25211
rect 1593 25109 1627 25143
rect 6285 25109 6319 25143
rect 7205 25109 7239 25143
rect 8953 25109 8987 25143
rect 9229 25109 9263 25143
rect 10057 25109 10091 25143
rect 12081 25109 12115 25143
rect 13737 25109 13771 25143
rect 14013 25109 14047 25143
rect 14841 25109 14875 25143
rect 15301 25109 15335 25143
rect 15669 25109 15703 25143
rect 16681 25109 16715 25143
rect 17049 25109 17083 25143
rect 17693 25109 17727 25143
rect 18153 25109 18187 25143
rect 18521 25109 18555 25143
rect 19533 25109 19567 25143
rect 2697 24905 2731 24939
rect 3801 24905 3835 24939
rect 4905 24905 4939 24939
rect 17785 24905 17819 24939
rect 18153 24905 18187 24939
rect 22937 24905 22971 24939
rect 24409 24905 24443 24939
rect 11897 24837 11931 24871
rect 6653 24769 6687 24803
rect 7389 24769 7423 24803
rect 7573 24769 7607 24803
rect 9045 24769 9079 24803
rect 9505 24769 9539 24803
rect 11253 24769 11287 24803
rect 13645 24769 13679 24803
rect 16405 24769 16439 24803
rect 18613 24769 18647 24803
rect 18705 24769 18739 24803
rect 19809 24769 19843 24803
rect 20637 24769 20671 24803
rect 21005 24769 21039 24803
rect 1409 24701 1443 24735
rect 2053 24701 2087 24735
rect 2513 24701 2547 24735
rect 3157 24701 3191 24735
rect 3617 24701 3651 24735
rect 4261 24701 4295 24735
rect 4721 24701 4755 24735
rect 6285 24701 6319 24735
rect 8309 24701 8343 24735
rect 8861 24701 8895 24735
rect 11069 24701 11103 24735
rect 13369 24701 13403 24735
rect 20361 24701 20395 24735
rect 22201 24701 22235 24735
rect 24593 24701 24627 24735
rect 25145 24701 25179 24735
rect 5825 24633 5859 24667
rect 8033 24633 8067 24667
rect 10057 24633 10091 24667
rect 13461 24633 13495 24667
rect 14381 24633 14415 24667
rect 15301 24633 15335 24667
rect 20453 24633 20487 24667
rect 22477 24633 22511 24667
rect 1593 24565 1627 24599
rect 2421 24565 2455 24599
rect 3525 24565 3559 24599
rect 5273 24565 5307 24599
rect 6929 24565 6963 24599
rect 7297 24565 7331 24599
rect 8493 24565 8527 24599
rect 8953 24565 8987 24599
rect 9965 24565 9999 24599
rect 10609 24565 10643 24599
rect 10977 24565 11011 24599
rect 12173 24565 12207 24599
rect 12817 24565 12851 24599
rect 13001 24565 13035 24599
rect 14105 24565 14139 24599
rect 14841 24565 14875 24599
rect 15577 24565 15611 24599
rect 15761 24565 15795 24599
rect 16129 24565 16163 24599
rect 16221 24565 16255 24599
rect 16773 24565 16807 24599
rect 17417 24565 17451 24599
rect 18521 24565 18555 24599
rect 19165 24565 19199 24599
rect 19993 24565 20027 24599
rect 21373 24565 21407 24599
rect 22109 24565 22143 24599
rect 24777 24565 24811 24599
rect 4261 24361 4295 24395
rect 7849 24361 7883 24395
rect 8217 24361 8251 24395
rect 9229 24361 9263 24395
rect 9689 24361 9723 24395
rect 10057 24361 10091 24395
rect 11253 24361 11287 24395
rect 13645 24361 13679 24395
rect 14657 24361 14691 24395
rect 15485 24361 15519 24395
rect 16589 24361 16623 24395
rect 18061 24361 18095 24395
rect 19533 24361 19567 24395
rect 19901 24361 19935 24395
rect 20269 24361 20303 24395
rect 25513 24361 25547 24395
rect 5908 24293 5942 24327
rect 8309 24293 8343 24327
rect 10149 24293 10183 24327
rect 16865 24293 16899 24327
rect 1409 24225 1443 24259
rect 2513 24225 2547 24259
rect 4077 24225 4111 24259
rect 5641 24225 5675 24259
rect 12081 24225 12115 24259
rect 13737 24225 13771 24259
rect 15853 24225 15887 24259
rect 17601 24225 17635 24259
rect 18429 24225 18463 24259
rect 19717 24225 19751 24259
rect 21281 24225 21315 24259
rect 22845 24225 22879 24259
rect 24041 24225 24075 24259
rect 25329 24225 25363 24259
rect 3065 24157 3099 24191
rect 8401 24157 8435 24191
rect 10241 24157 10275 24191
rect 12173 24157 12207 24191
rect 12265 24157 12299 24191
rect 13921 24157 13955 24191
rect 14381 24157 14415 24191
rect 15945 24157 15979 24191
rect 16037 24157 16071 24191
rect 17049 24157 17083 24191
rect 18521 24157 18555 24191
rect 18705 24157 18739 24191
rect 21373 24157 21407 24191
rect 21557 24157 21591 24191
rect 22937 24157 22971 24191
rect 23029 24157 23063 24191
rect 24225 24157 24259 24191
rect 7297 24089 7331 24123
rect 11529 24089 11563 24123
rect 20637 24089 20671 24123
rect 21925 24089 21959 24123
rect 1593 24021 1627 24055
rect 1961 24021 1995 24055
rect 2697 24021 2731 24055
rect 4905 24021 4939 24055
rect 5273 24021 5307 24055
rect 7021 24021 7055 24055
rect 7757 24021 7791 24055
rect 8953 24021 8987 24055
rect 10701 24021 10735 24055
rect 11713 24021 11747 24055
rect 13001 24021 13035 24055
rect 13277 24021 13311 24055
rect 15117 24021 15151 24055
rect 17969 24021 18003 24055
rect 19165 24021 19199 24055
rect 20913 24021 20947 24055
rect 22293 24021 22327 24055
rect 22477 24021 22511 24055
rect 23765 24021 23799 24055
rect 3157 23817 3191 23851
rect 3801 23817 3835 23851
rect 4629 23817 4663 23851
rect 8309 23817 8343 23851
rect 11069 23817 11103 23851
rect 11437 23817 11471 23851
rect 12265 23817 12299 23851
rect 15117 23817 15151 23851
rect 16865 23817 16899 23851
rect 17877 23817 17911 23851
rect 19441 23817 19475 23851
rect 22109 23817 22143 23851
rect 25421 23817 25455 23851
rect 25789 23817 25823 23851
rect 6837 23749 6871 23783
rect 8401 23749 8435 23783
rect 10057 23749 10091 23783
rect 23673 23749 23707 23783
rect 5641 23681 5675 23715
rect 5825 23681 5859 23715
rect 7297 23681 7331 23715
rect 7389 23681 7423 23715
rect 8953 23681 8987 23715
rect 9781 23681 9815 23715
rect 10701 23681 10735 23715
rect 15209 23681 15243 23715
rect 20361 23681 20395 23715
rect 24225 23681 24259 23715
rect 1409 23613 1443 23647
rect 2421 23613 2455 23647
rect 2513 23613 2547 23647
rect 3617 23613 3651 23647
rect 4261 23613 4295 23647
rect 5549 23613 5583 23647
rect 7941 23613 7975 23647
rect 8769 23613 8803 23647
rect 10425 23613 10459 23647
rect 12449 23613 12483 23647
rect 18061 23613 18095 23647
rect 25237 23613 25271 23647
rect 5089 23545 5123 23579
rect 8861 23545 8895 23579
rect 11897 23545 11931 23579
rect 12694 23545 12728 23579
rect 15476 23545 15510 23579
rect 18306 23545 18340 23579
rect 20606 23545 20640 23579
rect 23029 23545 23063 23579
rect 24685 23545 24719 23579
rect 1593 23477 1627 23511
rect 1961 23477 1995 23511
rect 2697 23477 2731 23511
rect 3525 23477 3559 23511
rect 5181 23477 5215 23511
rect 6285 23477 6319 23511
rect 6561 23477 6595 23511
rect 7205 23477 7239 23511
rect 10517 23477 10551 23511
rect 13829 23477 13863 23511
rect 14197 23477 14231 23511
rect 14565 23477 14599 23511
rect 16589 23477 16623 23511
rect 17509 23477 17543 23511
rect 19717 23477 19751 23511
rect 20269 23477 20303 23511
rect 21741 23477 21775 23511
rect 22385 23477 22419 23511
rect 22569 23477 22603 23511
rect 23489 23477 23523 23511
rect 24041 23477 24075 23511
rect 24133 23477 24167 23511
rect 25053 23477 25087 23511
rect 2513 23273 2547 23307
rect 4261 23273 4295 23307
rect 7297 23273 7331 23307
rect 9045 23273 9079 23307
rect 9505 23273 9539 23307
rect 9689 23273 9723 23307
rect 11253 23273 11287 23307
rect 12725 23273 12759 23307
rect 13369 23273 13403 23307
rect 13921 23273 13955 23307
rect 15117 23273 15151 23307
rect 15853 23273 15887 23307
rect 17693 23273 17727 23307
rect 18061 23273 18095 23307
rect 18521 23273 18555 23307
rect 19993 23273 20027 23307
rect 20453 23273 20487 23307
rect 22937 23273 22971 23307
rect 23213 23273 23247 23307
rect 23581 23273 23615 23307
rect 24225 23273 24259 23307
rect 24869 23273 24903 23307
rect 25513 23273 25547 23307
rect 3525 23205 3559 23239
rect 3893 23205 3927 23239
rect 16580 23205 16614 23239
rect 18858 23205 18892 23239
rect 21802 23205 21836 23239
rect 1685 23137 1719 23171
rect 1961 23137 1995 23171
rect 4077 23137 4111 23171
rect 4629 23137 4663 23171
rect 5181 23137 5215 23171
rect 5448 23137 5482 23171
rect 7656 23137 7690 23171
rect 10057 23137 10091 23171
rect 11612 23137 11646 23171
rect 14013 23137 14047 23171
rect 16313 23137 16347 23171
rect 18613 23137 18647 23171
rect 21557 23137 21591 23171
rect 24133 23137 24167 23171
rect 25329 23137 25363 23171
rect 2973 23069 3007 23103
rect 7389 23069 7423 23103
rect 10149 23069 10183 23103
rect 10241 23069 10275 23103
rect 11345 23069 11379 23103
rect 14105 23069 14139 23103
rect 15301 23069 15335 23103
rect 24317 23069 24351 23103
rect 2881 23001 2915 23035
rect 23765 23001 23799 23035
rect 5089 22933 5123 22967
rect 6561 22933 6595 22967
rect 6929 22933 6963 22967
rect 8769 22933 8803 22967
rect 10793 22933 10827 22967
rect 13553 22933 13587 22967
rect 14565 22933 14599 22967
rect 16221 22933 16255 22967
rect 21097 22933 21131 22967
rect 2237 22729 2271 22763
rect 5181 22729 5215 22763
rect 7849 22729 7883 22763
rect 9505 22729 9539 22763
rect 9873 22729 9907 22763
rect 10333 22729 10367 22763
rect 13553 22729 13587 22763
rect 15853 22729 15887 22763
rect 18061 22729 18095 22763
rect 19073 22729 19107 22763
rect 19901 22729 19935 22763
rect 20361 22729 20395 22763
rect 21557 22729 21591 22763
rect 22017 22729 22051 22763
rect 23029 22729 23063 22763
rect 26065 22729 26099 22763
rect 4997 22661 5031 22695
rect 6837 22661 6871 22695
rect 11345 22661 11379 22695
rect 21925 22661 21959 22695
rect 5641 22593 5675 22627
rect 5825 22593 5859 22627
rect 7481 22593 7515 22627
rect 8861 22593 8895 22627
rect 9045 22593 9079 22627
rect 10793 22593 10827 22627
rect 10885 22593 10919 22627
rect 11713 22593 11747 22627
rect 12909 22593 12943 22627
rect 13093 22593 13127 22627
rect 16865 22593 16899 22627
rect 18613 22593 18647 22627
rect 20269 22593 20303 22627
rect 21005 22593 21039 22627
rect 22661 22593 22695 22627
rect 24317 22593 24351 22627
rect 1409 22525 1443 22559
rect 1685 22525 1719 22559
rect 2697 22525 2731 22559
rect 5549 22525 5583 22559
rect 6285 22525 6319 22559
rect 8309 22525 8343 22559
rect 8769 22525 8803 22559
rect 10241 22525 10275 22559
rect 10701 22525 10735 22559
rect 12173 22525 12207 22559
rect 12817 22525 12851 22559
rect 14105 22525 14139 22559
rect 17877 22525 17911 22559
rect 18521 22525 18555 22559
rect 20821 22525 20855 22559
rect 22385 22525 22419 22559
rect 22477 22525 22511 22559
rect 24133 22525 24167 22559
rect 25329 22525 25363 22559
rect 2605 22457 2639 22491
rect 2964 22457 2998 22491
rect 4721 22457 4755 22491
rect 6653 22457 6687 22491
rect 7297 22457 7331 22491
rect 14013 22457 14047 22491
rect 14350 22457 14384 22491
rect 16773 22457 16807 22491
rect 17417 22457 17451 22491
rect 19533 22457 19567 22491
rect 20729 22457 20763 22491
rect 24777 22457 24811 22491
rect 25605 22457 25639 22491
rect 4077 22389 4111 22423
rect 7205 22389 7239 22423
rect 8401 22389 8435 22423
rect 12449 22389 12483 22423
rect 15485 22389 15519 22423
rect 16129 22389 16163 22423
rect 16313 22389 16347 22423
rect 16681 22389 16715 22423
rect 18429 22389 18463 22423
rect 23397 22389 23431 22423
rect 23765 22389 23799 22423
rect 24225 22389 24259 22423
rect 25145 22389 25179 22423
rect 2789 22185 2823 22219
rect 5457 22185 5491 22219
rect 5825 22185 5859 22219
rect 7021 22185 7055 22219
rect 7665 22185 7699 22219
rect 18061 22185 18095 22219
rect 18429 22185 18463 22219
rect 18613 22185 18647 22219
rect 20913 22185 20947 22219
rect 21281 22185 21315 22219
rect 22109 22185 22143 22219
rect 24133 22185 24167 22219
rect 11336 22117 11370 22151
rect 22477 22117 22511 22151
rect 22998 22117 23032 22151
rect 4333 22049 4367 22083
rect 8309 22049 8343 22083
rect 9689 22049 9723 22083
rect 9965 22049 9999 22083
rect 11069 22049 11103 22083
rect 12817 22049 12851 22083
rect 13645 22049 13679 22083
rect 13737 22049 13771 22083
rect 15301 22049 15335 22083
rect 16672 22049 16706 22083
rect 18981 22049 19015 22083
rect 22753 22049 22787 22083
rect 24869 22049 24903 22083
rect 24961 22049 24995 22083
rect 2881 21981 2915 22015
rect 3065 21981 3099 22015
rect 4077 21981 4111 22015
rect 7113 21981 7147 22015
rect 7297 21981 7331 22015
rect 8585 21981 8619 22015
rect 13093 21981 13127 22015
rect 13921 21981 13955 22015
rect 16405 21981 16439 22015
rect 19073 21981 19107 22015
rect 19165 21981 19199 22015
rect 21373 21981 21407 22015
rect 21465 21981 21499 22015
rect 25237 21981 25271 22015
rect 2329 21913 2363 21947
rect 6101 21913 6135 21947
rect 6653 21913 6687 21947
rect 9045 21913 9079 21947
rect 13277 21913 13311 21947
rect 14381 21913 14415 21947
rect 15485 21913 15519 21947
rect 19717 21913 19751 21947
rect 1593 21845 1627 21879
rect 2421 21845 2455 21879
rect 3433 21845 3467 21879
rect 3801 21845 3835 21879
rect 6561 21845 6595 21879
rect 8033 21845 8067 21879
rect 9413 21845 9447 21879
rect 10425 21845 10459 21879
rect 10885 21845 10919 21879
rect 12449 21845 12483 21879
rect 14657 21845 14691 21879
rect 15025 21845 15059 21879
rect 16129 21845 16163 21879
rect 17785 21845 17819 21879
rect 19993 21845 20027 21879
rect 20729 21845 20763 21879
rect 24501 21845 24535 21879
rect 2513 21641 2547 21675
rect 4169 21641 4203 21675
rect 4813 21641 4847 21675
rect 6193 21641 6227 21675
rect 8769 21641 8803 21675
rect 9137 21641 9171 21675
rect 10241 21641 10275 21675
rect 11345 21641 11379 21675
rect 12265 21641 12299 21675
rect 15393 21641 15427 21675
rect 19625 21641 19659 21675
rect 21189 21641 21223 21675
rect 22201 21641 22235 21675
rect 22845 21641 22879 21675
rect 4445 21573 4479 21607
rect 15301 21573 15335 21607
rect 1777 21505 1811 21539
rect 5457 21505 5491 21539
rect 5549 21505 5583 21539
rect 10793 21505 10827 21539
rect 11897 21505 11931 21539
rect 12725 21505 12759 21539
rect 17785 21573 17819 21607
rect 19073 21573 19107 21607
rect 16773 21505 16807 21539
rect 17509 21505 17543 21539
rect 18613 21505 18647 21539
rect 20269 21505 20303 21539
rect 21741 21505 21775 21539
rect 23489 21505 23523 21539
rect 1501 21437 1535 21471
rect 2789 21437 2823 21471
rect 5365 21437 5399 21471
rect 7389 21437 7423 21471
rect 7656 21437 7690 21471
rect 12449 21437 12483 21471
rect 13921 21437 13955 21471
rect 15393 21437 15427 21471
rect 15669 21437 15703 21471
rect 19993 21437 20027 21471
rect 23673 21437 23707 21471
rect 23940 21437 23974 21471
rect 3056 21369 3090 21403
rect 10701 21369 10735 21403
rect 14188 21369 14222 21403
rect 16589 21369 16623 21403
rect 18521 21369 18555 21403
rect 21649 21369 21683 21403
rect 25329 21369 25363 21403
rect 4997 21301 5031 21335
rect 6653 21301 6687 21335
rect 7113 21301 7147 21335
rect 9689 21301 9723 21335
rect 10057 21301 10091 21335
rect 10609 21301 10643 21335
rect 13277 21301 13311 21335
rect 13737 21301 13771 21335
rect 15945 21301 15979 21335
rect 16129 21301 16163 21335
rect 16497 21301 16531 21335
rect 18061 21301 18095 21335
rect 18429 21301 18463 21335
rect 19441 21301 19475 21335
rect 20085 21301 20119 21335
rect 20913 21301 20947 21335
rect 21557 21301 21591 21335
rect 25053 21301 25087 21335
rect 25697 21301 25731 21335
rect 2421 21097 2455 21131
rect 5181 21097 5215 21131
rect 6193 21097 6227 21131
rect 7573 21097 7607 21131
rect 8033 21097 8067 21131
rect 8401 21097 8435 21131
rect 12357 21097 12391 21131
rect 12817 21097 12851 21131
rect 13461 21097 13495 21131
rect 17233 21097 17267 21131
rect 19993 21097 20027 21131
rect 20729 21097 20763 21131
rect 21189 21097 21223 21131
rect 21557 21097 21591 21131
rect 22201 21097 22235 21131
rect 22845 21097 22879 21131
rect 23121 21097 23155 21131
rect 23213 21097 23247 21131
rect 24777 21097 24811 21131
rect 2881 21029 2915 21063
rect 3525 21029 3559 21063
rect 4537 21029 4571 21063
rect 7941 21029 7975 21063
rect 12173 21029 12207 21063
rect 15025 21029 15059 21063
rect 15669 21029 15703 21063
rect 16865 21029 16899 21063
rect 17601 21029 17635 21063
rect 18052 21029 18086 21063
rect 2329 20961 2363 20995
rect 2789 20961 2823 20995
rect 3709 20961 3743 20995
rect 4445 20961 4479 20995
rect 5457 20961 5491 20995
rect 6377 20961 6411 20995
rect 6837 20961 6871 20995
rect 10057 20961 10091 20995
rect 10324 20961 10358 20995
rect 12725 20961 12759 20995
rect 13921 20961 13955 20995
rect 16497 20961 16531 20995
rect 20177 20961 20211 20995
rect 1409 20893 1443 20927
rect 1961 20893 1995 20927
rect 3065 20893 3099 20927
rect 23653 20961 23687 20995
rect 4629 20893 4663 20927
rect 6929 20893 6963 20927
rect 7021 20893 7055 20927
rect 8493 20893 8527 20927
rect 8677 20893 8711 20927
rect 13001 20893 13035 20927
rect 14197 20893 14231 20927
rect 15761 20893 15795 20927
rect 15945 20893 15979 20927
rect 17785 20893 17819 20927
rect 22293 20893 22327 20927
rect 22477 20893 22511 20927
rect 23121 20893 23155 20927
rect 23397 20893 23431 20927
rect 3801 20825 3835 20859
rect 15301 20825 15335 20859
rect 19165 20825 19199 20859
rect 3709 20757 3743 20791
rect 4077 20757 4111 20791
rect 6101 20757 6135 20791
rect 6469 20757 6503 20791
rect 9137 20757 9171 20791
rect 9505 20757 9539 20791
rect 9965 20757 9999 20791
rect 11437 20757 11471 20791
rect 11897 20757 11931 20791
rect 13737 20757 13771 20791
rect 14749 20757 14783 20791
rect 19625 20757 19659 20791
rect 21833 20757 21867 20791
rect 25053 20757 25087 20791
rect 25421 20757 25455 20791
rect 2513 20553 2547 20587
rect 3985 20553 4019 20587
rect 5917 20553 5951 20587
rect 6561 20553 6595 20587
rect 7113 20553 7147 20587
rect 7573 20553 7607 20587
rect 11253 20553 11287 20587
rect 11989 20553 12023 20587
rect 13829 20553 13863 20587
rect 16313 20553 16347 20587
rect 23673 20553 23707 20587
rect 15485 20485 15519 20519
rect 16129 20485 16163 20519
rect 3157 20417 3191 20451
rect 4537 20417 4571 20451
rect 9873 20417 9907 20451
rect 11621 20417 11655 20451
rect 13001 20417 13035 20451
rect 16865 20417 16899 20451
rect 19073 20417 19107 20451
rect 21281 20417 21315 20451
rect 24133 20417 24167 20451
rect 24317 20417 24351 20451
rect 25421 20417 25455 20451
rect 1409 20349 1443 20383
rect 2421 20349 2455 20383
rect 2973 20349 3007 20383
rect 7665 20349 7699 20383
rect 9689 20349 9723 20383
rect 12265 20349 12299 20383
rect 12817 20349 12851 20383
rect 14105 20349 14139 20383
rect 14372 20349 14406 20383
rect 16681 20349 16715 20383
rect 17325 20349 17359 20383
rect 18981 20349 19015 20383
rect 19340 20349 19374 20383
rect 24041 20349 24075 20383
rect 24685 20349 24719 20383
rect 25237 20349 25271 20383
rect 25973 20349 26007 20383
rect 4782 20281 4816 20315
rect 7932 20281 7966 20315
rect 10118 20281 10152 20315
rect 12909 20281 12943 20315
rect 16773 20281 16807 20315
rect 17877 20281 17911 20315
rect 20821 20281 20855 20315
rect 21526 20281 21560 20315
rect 1593 20213 1627 20247
rect 2053 20213 2087 20247
rect 2881 20213 2915 20247
rect 3525 20213 3559 20247
rect 4353 20213 4387 20247
rect 9045 20213 9079 20247
rect 9413 20213 9447 20247
rect 12081 20213 12115 20247
rect 12449 20213 12483 20247
rect 13461 20213 13495 20247
rect 15853 20213 15887 20247
rect 18061 20213 18095 20247
rect 18521 20213 18555 20247
rect 20453 20213 20487 20247
rect 21097 20213 21131 20247
rect 22661 20213 22695 20247
rect 23029 20213 23063 20247
rect 23489 20213 23523 20247
rect 25053 20213 25087 20247
rect 1409 20009 1443 20043
rect 3525 20009 3559 20043
rect 3893 20009 3927 20043
rect 4353 20009 4387 20043
rect 6561 20009 6595 20043
rect 7389 20009 7423 20043
rect 8125 20009 8159 20043
rect 8493 20009 8527 20043
rect 10333 20009 10367 20043
rect 10793 20009 10827 20043
rect 11897 20009 11931 20043
rect 12357 20009 12391 20043
rect 12909 20009 12943 20043
rect 13461 20009 13495 20043
rect 14565 20009 14599 20043
rect 16681 20009 16715 20043
rect 17877 20009 17911 20043
rect 20913 20009 20947 20043
rect 22385 20009 22419 20043
rect 24317 20009 24351 20043
rect 24869 20009 24903 20043
rect 2329 19941 2363 19975
rect 4988 19941 5022 19975
rect 9505 19941 9539 19975
rect 13921 19941 13955 19975
rect 20269 19941 20303 19975
rect 22017 19941 22051 19975
rect 24685 19941 24719 19975
rect 2789 19873 2823 19907
rect 4721 19873 4755 19907
rect 7297 19873 7331 19907
rect 10149 19873 10183 19907
rect 10701 19873 10735 19907
rect 12265 19873 12299 19907
rect 13829 19873 13863 19907
rect 15301 19873 15335 19907
rect 15568 19873 15602 19907
rect 17969 19873 18003 19907
rect 19625 19873 19659 19907
rect 21281 19873 21315 19907
rect 21373 19873 21407 19907
rect 22661 19873 22695 19907
rect 22928 19873 22962 19907
rect 25237 19873 25271 19907
rect 2881 19805 2915 19839
rect 3065 19805 3099 19839
rect 7481 19805 7515 19839
rect 8585 19805 8619 19839
rect 10885 19805 10919 19839
rect 12541 19805 12575 19839
rect 13277 19805 13311 19839
rect 14013 19805 14047 19839
rect 18061 19805 18095 19839
rect 19717 19805 19751 19839
rect 19809 19805 19843 19839
rect 21465 19805 21499 19839
rect 25329 19805 25363 19839
rect 25513 19805 25547 19839
rect 2421 19737 2455 19771
rect 6101 19737 6135 19771
rect 6929 19737 6963 19771
rect 17049 19737 17083 19771
rect 17509 19737 17543 19771
rect 19165 19737 19199 19771
rect 24041 19737 24075 19771
rect 1869 19669 1903 19703
rect 9137 19669 9171 19703
rect 11437 19669 11471 19703
rect 11713 19669 11747 19703
rect 15025 19669 15059 19703
rect 17417 19669 17451 19703
rect 18521 19669 18555 19703
rect 19257 19669 19291 19703
rect 20729 19669 20763 19703
rect 2789 19465 2823 19499
rect 4445 19465 4479 19499
rect 6837 19465 6871 19499
rect 9689 19465 9723 19499
rect 11621 19465 11655 19499
rect 17601 19465 17635 19499
rect 19073 19465 19107 19499
rect 20545 19465 20579 19499
rect 20913 19465 20947 19499
rect 22845 19465 22879 19499
rect 2513 19397 2547 19431
rect 4077 19397 4111 19431
rect 11989 19397 12023 19431
rect 1961 19329 1995 19363
rect 3525 19329 3559 19363
rect 4537 19329 4571 19363
rect 7389 19329 7423 19363
rect 9137 19329 9171 19363
rect 10701 19329 10735 19363
rect 16957 19329 16991 19363
rect 21925 19329 21959 19363
rect 1777 19261 1811 19295
rect 3341 19261 3375 19295
rect 8125 19261 8159 19295
rect 9965 19261 9999 19295
rect 10609 19261 10643 19295
rect 12449 19261 12483 19295
rect 13369 19261 13403 19295
rect 13553 19261 13587 19295
rect 15393 19261 15427 19295
rect 16037 19261 16071 19295
rect 16773 19261 16807 19295
rect 18061 19261 18095 19295
rect 19165 19261 19199 19295
rect 21741 19261 21775 19295
rect 23673 19261 23707 19295
rect 3433 19193 3467 19227
rect 4804 19193 4838 19227
rect 6285 19193 6319 19227
rect 8493 19193 8527 19227
rect 10517 19193 10551 19227
rect 13820 19193 13854 19227
rect 15761 19193 15795 19227
rect 18613 19193 18647 19227
rect 19432 19193 19466 19227
rect 21833 19193 21867 19227
rect 23918 19193 23952 19227
rect 25421 19193 25455 19227
rect 1409 19125 1443 19159
rect 1869 19125 1903 19159
rect 2973 19125 3007 19159
rect 5917 19125 5951 19159
rect 6653 19125 6687 19159
rect 7205 19125 7239 19159
rect 7297 19125 7331 19159
rect 8585 19125 8619 19159
rect 8953 19125 8987 19159
rect 9045 19125 9079 19159
rect 10149 19125 10183 19159
rect 11253 19125 11287 19159
rect 12633 19125 12667 19159
rect 13093 19125 13127 19159
rect 14933 19125 14967 19159
rect 15853 19125 15887 19159
rect 16405 19125 16439 19159
rect 16865 19125 16899 19159
rect 18245 19125 18279 19159
rect 21189 19125 21223 19159
rect 21373 19125 21407 19159
rect 22385 19125 22419 19159
rect 23489 19125 23523 19159
rect 25053 19125 25087 19159
rect 25697 19125 25731 19159
rect 2329 18921 2363 18955
rect 3065 18921 3099 18955
rect 4905 18921 4939 18955
rect 6009 18921 6043 18955
rect 7481 18921 7515 18955
rect 7849 18921 7883 18955
rect 9505 18921 9539 18955
rect 11989 18921 12023 18955
rect 12357 18921 12391 18955
rect 13829 18921 13863 18955
rect 18889 18921 18923 18955
rect 19257 18921 19291 18955
rect 19993 18921 20027 18955
rect 20729 18921 20763 18955
rect 21281 18921 21315 18955
rect 21925 18921 21959 18955
rect 23397 18921 23431 18955
rect 24869 18921 24903 18955
rect 25329 18921 25363 18955
rect 4629 18853 4663 18887
rect 6285 18853 6319 18887
rect 9956 18853 9990 18887
rect 15669 18853 15703 18887
rect 18337 18853 18371 18887
rect 18705 18853 18739 18887
rect 19349 18853 19383 18887
rect 24961 18853 24995 18887
rect 5273 18785 5307 18819
rect 6837 18785 6871 18819
rect 8401 18785 8435 18819
rect 9689 18785 9723 18819
rect 12449 18785 12483 18819
rect 12716 18785 12750 18819
rect 14473 18785 14507 18819
rect 15117 18785 15151 18819
rect 15393 18785 15427 18819
rect 16497 18785 16531 18819
rect 16948 18785 16982 18819
rect 23305 18785 23339 18819
rect 24317 18785 24351 18819
rect 2421 18717 2455 18751
rect 2513 18717 2547 18751
rect 3893 18717 3927 18751
rect 5365 18717 5399 18751
rect 5549 18717 5583 18751
rect 6929 18717 6963 18751
rect 7021 18717 7055 18751
rect 8493 18717 8527 18751
rect 8585 18717 8619 18751
rect 16681 18717 16715 18751
rect 19441 18717 19475 18751
rect 21373 18717 21407 18751
rect 21465 18717 21499 18751
rect 23489 18717 23523 18751
rect 25053 18717 25087 18751
rect 25605 18853 25639 18887
rect 25881 18785 25915 18819
rect 9045 18649 9079 18683
rect 20913 18649 20947 18683
rect 22293 18649 22327 18683
rect 22845 18649 22879 18683
rect 24501 18649 24535 18683
rect 25329 18649 25363 18683
rect 1869 18581 1903 18615
rect 1961 18581 1995 18615
rect 3433 18581 3467 18615
rect 6469 18581 6503 18615
rect 8033 18581 8067 18615
rect 11069 18581 11103 18615
rect 11437 18581 11471 18615
rect 14105 18581 14139 18615
rect 18061 18581 18095 18615
rect 20361 18581 20395 18615
rect 22937 18581 22971 18615
rect 23949 18581 23983 18615
rect 1593 18377 1627 18411
rect 6561 18377 6595 18411
rect 10517 18377 10551 18411
rect 11897 18377 11931 18411
rect 12817 18377 12851 18411
rect 13829 18377 13863 18411
rect 14381 18377 14415 18411
rect 15485 18377 15519 18411
rect 16313 18377 16347 18411
rect 19533 18377 19567 18411
rect 21833 18377 21867 18411
rect 23305 18377 23339 18411
rect 25053 18377 25087 18411
rect 25789 18377 25823 18411
rect 5733 18309 5767 18343
rect 9689 18309 9723 18343
rect 9965 18309 9999 18343
rect 10241 18309 10275 18343
rect 16405 18309 16439 18343
rect 21281 18309 21315 18343
rect 21649 18309 21683 18343
rect 4353 18241 4387 18275
rect 11069 18241 11103 18275
rect 12265 18241 12299 18275
rect 13461 18241 13495 18275
rect 14933 18241 14967 18275
rect 17049 18241 17083 18275
rect 17877 18241 17911 18275
rect 18613 18241 18647 18275
rect 19625 18241 19659 18275
rect 22385 18241 22419 18275
rect 25329 18241 25363 18275
rect 2145 18173 2179 18207
rect 6101 18173 6135 18207
rect 6837 18173 6871 18207
rect 8309 18173 8343 18207
rect 10241 18173 10275 18207
rect 10977 18173 11011 18207
rect 14749 18173 14783 18207
rect 18429 18173 18463 18207
rect 18521 18173 18555 18207
rect 19165 18173 19199 18207
rect 22293 18173 22327 18207
rect 23673 18173 23707 18207
rect 2412 18105 2446 18139
rect 4169 18105 4203 18139
rect 4598 18105 4632 18139
rect 7113 18105 7147 18139
rect 8217 18105 8251 18139
rect 8554 18105 8588 18139
rect 10425 18105 10459 18139
rect 10885 18105 10919 18139
rect 13277 18105 13311 18139
rect 15945 18105 15979 18139
rect 16773 18105 16807 18139
rect 19892 18105 19926 18139
rect 22201 18105 22235 18139
rect 23918 18105 23952 18139
rect 26065 18105 26099 18139
rect 2053 18037 2087 18071
rect 3525 18037 3559 18071
rect 3801 18037 3835 18071
rect 7757 18037 7791 18071
rect 12633 18037 12667 18071
rect 13185 18037 13219 18071
rect 14197 18037 14231 18071
rect 14841 18037 14875 18071
rect 16865 18037 16899 18071
rect 17509 18037 17543 18071
rect 18061 18037 18095 18071
rect 21005 18037 21039 18071
rect 23029 18037 23063 18071
rect 3157 17833 3191 17867
rect 4261 17833 4295 17867
rect 4905 17833 4939 17867
rect 5273 17833 5307 17867
rect 6929 17833 6963 17867
rect 9045 17833 9079 17867
rect 9413 17833 9447 17867
rect 10609 17833 10643 17867
rect 13185 17833 13219 17867
rect 14381 17833 14415 17867
rect 15577 17833 15611 17867
rect 17877 17833 17911 17867
rect 18153 17833 18187 17867
rect 18705 17833 18739 17867
rect 20085 17833 20119 17867
rect 20637 17833 20671 17867
rect 20913 17833 20947 17867
rect 21373 17833 21407 17867
rect 22293 17833 22327 17867
rect 25053 17833 25087 17867
rect 25789 17833 25823 17867
rect 10149 17765 10183 17799
rect 13829 17765 13863 17799
rect 19073 17765 19107 17799
rect 21925 17765 21959 17799
rect 22845 17765 22879 17799
rect 25421 17765 25455 17799
rect 1777 17697 1811 17731
rect 2044 17697 2078 17731
rect 3893 17697 3927 17731
rect 4077 17697 4111 17731
rect 5641 17697 5675 17731
rect 7205 17697 7239 17731
rect 7389 17697 7423 17731
rect 7656 17697 7690 17731
rect 9873 17697 9907 17731
rect 11428 17697 11462 17731
rect 13737 17697 13771 17731
rect 15393 17697 15427 17731
rect 16313 17697 16347 17731
rect 16764 17697 16798 17731
rect 21281 17697 21315 17731
rect 24409 17697 24443 17731
rect 24501 17697 24535 17731
rect 5733 17629 5767 17663
rect 5917 17629 5951 17663
rect 11161 17629 11195 17663
rect 13921 17629 13955 17663
rect 16497 17629 16531 17663
rect 19165 17629 19199 17663
rect 19257 17629 19291 17663
rect 19717 17629 19751 17663
rect 21465 17629 21499 17663
rect 22937 17629 22971 17663
rect 23029 17629 23063 17663
rect 24685 17629 24719 17663
rect 8769 17561 8803 17595
rect 12817 17561 12851 17595
rect 13369 17561 13403 17595
rect 22477 17561 22511 17595
rect 1685 17493 1719 17527
rect 3433 17493 3467 17527
rect 6469 17493 6503 17527
rect 11069 17493 11103 17527
rect 12541 17493 12575 17527
rect 14841 17493 14875 17527
rect 18613 17493 18647 17527
rect 23765 17493 23799 17527
rect 24041 17493 24075 17527
rect 3617 17289 3651 17323
rect 5917 17289 5951 17323
rect 6653 17289 6687 17323
rect 7573 17289 7607 17323
rect 11621 17289 11655 17323
rect 14105 17289 14139 17323
rect 14565 17289 14599 17323
rect 17785 17289 17819 17323
rect 18337 17289 18371 17323
rect 18797 17289 18831 17323
rect 23489 17289 23523 17323
rect 23673 17289 23707 17323
rect 2973 17221 3007 17255
rect 4445 17221 4479 17255
rect 11345 17221 11379 17255
rect 14657 17221 14691 17255
rect 15669 17221 15703 17255
rect 17325 17221 17359 17255
rect 23029 17221 23063 17255
rect 1777 17153 1811 17187
rect 2513 17153 2547 17187
rect 4537 17153 4571 17187
rect 7021 17153 7055 17187
rect 7941 17153 7975 17187
rect 10149 17153 10183 17187
rect 10701 17153 10735 17187
rect 10885 17153 10919 17187
rect 15117 17153 15151 17187
rect 15209 17153 15243 17187
rect 16129 17153 16163 17187
rect 16773 17153 16807 17187
rect 24133 17153 24167 17187
rect 24225 17153 24259 17187
rect 25053 17153 25087 17187
rect 3433 17085 3467 17119
rect 8033 17085 8067 17119
rect 8300 17085 8334 17119
rect 12449 17085 12483 17119
rect 16589 17085 16623 17119
rect 18981 17085 19015 17119
rect 19237 17085 19271 17119
rect 21189 17085 21223 17119
rect 25237 17085 25271 17119
rect 25973 17085 26007 17119
rect 2329 17017 2363 17051
rect 3341 17017 3375 17051
rect 4804 17017 4838 17051
rect 9781 17017 9815 17051
rect 10609 17017 10643 17051
rect 12716 17017 12750 17051
rect 15025 17017 15059 17051
rect 16681 17017 16715 17051
rect 21005 17017 21039 17051
rect 21456 17017 21490 17051
rect 25513 17017 25547 17051
rect 1869 16949 1903 16983
rect 2237 16949 2271 16983
rect 4077 16949 4111 16983
rect 6285 16949 6319 16983
rect 9413 16949 9447 16983
rect 10241 16949 10275 16983
rect 12173 16949 12207 16983
rect 13829 16949 13863 16983
rect 16221 16949 16255 16983
rect 20361 16949 20395 16983
rect 22569 16949 22603 16983
rect 24041 16949 24075 16983
rect 24685 16949 24719 16983
rect 26341 16949 26375 16983
rect 1777 16745 1811 16779
rect 3617 16745 3651 16779
rect 4261 16745 4295 16779
rect 5181 16745 5215 16779
rect 5641 16745 5675 16779
rect 6929 16745 6963 16779
rect 8861 16745 8895 16779
rect 10701 16745 10735 16779
rect 12909 16745 12943 16779
rect 14657 16745 14691 16779
rect 15025 16745 15059 16779
rect 17693 16745 17727 16779
rect 18613 16745 18647 16779
rect 18797 16745 18831 16779
rect 19165 16745 19199 16779
rect 20269 16745 20303 16779
rect 20545 16745 20579 16779
rect 20913 16745 20947 16779
rect 21373 16745 21407 16779
rect 21925 16745 21959 16779
rect 22569 16745 22603 16779
rect 24133 16745 24167 16779
rect 24869 16745 24903 16779
rect 25145 16745 25179 16779
rect 2145 16677 2179 16711
rect 2881 16677 2915 16711
rect 3341 16677 3375 16711
rect 7665 16677 7699 16711
rect 9229 16677 9263 16711
rect 17601 16677 17635 16711
rect 19625 16677 19659 16711
rect 4077 16609 4111 16643
rect 5549 16609 5583 16643
rect 6561 16609 6595 16643
rect 6745 16609 6779 16643
rect 7297 16609 7331 16643
rect 8217 16609 8251 16643
rect 9873 16609 9907 16643
rect 10149 16609 10183 16643
rect 11161 16609 11195 16643
rect 11428 16609 11462 16643
rect 13185 16609 13219 16643
rect 13737 16609 13771 16643
rect 15485 16609 15519 16643
rect 15752 16609 15786 16643
rect 18061 16609 18095 16643
rect 18153 16609 18187 16643
rect 18613 16609 18647 16643
rect 25513 16677 25547 16711
rect 21281 16609 21315 16643
rect 22753 16609 22787 16643
rect 23020 16609 23054 16643
rect 24961 16609 24995 16643
rect 2237 16541 2271 16575
rect 2421 16541 2455 16575
rect 5825 16541 5859 16575
rect 8309 16541 8343 16575
rect 8493 16541 8527 16575
rect 13829 16541 13863 16575
rect 13921 16541 13955 16575
rect 18337 16541 18371 16575
rect 19717 16541 19751 16575
rect 19809 16541 19843 16575
rect 20545 16541 20579 16575
rect 21465 16541 21499 16575
rect 16865 16473 16899 16507
rect 19257 16473 19291 16507
rect 1685 16405 1719 16439
rect 4721 16405 4755 16439
rect 5089 16405 5123 16439
rect 6285 16405 6319 16439
rect 7849 16405 7883 16439
rect 11069 16405 11103 16439
rect 12541 16405 12575 16439
rect 13369 16405 13403 16439
rect 17233 16405 17267 16439
rect 20637 16405 20671 16439
rect 24501 16405 24535 16439
rect 2237 16201 2271 16235
rect 2697 16201 2731 16235
rect 4445 16201 4479 16235
rect 5089 16201 5123 16235
rect 6561 16201 6595 16235
rect 7849 16201 7883 16235
rect 9321 16201 9355 16235
rect 9689 16201 9723 16235
rect 10333 16201 10367 16235
rect 13553 16201 13587 16235
rect 14013 16201 14047 16235
rect 17049 16201 17083 16235
rect 20453 16201 20487 16235
rect 21465 16201 21499 16235
rect 22017 16201 22051 16235
rect 23673 16201 23707 16235
rect 24961 16201 24995 16235
rect 25421 16201 25455 16235
rect 26157 16201 26191 16235
rect 2881 16133 2915 16167
rect 6193 16133 6227 16167
rect 10701 16133 10735 16167
rect 19993 16133 20027 16167
rect 21925 16133 21959 16167
rect 3433 16065 3467 16099
rect 5825 16065 5859 16099
rect 11253 16065 11287 16099
rect 11345 16065 11379 16099
rect 11897 16065 11931 16099
rect 13001 16065 13035 16099
rect 14565 16065 14599 16099
rect 15025 16065 15059 16099
rect 15485 16065 15519 16099
rect 16221 16065 16255 16099
rect 21097 16065 21131 16099
rect 22569 16065 22603 16099
rect 24225 16065 24259 16099
rect 1409 15997 1443 16031
rect 3341 15997 3375 16031
rect 4629 15997 4663 16031
rect 5641 15997 5675 16031
rect 7941 15997 7975 16031
rect 14473 15997 14507 16031
rect 18061 15997 18095 16031
rect 23121 15997 23155 16031
rect 25237 15997 25271 16031
rect 25789 15997 25823 16031
rect 1685 15929 1719 15963
rect 7481 15929 7515 15963
rect 8208 15929 8242 15963
rect 12265 15929 12299 15963
rect 12817 15929 12851 15963
rect 13921 15929 13955 15963
rect 14381 15929 14415 15963
rect 17325 15929 17359 15963
rect 18306 15929 18340 15963
rect 20361 15929 20395 15963
rect 20821 15929 20855 15963
rect 24133 15929 24167 15963
rect 3249 15861 3283 15895
rect 4169 15861 4203 15895
rect 5181 15861 5215 15895
rect 5549 15861 5583 15895
rect 6837 15861 6871 15895
rect 10793 15861 10827 15895
rect 11161 15861 11195 15895
rect 12449 15861 12483 15895
rect 12909 15861 12943 15895
rect 15577 15861 15611 15895
rect 15945 15861 15979 15895
rect 16037 15861 16071 15895
rect 16681 15861 16715 15895
rect 17785 15861 17819 15895
rect 19441 15861 19475 15895
rect 20913 15861 20947 15895
rect 22385 15861 22419 15895
rect 22477 15861 22511 15895
rect 23489 15861 23523 15895
rect 24041 15861 24075 15895
rect 1961 15657 1995 15691
rect 3341 15657 3375 15691
rect 8033 15657 8067 15691
rect 8401 15657 8435 15691
rect 13001 15657 13035 15691
rect 13461 15657 13495 15691
rect 14381 15657 14415 15691
rect 16681 15657 16715 15691
rect 17417 15657 17451 15691
rect 17693 15657 17727 15691
rect 18153 15657 18187 15691
rect 18521 15657 18555 15691
rect 19993 15657 20027 15691
rect 22109 15657 22143 15691
rect 23857 15657 23891 15691
rect 24133 15657 24167 15691
rect 24501 15657 24535 15691
rect 25145 15657 25179 15691
rect 2421 15589 2455 15623
rect 7941 15589 7975 15623
rect 10701 15589 10735 15623
rect 13369 15589 13403 15623
rect 14749 15589 14783 15623
rect 21281 15589 21315 15623
rect 22722 15589 22756 15623
rect 2329 15521 2363 15555
rect 4077 15521 4111 15555
rect 4333 15521 4367 15555
rect 6653 15521 6687 15555
rect 8493 15521 8527 15555
rect 11060 15521 11094 15555
rect 12909 15521 12943 15555
rect 14105 15521 14139 15555
rect 15568 15521 15602 15555
rect 17509 15521 17543 15555
rect 18880 15521 18914 15555
rect 21373 15521 21407 15555
rect 22477 15521 22511 15555
rect 25053 15521 25087 15555
rect 2513 15453 2547 15487
rect 3893 15453 3927 15487
rect 6745 15453 6779 15487
rect 6929 15453 6963 15487
rect 8677 15453 8711 15487
rect 9781 15453 9815 15487
rect 10333 15453 10367 15487
rect 10793 15453 10827 15487
rect 13645 15453 13679 15487
rect 15301 15453 15335 15487
rect 18613 15453 18647 15487
rect 21465 15453 21499 15487
rect 25329 15453 25363 15487
rect 6285 15385 6319 15419
rect 24685 15385 24719 15419
rect 1685 15317 1719 15351
rect 3065 15317 3099 15351
rect 5457 15317 5491 15351
rect 5825 15317 5859 15351
rect 6101 15317 6135 15351
rect 7389 15317 7423 15351
rect 9137 15317 9171 15351
rect 9505 15317 9539 15351
rect 12173 15317 12207 15351
rect 12541 15317 12575 15351
rect 16957 15317 16991 15351
rect 20545 15317 20579 15351
rect 20913 15317 20947 15351
rect 2513 15113 2547 15147
rect 2697 15113 2731 15147
rect 5181 15113 5215 15147
rect 6561 15113 6595 15147
rect 6837 15113 6871 15147
rect 7021 15113 7055 15147
rect 8493 15113 8527 15147
rect 9137 15113 9171 15147
rect 11161 15113 11195 15147
rect 11437 15113 11471 15147
rect 12173 15113 12207 15147
rect 12449 15113 12483 15147
rect 13553 15113 13587 15147
rect 13829 15113 13863 15147
rect 17049 15113 17083 15147
rect 17877 15113 17911 15147
rect 19533 15113 19567 15147
rect 20269 15113 20303 15147
rect 22661 15113 22695 15147
rect 23673 15113 23707 15147
rect 24777 15113 24811 15147
rect 24961 15113 24995 15147
rect 25053 15113 25087 15147
rect 2237 15045 2271 15079
rect 1409 14909 1443 14943
rect 1685 14841 1719 14875
rect 2789 14977 2823 15011
rect 5089 14977 5123 15011
rect 5733 14977 5767 15011
rect 3056 14909 3090 14943
rect 5549 14909 5583 14943
rect 6285 14909 6319 14943
rect 8125 15045 8159 15079
rect 25421 15045 25455 15079
rect 7665 14977 7699 15011
rect 8585 14977 8619 15011
rect 11897 14977 11931 15011
rect 13093 14977 13127 15011
rect 19901 14977 19935 15011
rect 20821 14977 20855 15011
rect 20913 14977 20947 15011
rect 23121 14977 23155 15011
rect 24225 14977 24259 15011
rect 24961 14977 24995 15011
rect 9781 14909 9815 14943
rect 12909 14909 12943 14943
rect 14657 14909 14691 14943
rect 16865 14909 16899 14943
rect 18153 14909 18187 14943
rect 21373 14909 21407 14943
rect 21925 14909 21959 14943
rect 24041 14909 24075 14943
rect 25237 14909 25271 14943
rect 25789 14909 25823 14943
rect 6837 14841 6871 14875
rect 7389 14841 7423 14875
rect 9689 14841 9723 14875
rect 10048 14841 10082 14875
rect 14565 14841 14599 14875
rect 14902 14841 14936 14875
rect 17509 14841 17543 14875
rect 18420 14841 18454 14875
rect 20729 14841 20763 14875
rect 21741 14841 21775 14875
rect 22201 14841 22235 14875
rect 23489 14841 23523 14875
rect 24133 14841 24167 14875
rect 2697 14773 2731 14807
rect 4169 14773 4203 14807
rect 4445 14773 4479 14807
rect 5641 14773 5675 14807
rect 7481 14773 7515 14807
rect 12817 14773 12851 14807
rect 16037 14773 16071 14807
rect 16313 14773 16347 14807
rect 16681 14773 16715 14807
rect 20361 14773 20395 14807
rect 1961 14569 1995 14603
rect 2421 14569 2455 14603
rect 2881 14569 2915 14603
rect 3249 14569 3283 14603
rect 3893 14569 3927 14603
rect 4261 14569 4295 14603
rect 5733 14569 5767 14603
rect 8033 14569 8067 14603
rect 8401 14569 8435 14603
rect 9045 14569 9079 14603
rect 9505 14569 9539 14603
rect 10609 14569 10643 14603
rect 10977 14569 11011 14603
rect 12725 14569 12759 14603
rect 13277 14569 13311 14603
rect 15117 14569 15151 14603
rect 16221 14569 16255 14603
rect 16681 14569 16715 14603
rect 17509 14569 17543 14603
rect 19257 14569 19291 14603
rect 20453 14569 20487 14603
rect 21097 14569 21131 14603
rect 21557 14569 21591 14603
rect 22017 14569 22051 14603
rect 22385 14569 22419 14603
rect 22661 14569 22695 14603
rect 24041 14569 24075 14603
rect 25053 14569 25087 14603
rect 2789 14433 2823 14467
rect 1409 14365 1443 14399
rect 2329 14365 2363 14399
rect 3065 14365 3099 14399
rect 4629 14501 4663 14535
rect 5365 14501 5399 14535
rect 6092 14501 6126 14535
rect 11336 14501 11370 14535
rect 13645 14501 13679 14535
rect 13737 14501 13771 14535
rect 16773 14501 16807 14535
rect 18144 14501 18178 14535
rect 19717 14501 19751 14535
rect 4721 14433 4755 14467
rect 5825 14433 5859 14467
rect 8493 14433 8527 14467
rect 9781 14433 9815 14467
rect 10057 14433 10091 14467
rect 11069 14433 11103 14467
rect 20729 14433 20763 14467
rect 20913 14433 20947 14467
rect 23029 14433 23063 14467
rect 24225 14433 24259 14467
rect 4905 14365 4939 14399
rect 7481 14365 7515 14399
rect 8677 14365 8711 14399
rect 13185 14365 13219 14399
rect 13829 14365 13863 14399
rect 15301 14365 15335 14399
rect 16957 14365 16991 14399
rect 17877 14365 17911 14399
rect 19993 14365 20027 14399
rect 23121 14365 23155 14399
rect 23213 14365 23247 14399
rect 24501 14365 24535 14399
rect 3433 14297 3467 14331
rect 7941 14297 7975 14331
rect 16313 14297 16347 14331
rect 3249 14229 3283 14263
rect 7205 14229 7239 14263
rect 12449 14229 12483 14263
rect 14289 14229 14323 14263
rect 14657 14229 14691 14263
rect 15853 14229 15887 14263
rect 20545 14229 20579 14263
rect 23673 14229 23707 14263
rect 2513 14025 2547 14059
rect 4261 14025 4295 14059
rect 4629 14025 4663 14059
rect 4905 14025 4939 14059
rect 5181 14025 5215 14059
rect 6285 14025 6319 14059
rect 6561 14025 6595 14059
rect 8861 14025 8895 14059
rect 10425 14025 10459 14059
rect 15761 14025 15795 14059
rect 16405 14025 16439 14059
rect 17509 14025 17543 14059
rect 17877 14025 17911 14059
rect 19165 14025 19199 14059
rect 21005 14025 21039 14059
rect 21833 14025 21867 14059
rect 22109 14025 22143 14059
rect 23121 14025 23155 14059
rect 23489 14025 23523 14059
rect 12449 13957 12483 13991
rect 18061 13957 18095 13991
rect 21465 13957 21499 13991
rect 1685 13889 1719 13923
rect 5825 13889 5859 13923
rect 8493 13889 8527 13923
rect 10793 13889 10827 13923
rect 12173 13889 12207 13923
rect 13001 13889 13035 13923
rect 14013 13889 14047 13923
rect 16957 13889 16991 13923
rect 18521 13889 18555 13923
rect 18613 13889 18647 13923
rect 20177 13889 20211 13923
rect 1409 13821 1443 13855
rect 2881 13821 2915 13855
rect 6837 13821 6871 13855
rect 7093 13821 7127 13855
rect 9045 13821 9079 13855
rect 11897 13821 11931 13855
rect 12909 13821 12943 13855
rect 14381 13821 14415 13855
rect 14648 13821 14682 13855
rect 16681 13821 16715 13855
rect 19533 13821 19567 13855
rect 20085 13821 20119 13855
rect 21925 13821 21959 13855
rect 22753 13821 22787 13855
rect 23673 13821 23707 13855
rect 23929 13821 23963 13855
rect 3148 13753 3182 13787
rect 5549 13753 5583 13787
rect 9290 13753 9324 13787
rect 11253 13753 11287 13787
rect 13921 13753 13955 13787
rect 19993 13753 20027 13787
rect 5641 13685 5675 13719
rect 8217 13685 8251 13719
rect 11161 13685 11195 13719
rect 12817 13685 12851 13719
rect 13461 13685 13495 13719
rect 13829 13685 13863 13719
rect 18429 13685 18463 13719
rect 19625 13685 19659 13719
rect 25053 13685 25087 13719
rect 2421 13481 2455 13515
rect 2881 13481 2915 13515
rect 4445 13481 4479 13515
rect 5181 13481 5215 13515
rect 5641 13481 5675 13515
rect 7113 13481 7147 13515
rect 9137 13481 9171 13515
rect 9505 13481 9539 13515
rect 10057 13481 10091 13515
rect 11897 13481 11931 13515
rect 12633 13481 12667 13515
rect 15301 13481 15335 13515
rect 16405 13481 16439 13515
rect 16773 13481 16807 13515
rect 16865 13481 16899 13515
rect 17417 13481 17451 13515
rect 17785 13481 17819 13515
rect 18245 13481 18279 13515
rect 18613 13481 18647 13515
rect 19809 13481 19843 13515
rect 21649 13481 21683 13515
rect 22753 13481 22787 13515
rect 23673 13481 23707 13515
rect 24869 13481 24903 13515
rect 25513 13481 25547 13515
rect 2329 13413 2363 13447
rect 3893 13413 3927 13447
rect 4537 13413 4571 13447
rect 8309 13413 8343 13447
rect 15669 13413 15703 13447
rect 2789 13345 2823 13379
rect 5733 13345 5767 13379
rect 6000 13345 6034 13379
rect 10773 13345 10807 13379
rect 12725 13345 12759 13379
rect 18061 13345 18095 13379
rect 20545 13345 20579 13379
rect 21465 13345 21499 13379
rect 22569 13345 22603 13379
rect 24041 13345 24075 13379
rect 25329 13345 25363 13379
rect 2973 13277 3007 13311
rect 4721 13277 4755 13311
rect 8401 13277 8435 13311
rect 8493 13277 8527 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 10517 13277 10551 13311
rect 15761 13277 15795 13311
rect 15853 13277 15887 13311
rect 18705 13277 18739 13311
rect 18889 13277 18923 13311
rect 24225 13277 24259 13311
rect 4077 13209 4111 13243
rect 7481 13209 7515 13243
rect 7849 13209 7883 13243
rect 14013 13209 14047 13243
rect 17877 13209 17911 13243
rect 19257 13209 19291 13243
rect 1961 13141 1995 13175
rect 3525 13141 3559 13175
rect 7941 13141 7975 13175
rect 9689 13141 9723 13175
rect 12265 13141 12299 13175
rect 15025 13141 15059 13175
rect 19625 13141 19659 13175
rect 1593 12937 1627 12971
rect 4261 12937 4295 12971
rect 5825 12937 5859 12971
rect 6837 12937 6871 12971
rect 8033 12937 8067 12971
rect 9321 12937 9355 12971
rect 10333 12937 10367 12971
rect 14749 12937 14783 12971
rect 15025 12937 15059 12971
rect 15209 12937 15243 12971
rect 17509 12937 17543 12971
rect 18889 12937 18923 12971
rect 19901 12937 19935 12971
rect 21281 12937 21315 12971
rect 22661 12937 22695 12971
rect 23029 12937 23063 12971
rect 2513 12869 2547 12903
rect 5273 12869 5307 12903
rect 9597 12869 9631 12903
rect 17877 12869 17911 12903
rect 21557 12869 21591 12903
rect 22385 12869 22419 12903
rect 2145 12801 2179 12835
rect 3249 12801 3283 12835
rect 3801 12801 3835 12835
rect 4169 12801 4203 12835
rect 4721 12801 4755 12835
rect 4813 12801 4847 12835
rect 6285 12801 6319 12835
rect 7481 12801 7515 12835
rect 8677 12801 8711 12835
rect 11345 12801 11379 12835
rect 11805 12801 11839 12835
rect 13001 12801 13035 12835
rect 15761 12801 15795 12835
rect 16773 12801 16807 12835
rect 19441 12801 19475 12835
rect 23489 12801 23523 12835
rect 1409 12733 1443 12767
rect 4629 12733 4663 12767
rect 7297 12733 7331 12767
rect 8585 12733 8619 12767
rect 10701 12733 10735 12767
rect 13268 12733 13302 12767
rect 21373 12733 21407 12767
rect 21925 12733 21959 12767
rect 22477 12733 22511 12767
rect 23673 12733 23707 12767
rect 23940 12733 23974 12767
rect 3065 12665 3099 12699
rect 6653 12665 6687 12699
rect 7205 12665 7239 12699
rect 9781 12665 9815 12699
rect 11161 12665 11195 12699
rect 12265 12665 12299 12699
rect 15577 12665 15611 12699
rect 16589 12665 16623 12699
rect 18429 12665 18463 12699
rect 19257 12665 19291 12699
rect 2697 12597 2731 12631
rect 3157 12597 3191 12631
rect 8401 12597 8435 12631
rect 10793 12597 10827 12631
rect 11253 12597 11287 12631
rect 12725 12597 12759 12631
rect 14381 12597 14415 12631
rect 15669 12597 15703 12631
rect 16221 12597 16255 12631
rect 18705 12597 18739 12631
rect 19349 12597 19383 12631
rect 25053 12597 25087 12631
rect 25329 12597 25363 12631
rect 1593 12393 1627 12427
rect 2421 12393 2455 12427
rect 4077 12393 4111 12427
rect 4537 12393 4571 12427
rect 5181 12393 5215 12427
rect 6285 12393 6319 12427
rect 6929 12393 6963 12427
rect 8033 12393 8067 12427
rect 8401 12393 8435 12427
rect 8677 12393 8711 12427
rect 10425 12393 10459 12427
rect 11437 12393 11471 12427
rect 13001 12393 13035 12427
rect 14657 12393 14691 12427
rect 15025 12393 15059 12427
rect 15301 12393 15335 12427
rect 16681 12393 16715 12427
rect 17969 12393 18003 12427
rect 18337 12393 18371 12427
rect 19533 12393 19567 12427
rect 21833 12393 21867 12427
rect 22937 12393 22971 12427
rect 2789 12325 2823 12359
rect 3525 12325 3559 12359
rect 9965 12325 9999 12359
rect 11897 12325 11931 12359
rect 18613 12325 18647 12359
rect 23673 12325 23707 12359
rect 2881 12257 2915 12291
rect 4445 12257 4479 12291
rect 11805 12257 11839 12291
rect 13369 12257 13403 12291
rect 13461 12257 13495 12291
rect 15669 12257 15703 12291
rect 17233 12257 17267 12291
rect 19165 12257 19199 12291
rect 21649 12257 21683 12291
rect 22753 12257 22787 12291
rect 24225 12257 24259 12291
rect 25421 12257 25455 12291
rect 3065 12189 3099 12223
rect 4721 12189 4755 12223
rect 5549 12189 5583 12223
rect 5825 12189 5859 12223
rect 11253 12189 11287 12223
rect 11989 12189 12023 12223
rect 13553 12189 13587 12223
rect 15761 12189 15795 12223
rect 15853 12189 15887 12223
rect 16313 12189 16347 12223
rect 17325 12189 17359 12223
rect 17417 12189 17451 12223
rect 19809 12189 19843 12223
rect 24317 12189 24351 12223
rect 24501 12189 24535 12223
rect 2329 12121 2363 12155
rect 3893 12121 3927 12155
rect 10885 12121 10919 12155
rect 23857 12121 23891 12155
rect 24869 12121 24903 12155
rect 12817 12053 12851 12087
rect 14105 12053 14139 12087
rect 16865 12053 16899 12087
rect 1593 11849 1627 11883
rect 2053 11849 2087 11883
rect 2421 11849 2455 11883
rect 3065 11849 3099 11883
rect 4445 11849 4479 11883
rect 4813 11849 4847 11883
rect 11161 11849 11195 11883
rect 11529 11849 11563 11883
rect 12725 11849 12759 11883
rect 14565 11849 14599 11883
rect 16129 11849 16163 11883
rect 17233 11849 17267 11883
rect 17509 11849 17543 11883
rect 18245 11849 18279 11883
rect 18613 11849 18647 11883
rect 21925 11849 21959 11883
rect 22661 11849 22695 11883
rect 23029 11849 23063 11883
rect 23489 11849 23523 11883
rect 25053 11849 25087 11883
rect 4169 11781 4203 11815
rect 12173 11781 12207 11815
rect 3617 11713 3651 11747
rect 11805 11713 11839 11747
rect 13277 11713 13311 11747
rect 15117 11713 15151 11747
rect 16589 11713 16623 11747
rect 16681 11713 16715 11747
rect 21465 11713 21499 11747
rect 22293 11713 22327 11747
rect 24685 11713 24719 11747
rect 25605 11713 25639 11747
rect 1409 11645 1443 11679
rect 3433 11645 3467 11679
rect 13737 11645 13771 11679
rect 22477 11645 22511 11679
rect 24409 11645 24443 11679
rect 15025 11577 15059 11611
rect 15669 11577 15703 11611
rect 25421 11577 25455 11611
rect 2973 11509 3007 11543
rect 3525 11509 3559 11543
rect 13093 11509 13127 11543
rect 13185 11509 13219 11543
rect 14381 11509 14415 11543
rect 14933 11509 14967 11543
rect 16037 11509 16071 11543
rect 16497 11509 16531 11543
rect 23857 11509 23891 11543
rect 24041 11509 24075 11543
rect 24501 11509 24535 11543
rect 1685 11305 1719 11339
rect 2145 11305 2179 11339
rect 3157 11305 3191 11339
rect 3525 11305 3559 11339
rect 11437 11305 11471 11339
rect 12357 11305 12391 11339
rect 13001 11305 13035 11339
rect 15301 11305 15335 11339
rect 16405 11305 16439 11339
rect 17233 11305 17267 11339
rect 22569 11305 22603 11339
rect 23673 11305 23707 11339
rect 24501 11305 24535 11339
rect 2513 11237 2547 11271
rect 12817 11237 12851 11271
rect 13369 11237 13403 11271
rect 15117 11237 15151 11271
rect 15761 11237 15795 11271
rect 14657 11169 14691 11203
rect 15669 11169 15703 11203
rect 22385 11169 22419 11203
rect 23489 11169 23523 11203
rect 24593 11169 24627 11203
rect 13461 11101 13495 11135
rect 13645 11101 13679 11135
rect 15945 11101 15979 11135
rect 24133 11101 24167 11135
rect 14289 11033 14323 11067
rect 16865 11033 16899 11067
rect 24777 11033 24811 11067
rect 2513 10761 2547 10795
rect 13737 10761 13771 10795
rect 15393 10761 15427 10795
rect 15761 10761 15795 10795
rect 16129 10761 16163 10795
rect 22385 10761 22419 10795
rect 23857 10761 23891 10795
rect 24777 10761 24811 10795
rect 25145 10761 25179 10795
rect 24409 10625 24443 10659
rect 1409 10557 1443 10591
rect 1961 10557 1995 10591
rect 24593 10557 24627 10591
rect 1593 10421 1627 10455
rect 13093 10421 13127 10455
rect 13461 10421 13495 10455
rect 14657 10421 14691 10455
rect 24777 10217 24811 10251
rect 24593 10081 24627 10115
rect 24409 9605 24443 9639
rect 24593 9469 24627 9503
rect 25145 9469 25179 9503
rect 24777 9333 24811 9367
rect 1593 8585 1627 8619
rect 1409 8381 1443 8415
rect 1961 8381 1995 8415
rect 1593 5865 1627 5899
rect 1409 5729 1443 5763
rect 1593 5321 1627 5355
rect 12449 2601 12483 2635
rect 14105 2601 14139 2635
rect 12970 2533 13004 2567
rect 12081 2465 12115 2499
rect 12725 2465 12759 2499
rect 24225 2261 24259 2295
<< metal1 >>
rect 9214 27412 9220 27464
rect 9272 27452 9278 27464
rect 9398 27452 9404 27464
rect 9272 27424 9404 27452
rect 9272 27412 9278 27424
rect 9398 27412 9404 27424
rect 9456 27412 9462 27464
rect 26418 27412 26424 27464
rect 26476 27452 26482 27464
rect 26510 27452 26516 27464
rect 26476 27424 26516 27452
rect 26476 27412 26482 27424
rect 26510 27412 26516 27424
rect 26568 27412 26574 27464
rect 3510 27276 3516 27328
rect 3568 27316 3574 27328
rect 4890 27316 4896 27328
rect 3568 27288 4896 27316
rect 3568 27276 3574 27288
rect 4890 27276 4896 27288
rect 4948 27276 4954 27328
rect 11606 26188 11612 26240
rect 11664 26228 11670 26240
rect 18138 26228 18144 26240
rect 11664 26200 18144 26228
rect 11664 26188 11670 26200
rect 18138 26188 18144 26200
rect 18196 26188 18202 26240
rect 13446 26120 13452 26172
rect 13504 26160 13510 26172
rect 22738 26160 22744 26172
rect 13504 26132 22744 26160
rect 13504 26120 13510 26132
rect 22738 26120 22744 26132
rect 22796 26120 22802 26172
rect 10962 25984 10968 26036
rect 11020 26024 11026 26036
rect 24578 26024 24584 26036
rect 11020 25996 24584 26024
rect 11020 25984 11026 25996
rect 24578 25984 24584 25996
rect 24636 25984 24642 26036
rect 4614 25916 4620 25968
rect 4672 25956 4678 25968
rect 19334 25956 19340 25968
rect 4672 25928 19340 25956
rect 4672 25916 4678 25928
rect 19334 25916 19340 25928
rect 19392 25916 19398 25968
rect 12618 25848 12624 25900
rect 12676 25888 12682 25900
rect 25866 25888 25872 25900
rect 12676 25860 25872 25888
rect 12676 25848 12682 25860
rect 25866 25848 25872 25860
rect 25924 25848 25930 25900
rect 10686 25780 10692 25832
rect 10744 25820 10750 25832
rect 18690 25820 18696 25832
rect 10744 25792 18696 25820
rect 10744 25780 10750 25792
rect 18690 25780 18696 25792
rect 18748 25780 18754 25832
rect 1946 25712 1952 25764
rect 2004 25752 2010 25764
rect 20806 25752 20812 25764
rect 2004 25724 20812 25752
rect 2004 25712 2010 25724
rect 20806 25712 20812 25724
rect 20864 25712 20870 25764
rect 8754 25644 8760 25696
rect 8812 25684 8818 25696
rect 19242 25684 19248 25696
rect 8812 25656 19248 25684
rect 8812 25644 8818 25656
rect 19242 25644 19248 25656
rect 19300 25644 19306 25696
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 2685 25483 2743 25489
rect 2685 25449 2697 25483
rect 2731 25480 2743 25483
rect 2774 25480 2780 25492
rect 2731 25452 2780 25480
rect 2731 25449 2743 25452
rect 2685 25443 2743 25449
rect 2774 25440 2780 25452
rect 2832 25440 2838 25492
rect 8754 25480 8760 25492
rect 8715 25452 8760 25480
rect 8754 25440 8760 25452
rect 8812 25440 8818 25492
rect 10505 25483 10563 25489
rect 10505 25449 10517 25483
rect 10551 25480 10563 25483
rect 10686 25480 10692 25492
rect 10551 25452 10692 25480
rect 10551 25449 10563 25452
rect 10505 25443 10563 25449
rect 10686 25440 10692 25452
rect 10744 25440 10750 25492
rect 11606 25480 11612 25492
rect 11567 25452 11612 25480
rect 11606 25440 11612 25452
rect 11664 25440 11670 25492
rect 11885 25483 11943 25489
rect 11885 25449 11897 25483
rect 11931 25480 11943 25483
rect 24762 25480 24768 25492
rect 11931 25452 24624 25480
rect 24723 25452 24768 25480
rect 11931 25449 11943 25452
rect 11885 25443 11943 25449
rect 8113 25415 8171 25421
rect 8113 25412 8125 25415
rect 7484 25384 8125 25412
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 2314 25344 2320 25356
rect 1443 25316 2320 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 2314 25304 2320 25316
rect 2372 25304 2378 25356
rect 2501 25347 2559 25353
rect 2501 25313 2513 25347
rect 2547 25344 2559 25347
rect 2590 25344 2596 25356
rect 2547 25316 2596 25344
rect 2547 25313 2559 25316
rect 2501 25307 2559 25313
rect 2590 25304 2596 25316
rect 2648 25304 2654 25356
rect 4065 25347 4123 25353
rect 4065 25313 4077 25347
rect 4111 25344 4123 25347
rect 4338 25344 4344 25356
rect 4111 25316 4344 25344
rect 4111 25313 4123 25316
rect 4065 25307 4123 25313
rect 4338 25304 4344 25316
rect 4396 25304 4402 25356
rect 5721 25347 5779 25353
rect 5721 25313 5733 25347
rect 5767 25344 5779 25347
rect 5994 25344 6000 25356
rect 5767 25316 6000 25344
rect 5767 25313 5779 25316
rect 5721 25307 5779 25313
rect 5994 25304 6000 25316
rect 6052 25304 6058 25356
rect 7484 25353 7512 25384
rect 8113 25381 8125 25384
rect 8159 25412 8171 25415
rect 11238 25412 11244 25424
rect 8159 25384 11244 25412
rect 8159 25381 8171 25384
rect 8113 25375 8171 25381
rect 11238 25372 11244 25384
rect 11296 25372 11302 25424
rect 11793 25415 11851 25421
rect 11793 25381 11805 25415
rect 11839 25412 11851 25415
rect 20073 25415 20131 25421
rect 11839 25384 19012 25412
rect 11839 25381 11851 25384
rect 11793 25375 11851 25381
rect 7469 25347 7527 25353
rect 7469 25313 7481 25347
rect 7515 25313 7527 25347
rect 7469 25307 7527 25313
rect 8573 25347 8631 25353
rect 8573 25313 8585 25347
rect 8619 25344 8631 25347
rect 8941 25347 8999 25353
rect 8941 25344 8953 25347
rect 8619 25316 8953 25344
rect 8619 25313 8631 25316
rect 8573 25307 8631 25313
rect 8941 25313 8953 25316
rect 8987 25313 8999 25347
rect 8941 25307 8999 25313
rect 9950 25304 9956 25356
rect 10008 25344 10014 25356
rect 10321 25347 10379 25353
rect 10321 25344 10333 25347
rect 10008 25316 10333 25344
rect 10008 25304 10014 25316
rect 10321 25313 10333 25316
rect 10367 25313 10379 25347
rect 10321 25307 10379 25313
rect 11450 25347 11508 25353
rect 11450 25313 11462 25347
rect 11496 25344 11508 25347
rect 11496 25316 12112 25344
rect 11496 25313 11508 25316
rect 11450 25307 11508 25313
rect 11885 25279 11943 25285
rect 11885 25276 11897 25279
rect 5920 25248 11897 25276
rect 290 25168 296 25220
rect 348 25208 354 25220
rect 5920 25217 5948 25248
rect 11885 25245 11897 25248
rect 11931 25245 11943 25279
rect 11885 25239 11943 25245
rect 4249 25211 4307 25217
rect 4249 25208 4261 25211
rect 348 25180 4261 25208
rect 348 25168 354 25180
rect 4249 25177 4261 25180
rect 4295 25177 4307 25211
rect 4249 25171 4307 25177
rect 5905 25211 5963 25217
rect 5905 25177 5917 25211
rect 5951 25177 5963 25211
rect 5905 25171 5963 25177
rect 7653 25211 7711 25217
rect 7653 25177 7665 25211
rect 7699 25208 7711 25211
rect 11793 25211 11851 25217
rect 11793 25208 11805 25211
rect 7699 25180 11805 25208
rect 7699 25177 7711 25180
rect 7653 25171 7711 25177
rect 11793 25177 11805 25180
rect 11839 25177 11851 25211
rect 11793 25171 11851 25177
rect 1578 25140 1584 25152
rect 1539 25112 1584 25140
rect 1578 25100 1584 25112
rect 1636 25100 1642 25152
rect 6270 25140 6276 25152
rect 6231 25112 6276 25140
rect 6270 25100 6276 25112
rect 6328 25100 6334 25152
rect 7190 25140 7196 25152
rect 7151 25112 7196 25140
rect 7190 25100 7196 25112
rect 7248 25100 7254 25152
rect 8941 25143 8999 25149
rect 8941 25109 8953 25143
rect 8987 25140 8999 25143
rect 9217 25143 9275 25149
rect 9217 25140 9229 25143
rect 8987 25112 9229 25140
rect 8987 25109 8999 25112
rect 8941 25103 8999 25109
rect 9217 25109 9229 25112
rect 9263 25140 9275 25143
rect 9306 25140 9312 25152
rect 9263 25112 9312 25140
rect 9263 25109 9275 25112
rect 9217 25103 9275 25109
rect 9306 25100 9312 25112
rect 9364 25100 9370 25152
rect 10045 25143 10103 25149
rect 10045 25109 10057 25143
rect 10091 25140 10103 25143
rect 11330 25140 11336 25152
rect 10091 25112 11336 25140
rect 10091 25109 10103 25112
rect 10045 25103 10103 25109
rect 11330 25100 11336 25112
rect 11388 25100 11394 25152
rect 12084 25149 12112 25316
rect 12894 25304 12900 25356
rect 12952 25344 12958 25356
rect 12989 25347 13047 25353
rect 12989 25344 13001 25347
rect 12952 25316 13001 25344
rect 12952 25304 12958 25316
rect 12989 25313 13001 25316
rect 13035 25313 13047 25347
rect 12989 25307 13047 25313
rect 13081 25347 13139 25353
rect 13081 25313 13093 25347
rect 13127 25344 13139 25347
rect 13262 25344 13268 25356
rect 13127 25316 13268 25344
rect 13127 25313 13139 25316
rect 13081 25307 13139 25313
rect 13262 25304 13268 25316
rect 13320 25304 13326 25356
rect 14182 25304 14188 25356
rect 14240 25344 14246 25356
rect 14277 25347 14335 25353
rect 14277 25344 14289 25347
rect 14240 25316 14289 25344
rect 14240 25304 14246 25316
rect 14277 25313 14289 25316
rect 14323 25313 14335 25347
rect 14277 25307 14335 25313
rect 16025 25347 16083 25353
rect 16025 25313 16037 25347
rect 16071 25344 16083 25347
rect 16574 25344 16580 25356
rect 16071 25316 16580 25344
rect 16071 25313 16083 25316
rect 16025 25307 16083 25313
rect 16574 25304 16580 25316
rect 16632 25344 16638 25356
rect 17221 25347 17279 25353
rect 17221 25344 17233 25347
rect 16632 25316 17233 25344
rect 16632 25304 16638 25316
rect 17221 25313 17233 25316
rect 17267 25313 17279 25347
rect 17221 25307 17279 25313
rect 18782 25304 18788 25356
rect 18840 25344 18846 25356
rect 18877 25347 18935 25353
rect 18877 25344 18889 25347
rect 18840 25316 18889 25344
rect 18840 25304 18846 25316
rect 18877 25313 18889 25316
rect 18923 25313 18935 25347
rect 18984 25344 19012 25384
rect 20073 25381 20085 25415
rect 20119 25412 20131 25415
rect 22186 25412 22192 25424
rect 20119 25384 22192 25412
rect 20119 25381 20131 25384
rect 20073 25375 20131 25381
rect 22186 25372 22192 25384
rect 22244 25372 22250 25424
rect 22738 25412 22744 25424
rect 22699 25384 22744 25412
rect 22738 25372 22744 25384
rect 22796 25372 22802 25424
rect 24596 25412 24624 25452
rect 24762 25440 24768 25452
rect 24820 25440 24826 25492
rect 27062 25412 27068 25424
rect 24596 25384 27068 25412
rect 27062 25372 27068 25384
rect 27120 25372 27126 25424
rect 20898 25344 20904 25356
rect 18984 25316 20904 25344
rect 18877 25307 18935 25313
rect 20898 25304 20904 25316
rect 20956 25304 20962 25356
rect 21174 25344 21180 25356
rect 21135 25316 21180 25344
rect 21174 25304 21180 25316
rect 21232 25304 21238 25356
rect 22462 25344 22468 25356
rect 22423 25316 22468 25344
rect 22462 25304 22468 25316
rect 22520 25304 22526 25356
rect 24118 25304 24124 25356
rect 24176 25344 24182 25356
rect 24578 25344 24584 25356
rect 24176 25316 24584 25344
rect 24176 25304 24182 25316
rect 24578 25304 24584 25316
rect 24636 25304 24642 25356
rect 12158 25236 12164 25288
rect 12216 25276 12222 25288
rect 13173 25279 13231 25285
rect 13173 25276 13185 25279
rect 12216 25248 13185 25276
rect 12216 25236 12222 25248
rect 13173 25245 13185 25248
rect 13219 25245 13231 25279
rect 13173 25239 13231 25245
rect 15562 25236 15568 25288
rect 15620 25276 15626 25288
rect 16117 25279 16175 25285
rect 16117 25276 16129 25279
rect 15620 25248 16129 25276
rect 15620 25236 15626 25248
rect 16117 25245 16129 25248
rect 16163 25245 16175 25279
rect 16117 25239 16175 25245
rect 16301 25279 16359 25285
rect 16301 25245 16313 25279
rect 16347 25276 16359 25279
rect 16390 25276 16396 25288
rect 16347 25248 16396 25276
rect 16347 25245 16359 25248
rect 16301 25239 16359 25245
rect 16390 25236 16396 25248
rect 16448 25236 16454 25288
rect 17034 25236 17040 25288
rect 17092 25236 17098 25288
rect 18046 25236 18052 25288
rect 18104 25276 18110 25288
rect 18969 25279 19027 25285
rect 18969 25276 18981 25279
rect 18104 25248 18981 25276
rect 18104 25236 18110 25248
rect 18969 25245 18981 25248
rect 19015 25245 19027 25279
rect 19150 25276 19156 25288
rect 19111 25248 19156 25276
rect 18969 25239 19027 25245
rect 19150 25236 19156 25248
rect 19208 25236 19214 25288
rect 21450 25276 21456 25288
rect 21411 25248 21456 25276
rect 21450 25236 21456 25248
rect 21508 25236 21514 25288
rect 12618 25208 12624 25220
rect 12579 25180 12624 25208
rect 12618 25168 12624 25180
rect 12676 25168 12682 25220
rect 14461 25211 14519 25217
rect 14461 25177 14473 25211
rect 14507 25208 14519 25211
rect 17052 25208 17080 25236
rect 14507 25180 17080 25208
rect 14507 25177 14519 25180
rect 14461 25171 14519 25177
rect 17218 25168 17224 25220
rect 17276 25208 17282 25220
rect 25038 25208 25044 25220
rect 17276 25180 25044 25208
rect 17276 25168 17282 25180
rect 25038 25168 25044 25180
rect 25096 25168 25102 25220
rect 12069 25143 12127 25149
rect 12069 25109 12081 25143
rect 12115 25140 12127 25143
rect 12434 25140 12440 25152
rect 12115 25112 12440 25140
rect 12115 25109 12127 25112
rect 12069 25103 12127 25109
rect 12434 25100 12440 25112
rect 12492 25100 12498 25152
rect 13725 25143 13783 25149
rect 13725 25109 13737 25143
rect 13771 25140 13783 25143
rect 14001 25143 14059 25149
rect 14001 25140 14013 25143
rect 13771 25112 14013 25140
rect 13771 25109 13783 25112
rect 13725 25103 13783 25109
rect 14001 25109 14013 25112
rect 14047 25140 14059 25143
rect 14090 25140 14096 25152
rect 14047 25112 14096 25140
rect 14047 25109 14059 25112
rect 14001 25103 14059 25109
rect 14090 25100 14096 25112
rect 14148 25140 14154 25152
rect 14829 25143 14887 25149
rect 14829 25140 14841 25143
rect 14148 25112 14841 25140
rect 14148 25100 14154 25112
rect 14829 25109 14841 25112
rect 14875 25109 14887 25143
rect 14829 25103 14887 25109
rect 15289 25143 15347 25149
rect 15289 25109 15301 25143
rect 15335 25140 15347 25143
rect 15378 25140 15384 25152
rect 15335 25112 15384 25140
rect 15335 25109 15347 25112
rect 15289 25103 15347 25109
rect 15378 25100 15384 25112
rect 15436 25100 15442 25152
rect 15654 25140 15660 25152
rect 15615 25112 15660 25140
rect 15654 25100 15660 25112
rect 15712 25100 15718 25152
rect 16666 25140 16672 25152
rect 16627 25112 16672 25140
rect 16666 25100 16672 25112
rect 16724 25140 16730 25152
rect 17037 25143 17095 25149
rect 17037 25140 17049 25143
rect 16724 25112 17049 25140
rect 16724 25100 16730 25112
rect 17037 25109 17049 25112
rect 17083 25140 17095 25143
rect 17681 25143 17739 25149
rect 17681 25140 17693 25143
rect 17083 25112 17693 25140
rect 17083 25109 17095 25112
rect 17037 25103 17095 25109
rect 17681 25109 17693 25112
rect 17727 25109 17739 25143
rect 17681 25103 17739 25109
rect 18141 25143 18199 25149
rect 18141 25109 18153 25143
rect 18187 25140 18199 25143
rect 18509 25143 18567 25149
rect 18509 25140 18521 25143
rect 18187 25112 18521 25140
rect 18187 25109 18199 25112
rect 18141 25103 18199 25109
rect 18509 25109 18521 25112
rect 18555 25140 18567 25143
rect 18598 25140 18604 25152
rect 18555 25112 18604 25140
rect 18555 25109 18567 25112
rect 18509 25103 18567 25109
rect 18598 25100 18604 25112
rect 18656 25100 18662 25152
rect 19518 25140 19524 25152
rect 19479 25112 19524 25140
rect 19518 25100 19524 25112
rect 19576 25100 19582 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 2682 24936 2688 24948
rect 2643 24908 2688 24936
rect 2682 24896 2688 24908
rect 2740 24896 2746 24948
rect 3786 24936 3792 24948
rect 3747 24908 3792 24936
rect 3786 24896 3792 24908
rect 3844 24896 3850 24948
rect 4890 24936 4896 24948
rect 4851 24908 4896 24936
rect 4890 24896 4896 24908
rect 4948 24896 4954 24948
rect 9306 24896 9312 24948
rect 9364 24936 9370 24948
rect 17218 24936 17224 24948
rect 9364 24908 17224 24936
rect 9364 24896 9370 24908
rect 17218 24896 17224 24908
rect 17276 24896 17282 24948
rect 17773 24939 17831 24945
rect 17773 24936 17785 24939
rect 17328 24908 17785 24936
rect 11885 24871 11943 24877
rect 6840 24840 7604 24868
rect 6641 24803 6699 24809
rect 6641 24769 6653 24803
rect 6687 24800 6699 24803
rect 6840 24800 6868 24840
rect 6687 24772 6868 24800
rect 6687 24769 6699 24772
rect 6641 24763 6699 24769
rect 7190 24760 7196 24812
rect 7248 24800 7254 24812
rect 7576 24809 7604 24840
rect 11885 24837 11897 24871
rect 11931 24868 11943 24871
rect 13354 24868 13360 24880
rect 11931 24840 13360 24868
rect 11931 24837 11943 24840
rect 11885 24831 11943 24837
rect 13354 24828 13360 24840
rect 13412 24828 13418 24880
rect 14918 24828 14924 24880
rect 14976 24868 14982 24880
rect 17328 24868 17356 24908
rect 17773 24905 17785 24908
rect 17819 24936 17831 24939
rect 18046 24936 18052 24948
rect 17819 24908 18052 24936
rect 17819 24905 17831 24908
rect 17773 24899 17831 24905
rect 18046 24896 18052 24908
rect 18104 24896 18110 24948
rect 18141 24939 18199 24945
rect 18141 24905 18153 24939
rect 18187 24936 18199 24939
rect 22462 24936 22468 24948
rect 18187 24908 22468 24936
rect 18187 24905 18199 24908
rect 18141 24899 18199 24905
rect 22462 24896 22468 24908
rect 22520 24936 22526 24948
rect 22925 24939 22983 24945
rect 22925 24936 22937 24939
rect 22520 24908 22937 24936
rect 22520 24896 22526 24908
rect 22925 24905 22937 24908
rect 22971 24905 22983 24939
rect 22925 24899 22983 24905
rect 24118 24896 24124 24948
rect 24176 24936 24182 24948
rect 24397 24939 24455 24945
rect 24397 24936 24409 24939
rect 24176 24908 24409 24936
rect 24176 24896 24182 24908
rect 24397 24905 24409 24908
rect 24443 24905 24455 24939
rect 24397 24899 24455 24905
rect 14976 24840 17356 24868
rect 17420 24840 18736 24868
rect 14976 24828 14982 24840
rect 7377 24803 7435 24809
rect 7377 24800 7389 24803
rect 7248 24772 7389 24800
rect 7248 24760 7254 24772
rect 7377 24769 7389 24772
rect 7423 24769 7435 24803
rect 7377 24763 7435 24769
rect 7561 24803 7619 24809
rect 7561 24769 7573 24803
rect 7607 24800 7619 24803
rect 7607 24772 7972 24800
rect 7607 24769 7619 24772
rect 7561 24763 7619 24769
rect 7944 24744 7972 24772
rect 8386 24760 8392 24812
rect 8444 24800 8450 24812
rect 9033 24803 9091 24809
rect 9033 24800 9045 24803
rect 8444 24772 9045 24800
rect 8444 24760 8450 24772
rect 9033 24769 9045 24772
rect 9079 24800 9091 24803
rect 9490 24800 9496 24812
rect 9079 24772 9496 24800
rect 9079 24769 9091 24772
rect 9033 24763 9091 24769
rect 9490 24760 9496 24772
rect 9548 24760 9554 24812
rect 11238 24800 11244 24812
rect 11199 24772 11244 24800
rect 11238 24760 11244 24772
rect 11296 24760 11302 24812
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24800 13691 24803
rect 16393 24803 16451 24809
rect 13679 24772 14136 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24701 1455 24735
rect 1397 24695 1455 24701
rect 2041 24735 2099 24741
rect 2041 24701 2053 24735
rect 2087 24732 2099 24735
rect 2314 24732 2320 24744
rect 2087 24704 2320 24732
rect 2087 24701 2099 24704
rect 2041 24695 2099 24701
rect 1412 24664 1440 24695
rect 2314 24692 2320 24704
rect 2372 24692 2378 24744
rect 2501 24735 2559 24741
rect 2501 24701 2513 24735
rect 2547 24732 2559 24735
rect 3142 24732 3148 24744
rect 2547 24704 3148 24732
rect 2547 24701 2559 24704
rect 2501 24695 2559 24701
rect 3142 24692 3148 24704
rect 3200 24692 3206 24744
rect 3605 24735 3663 24741
rect 3605 24701 3617 24735
rect 3651 24701 3663 24735
rect 3605 24695 3663 24701
rect 4249 24735 4307 24741
rect 4249 24701 4261 24735
rect 4295 24732 4307 24735
rect 4338 24732 4344 24744
rect 4295 24704 4344 24732
rect 4295 24701 4307 24704
rect 4249 24695 4307 24701
rect 1412 24636 2452 24664
rect 2424 24608 2452 24636
rect 1578 24596 1584 24608
rect 1539 24568 1584 24596
rect 1578 24556 1584 24568
rect 1636 24556 1642 24608
rect 2406 24596 2412 24608
rect 2367 24568 2412 24596
rect 2406 24556 2412 24568
rect 2464 24556 2470 24608
rect 3513 24599 3571 24605
rect 3513 24565 3525 24599
rect 3559 24596 3571 24599
rect 3620 24596 3648 24695
rect 4338 24692 4344 24704
rect 4396 24692 4402 24744
rect 4709 24735 4767 24741
rect 4709 24701 4721 24735
rect 4755 24732 4767 24735
rect 6273 24735 6331 24741
rect 4755 24704 5488 24732
rect 4755 24701 4767 24704
rect 4709 24695 4767 24701
rect 5460 24608 5488 24704
rect 6273 24701 6285 24735
rect 6319 24732 6331 24735
rect 6319 24704 7328 24732
rect 6319 24701 6331 24704
rect 6273 24695 6331 24701
rect 5813 24667 5871 24673
rect 5813 24633 5825 24667
rect 5859 24664 5871 24667
rect 5994 24664 6000 24676
rect 5859 24636 6000 24664
rect 5859 24633 5871 24636
rect 5813 24627 5871 24633
rect 5994 24624 6000 24636
rect 6052 24664 6058 24676
rect 6362 24664 6368 24676
rect 6052 24636 6368 24664
rect 6052 24624 6058 24636
rect 6362 24624 6368 24636
rect 6420 24624 6426 24676
rect 3694 24596 3700 24608
rect 3559 24568 3700 24596
rect 3559 24565 3571 24568
rect 3513 24559 3571 24565
rect 3694 24556 3700 24568
rect 3752 24556 3758 24608
rect 4246 24556 4252 24608
rect 4304 24596 4310 24608
rect 4706 24596 4712 24608
rect 4304 24568 4712 24596
rect 4304 24556 4310 24568
rect 4706 24556 4712 24568
rect 4764 24556 4770 24608
rect 5261 24599 5319 24605
rect 5261 24565 5273 24599
rect 5307 24596 5319 24599
rect 5442 24596 5448 24608
rect 5307 24568 5448 24596
rect 5307 24565 5319 24568
rect 5261 24559 5319 24565
rect 5442 24556 5448 24568
rect 5500 24556 5506 24608
rect 6914 24596 6920 24608
rect 6875 24568 6920 24596
rect 6914 24556 6920 24568
rect 6972 24556 6978 24608
rect 7300 24605 7328 24704
rect 7926 24692 7932 24744
rect 7984 24692 7990 24744
rect 8294 24732 8300 24744
rect 8207 24704 8300 24732
rect 8294 24692 8300 24704
rect 8352 24732 8358 24744
rect 8849 24735 8907 24741
rect 8849 24732 8861 24735
rect 8352 24704 8861 24732
rect 8352 24692 8358 24704
rect 8849 24701 8861 24704
rect 8895 24732 8907 24735
rect 9122 24732 9128 24744
rect 8895 24704 9128 24732
rect 8895 24701 8907 24704
rect 8849 24695 8907 24701
rect 9122 24692 9128 24704
rect 9180 24692 9186 24744
rect 11057 24735 11115 24741
rect 11057 24732 11069 24735
rect 10980 24704 11069 24732
rect 8021 24667 8079 24673
rect 8021 24633 8033 24667
rect 8067 24664 8079 24667
rect 10045 24667 10103 24673
rect 8067 24636 8984 24664
rect 8067 24633 8079 24636
rect 8021 24627 8079 24633
rect 8956 24608 8984 24636
rect 10045 24633 10057 24667
rect 10091 24664 10103 24667
rect 10870 24664 10876 24676
rect 10091 24636 10876 24664
rect 10091 24633 10103 24636
rect 10045 24627 10103 24633
rect 10870 24624 10876 24636
rect 10928 24624 10934 24676
rect 10980 24608 11008 24704
rect 11057 24701 11069 24704
rect 11103 24701 11115 24735
rect 11057 24695 11115 24701
rect 12986 24692 12992 24744
rect 13044 24732 13050 24744
rect 13357 24735 13415 24741
rect 13357 24732 13369 24735
rect 13044 24704 13369 24732
rect 13044 24692 13050 24704
rect 13357 24701 13369 24704
rect 13403 24701 13415 24735
rect 13357 24695 13415 24701
rect 13449 24667 13507 24673
rect 13449 24664 13461 24667
rect 12820 24636 13461 24664
rect 12820 24608 12848 24636
rect 13449 24633 13461 24636
rect 13495 24633 13507 24667
rect 13449 24627 13507 24633
rect 7285 24599 7343 24605
rect 7285 24565 7297 24599
rect 7331 24596 7343 24599
rect 7742 24596 7748 24608
rect 7331 24568 7748 24596
rect 7331 24565 7343 24568
rect 7285 24559 7343 24565
rect 7742 24556 7748 24568
rect 7800 24556 7806 24608
rect 8478 24596 8484 24608
rect 8439 24568 8484 24596
rect 8478 24556 8484 24568
rect 8536 24556 8542 24608
rect 8938 24556 8944 24608
rect 8996 24596 9002 24608
rect 9950 24596 9956 24608
rect 8996 24568 9041 24596
rect 9911 24568 9956 24596
rect 8996 24556 9002 24568
rect 9950 24556 9956 24568
rect 10008 24556 10014 24608
rect 10597 24599 10655 24605
rect 10597 24565 10609 24599
rect 10643 24596 10655 24599
rect 10778 24596 10784 24608
rect 10643 24568 10784 24596
rect 10643 24565 10655 24568
rect 10597 24559 10655 24565
rect 10778 24556 10784 24568
rect 10836 24556 10842 24608
rect 10962 24596 10968 24608
rect 10923 24568 10968 24596
rect 10962 24556 10968 24568
rect 11020 24556 11026 24608
rect 11882 24556 11888 24608
rect 11940 24596 11946 24608
rect 12158 24596 12164 24608
rect 11940 24568 12164 24596
rect 11940 24556 11946 24568
rect 12158 24556 12164 24568
rect 12216 24556 12222 24608
rect 12802 24596 12808 24608
rect 12763 24568 12808 24596
rect 12802 24556 12808 24568
rect 12860 24556 12866 24608
rect 12989 24599 13047 24605
rect 12989 24565 13001 24599
rect 13035 24596 13047 24599
rect 13262 24596 13268 24608
rect 13035 24568 13268 24596
rect 13035 24565 13047 24568
rect 12989 24559 13047 24565
rect 13262 24556 13268 24568
rect 13320 24556 13326 24608
rect 14108 24605 14136 24772
rect 16393 24769 16405 24803
rect 16439 24769 16451 24803
rect 16393 24763 16451 24769
rect 16408 24732 16436 24763
rect 16482 24732 16488 24744
rect 16408 24704 16488 24732
rect 16482 24692 16488 24704
rect 16540 24692 16546 24744
rect 14366 24664 14372 24676
rect 14327 24636 14372 24664
rect 14366 24624 14372 24636
rect 14424 24624 14430 24676
rect 15289 24667 15347 24673
rect 15289 24633 15301 24667
rect 15335 24664 15347 24667
rect 15335 24636 16068 24664
rect 15335 24633 15347 24636
rect 15289 24627 15347 24633
rect 16040 24608 16068 24636
rect 14093 24599 14151 24605
rect 14093 24565 14105 24599
rect 14139 24596 14151 24599
rect 14274 24596 14280 24608
rect 14139 24568 14280 24596
rect 14139 24565 14151 24568
rect 14093 24559 14151 24565
rect 14274 24556 14280 24568
rect 14332 24556 14338 24608
rect 14829 24599 14887 24605
rect 14829 24565 14841 24599
rect 14875 24596 14887 24599
rect 15102 24596 15108 24608
rect 14875 24568 15108 24596
rect 14875 24565 14887 24568
rect 14829 24559 14887 24565
rect 15102 24556 15108 24568
rect 15160 24556 15166 24608
rect 15562 24596 15568 24608
rect 15523 24568 15568 24596
rect 15562 24556 15568 24568
rect 15620 24556 15626 24608
rect 15749 24599 15807 24605
rect 15749 24565 15761 24599
rect 15795 24596 15807 24599
rect 15930 24596 15936 24608
rect 15795 24568 15936 24596
rect 15795 24565 15807 24568
rect 15749 24559 15807 24565
rect 15930 24556 15936 24568
rect 15988 24556 15994 24608
rect 16022 24556 16028 24608
rect 16080 24596 16086 24608
rect 16117 24599 16175 24605
rect 16117 24596 16129 24599
rect 16080 24568 16129 24596
rect 16080 24556 16086 24568
rect 16117 24565 16129 24568
rect 16163 24565 16175 24599
rect 16117 24559 16175 24565
rect 16209 24599 16267 24605
rect 16209 24565 16221 24599
rect 16255 24596 16267 24599
rect 16390 24596 16396 24608
rect 16255 24568 16396 24596
rect 16255 24565 16267 24568
rect 16209 24559 16267 24565
rect 16390 24556 16396 24568
rect 16448 24596 16454 24608
rect 16761 24599 16819 24605
rect 16761 24596 16773 24599
rect 16448 24568 16773 24596
rect 16448 24556 16454 24568
rect 16761 24565 16773 24568
rect 16807 24565 16819 24599
rect 16761 24559 16819 24565
rect 17034 24556 17040 24608
rect 17092 24596 17098 24608
rect 17420 24605 17448 24840
rect 18598 24800 18604 24812
rect 18559 24772 18604 24800
rect 18598 24760 18604 24772
rect 18656 24760 18662 24812
rect 18708 24809 18736 24840
rect 20070 24828 20076 24880
rect 20128 24868 20134 24880
rect 24762 24868 24768 24880
rect 20128 24840 24768 24868
rect 20128 24828 20134 24840
rect 24762 24828 24768 24840
rect 24820 24828 24826 24880
rect 18693 24803 18751 24809
rect 18693 24769 18705 24803
rect 18739 24769 18751 24803
rect 18693 24763 18751 24769
rect 19334 24760 19340 24812
rect 19392 24800 19398 24812
rect 19797 24803 19855 24809
rect 19797 24800 19809 24803
rect 19392 24772 19809 24800
rect 19392 24760 19398 24772
rect 19797 24769 19809 24772
rect 19843 24800 19855 24803
rect 20438 24800 20444 24812
rect 19843 24772 20444 24800
rect 19843 24769 19855 24772
rect 19797 24763 19855 24769
rect 20364 24741 20392 24772
rect 20438 24760 20444 24772
rect 20496 24760 20502 24812
rect 20530 24760 20536 24812
rect 20588 24800 20594 24812
rect 20625 24803 20683 24809
rect 20625 24800 20637 24803
rect 20588 24772 20637 24800
rect 20588 24760 20594 24772
rect 20625 24769 20637 24772
rect 20671 24800 20683 24803
rect 20993 24803 21051 24809
rect 20993 24800 21005 24803
rect 20671 24772 21005 24800
rect 20671 24769 20683 24772
rect 20625 24763 20683 24769
rect 20993 24769 21005 24772
rect 21039 24769 21051 24803
rect 20993 24763 21051 24769
rect 24854 24760 24860 24812
rect 24912 24800 24918 24812
rect 26050 24800 26056 24812
rect 24912 24772 26056 24800
rect 24912 24760 24918 24772
rect 26050 24760 26056 24772
rect 26108 24760 26114 24812
rect 20349 24735 20407 24741
rect 20349 24701 20361 24735
rect 20395 24701 20407 24735
rect 20349 24695 20407 24701
rect 22189 24735 22247 24741
rect 22189 24701 22201 24735
rect 22235 24701 22247 24735
rect 22189 24695 22247 24701
rect 20162 24624 20168 24676
rect 20220 24664 20226 24676
rect 20441 24667 20499 24673
rect 20441 24664 20453 24667
rect 20220 24636 20453 24664
rect 20220 24624 20226 24636
rect 20441 24633 20453 24636
rect 20487 24633 20499 24667
rect 20441 24627 20499 24633
rect 17405 24599 17463 24605
rect 17405 24596 17417 24599
rect 17092 24568 17417 24596
rect 17092 24556 17098 24568
rect 17405 24565 17417 24568
rect 17451 24565 17463 24599
rect 17405 24559 17463 24565
rect 18509 24599 18567 24605
rect 18509 24565 18521 24599
rect 18555 24596 18567 24599
rect 18598 24596 18604 24608
rect 18555 24568 18604 24596
rect 18555 24565 18567 24568
rect 18509 24559 18567 24565
rect 18598 24556 18604 24568
rect 18656 24556 18662 24608
rect 18782 24556 18788 24608
rect 18840 24596 18846 24608
rect 19153 24599 19211 24605
rect 19153 24596 19165 24599
rect 18840 24568 19165 24596
rect 18840 24556 18846 24568
rect 19153 24565 19165 24568
rect 19199 24565 19211 24599
rect 19978 24596 19984 24608
rect 19939 24568 19984 24596
rect 19153 24559 19211 24565
rect 19978 24556 19984 24568
rect 20036 24556 20042 24608
rect 20714 24556 20720 24608
rect 20772 24596 20778 24608
rect 21174 24596 21180 24608
rect 20772 24568 21180 24596
rect 20772 24556 20778 24568
rect 21174 24556 21180 24568
rect 21232 24596 21238 24608
rect 21361 24599 21419 24605
rect 21361 24596 21373 24599
rect 21232 24568 21373 24596
rect 21232 24556 21238 24568
rect 21361 24565 21373 24568
rect 21407 24565 21419 24599
rect 21361 24559 21419 24565
rect 22097 24599 22155 24605
rect 22097 24565 22109 24599
rect 22143 24596 22155 24599
rect 22204 24596 22232 24695
rect 24026 24692 24032 24744
rect 24084 24732 24090 24744
rect 24581 24735 24639 24741
rect 24581 24732 24593 24735
rect 24084 24704 24593 24732
rect 24084 24692 24090 24704
rect 24581 24701 24593 24704
rect 24627 24732 24639 24735
rect 25133 24735 25191 24741
rect 25133 24732 25145 24735
rect 24627 24704 25145 24732
rect 24627 24701 24639 24704
rect 24581 24695 24639 24701
rect 25133 24701 25145 24704
rect 25179 24701 25191 24735
rect 25133 24695 25191 24701
rect 22465 24667 22523 24673
rect 22465 24633 22477 24667
rect 22511 24664 22523 24667
rect 23106 24664 23112 24676
rect 22511 24636 23112 24664
rect 22511 24633 22523 24636
rect 22465 24627 22523 24633
rect 23106 24624 23112 24636
rect 23164 24624 23170 24676
rect 23382 24596 23388 24608
rect 22143 24568 23388 24596
rect 22143 24565 22155 24568
rect 22097 24559 22155 24565
rect 23382 24556 23388 24568
rect 23440 24556 23446 24608
rect 24670 24556 24676 24608
rect 24728 24596 24734 24608
rect 24765 24599 24823 24605
rect 24765 24596 24777 24599
rect 24728 24568 24777 24596
rect 24728 24556 24734 24568
rect 24765 24565 24777 24568
rect 24811 24565 24823 24599
rect 24765 24559 24823 24565
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 4154 24352 4160 24404
rect 4212 24392 4218 24404
rect 4249 24395 4307 24401
rect 4249 24392 4261 24395
rect 4212 24364 4261 24392
rect 4212 24352 4218 24364
rect 4249 24361 4261 24364
rect 4295 24361 4307 24395
rect 4249 24355 4307 24361
rect 7190 24352 7196 24404
rect 7248 24392 7254 24404
rect 7837 24395 7895 24401
rect 7837 24392 7849 24395
rect 7248 24364 7849 24392
rect 7248 24352 7254 24364
rect 7837 24361 7849 24364
rect 7883 24361 7895 24395
rect 7837 24355 7895 24361
rect 8205 24395 8263 24401
rect 8205 24361 8217 24395
rect 8251 24392 8263 24395
rect 8478 24392 8484 24404
rect 8251 24364 8484 24392
rect 8251 24361 8263 24364
rect 8205 24355 8263 24361
rect 8478 24352 8484 24364
rect 8536 24392 8542 24404
rect 9217 24395 9275 24401
rect 9217 24392 9229 24395
rect 8536 24364 9229 24392
rect 8536 24352 8542 24364
rect 9217 24361 9229 24364
rect 9263 24361 9275 24395
rect 9217 24355 9275 24361
rect 9677 24395 9735 24401
rect 9677 24361 9689 24395
rect 9723 24361 9735 24395
rect 9677 24355 9735 24361
rect 5896 24327 5954 24333
rect 5896 24293 5908 24327
rect 5942 24324 5954 24327
rect 6546 24324 6552 24336
rect 5942 24296 6552 24324
rect 5942 24293 5954 24296
rect 5896 24287 5954 24293
rect 6546 24284 6552 24296
rect 6604 24284 6610 24336
rect 8297 24327 8355 24333
rect 8297 24293 8309 24327
rect 8343 24324 8355 24327
rect 9030 24324 9036 24336
rect 8343 24296 9036 24324
rect 8343 24293 8355 24296
rect 8297 24287 8355 24293
rect 9030 24284 9036 24296
rect 9088 24324 9094 24336
rect 9692 24324 9720 24355
rect 9766 24352 9772 24404
rect 9824 24392 9830 24404
rect 10045 24395 10103 24401
rect 10045 24392 10057 24395
rect 9824 24364 10057 24392
rect 9824 24352 9830 24364
rect 10045 24361 10057 24364
rect 10091 24361 10103 24395
rect 10045 24355 10103 24361
rect 11241 24395 11299 24401
rect 11241 24361 11253 24395
rect 11287 24392 11299 24395
rect 11330 24392 11336 24404
rect 11287 24364 11336 24392
rect 11287 24361 11299 24364
rect 11241 24355 11299 24361
rect 11330 24352 11336 24364
rect 11388 24352 11394 24404
rect 13630 24392 13636 24404
rect 13591 24364 13636 24392
rect 13630 24352 13636 24364
rect 13688 24352 13694 24404
rect 14090 24352 14096 24404
rect 14148 24392 14154 24404
rect 14645 24395 14703 24401
rect 14645 24392 14657 24395
rect 14148 24364 14657 24392
rect 14148 24352 14154 24364
rect 14645 24361 14657 24364
rect 14691 24392 14703 24395
rect 14826 24392 14832 24404
rect 14691 24364 14832 24392
rect 14691 24361 14703 24364
rect 14645 24355 14703 24361
rect 14826 24352 14832 24364
rect 14884 24352 14890 24404
rect 15470 24392 15476 24404
rect 15431 24364 15476 24392
rect 15470 24352 15476 24364
rect 15528 24352 15534 24404
rect 16574 24392 16580 24404
rect 16535 24364 16580 24392
rect 16574 24352 16580 24364
rect 16632 24352 16638 24404
rect 18049 24395 18107 24401
rect 18049 24361 18061 24395
rect 18095 24392 18107 24395
rect 19242 24392 19248 24404
rect 18095 24364 19248 24392
rect 18095 24361 18107 24364
rect 18049 24355 18107 24361
rect 19242 24352 19248 24364
rect 19300 24352 19306 24404
rect 19518 24392 19524 24404
rect 19479 24364 19524 24392
rect 19518 24352 19524 24364
rect 19576 24352 19582 24404
rect 19889 24395 19947 24401
rect 19889 24361 19901 24395
rect 19935 24392 19947 24395
rect 20070 24392 20076 24404
rect 19935 24364 20076 24392
rect 19935 24361 19947 24364
rect 19889 24355 19947 24361
rect 20070 24352 20076 24364
rect 20128 24352 20134 24404
rect 20162 24352 20168 24404
rect 20220 24392 20226 24404
rect 20257 24395 20315 24401
rect 20257 24392 20269 24395
rect 20220 24364 20269 24392
rect 20220 24352 20226 24364
rect 20257 24361 20269 24364
rect 20303 24361 20315 24395
rect 25498 24392 25504 24404
rect 25459 24364 25504 24392
rect 20257 24355 20315 24361
rect 25498 24352 25504 24364
rect 25556 24352 25562 24404
rect 9088 24296 9720 24324
rect 9088 24284 9094 24296
rect 9858 24284 9864 24336
rect 9916 24324 9922 24336
rect 10137 24327 10195 24333
rect 10137 24324 10149 24327
rect 9916 24296 10149 24324
rect 9916 24284 9922 24296
rect 10137 24293 10149 24296
rect 10183 24293 10195 24327
rect 14844 24324 14872 24352
rect 16390 24324 16396 24336
rect 14844 24296 16396 24324
rect 10137 24287 10195 24293
rect 16390 24284 16396 24296
rect 16448 24324 16454 24336
rect 16666 24324 16672 24336
rect 16448 24296 16672 24324
rect 16448 24284 16454 24296
rect 16666 24284 16672 24296
rect 16724 24324 16730 24336
rect 16853 24327 16911 24333
rect 16853 24324 16865 24327
rect 16724 24296 16865 24324
rect 16724 24284 16730 24296
rect 16853 24293 16865 24296
rect 16899 24293 16911 24327
rect 16853 24287 16911 24293
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 1762 24256 1768 24268
rect 1443 24228 1768 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 1762 24216 1768 24228
rect 1820 24216 1826 24268
rect 2501 24259 2559 24265
rect 2501 24225 2513 24259
rect 2547 24256 2559 24259
rect 3234 24256 3240 24268
rect 2547 24228 3240 24256
rect 2547 24225 2559 24228
rect 2501 24219 2559 24225
rect 3234 24216 3240 24228
rect 3292 24216 3298 24268
rect 4065 24259 4123 24265
rect 4065 24225 4077 24259
rect 4111 24256 4123 24259
rect 4614 24256 4620 24268
rect 4111 24228 4620 24256
rect 4111 24225 4123 24228
rect 4065 24219 4123 24225
rect 4614 24216 4620 24228
rect 4672 24216 4678 24268
rect 5534 24216 5540 24268
rect 5592 24256 5598 24268
rect 5629 24259 5687 24265
rect 5629 24256 5641 24259
rect 5592 24228 5641 24256
rect 5592 24216 5598 24228
rect 5629 24225 5641 24228
rect 5675 24256 5687 24259
rect 6270 24256 6276 24268
rect 5675 24228 6276 24256
rect 5675 24225 5687 24228
rect 5629 24219 5687 24225
rect 6270 24216 6276 24228
rect 6328 24216 6334 24268
rect 12066 24256 12072 24268
rect 12027 24228 12072 24256
rect 12066 24216 12072 24228
rect 12124 24216 12130 24268
rect 13725 24259 13783 24265
rect 13725 24225 13737 24259
rect 13771 24256 13783 24259
rect 14090 24256 14096 24268
rect 13771 24228 14096 24256
rect 13771 24225 13783 24228
rect 13725 24219 13783 24225
rect 14090 24216 14096 24228
rect 14148 24216 14154 24268
rect 15286 24216 15292 24268
rect 15344 24256 15350 24268
rect 15654 24256 15660 24268
rect 15344 24228 15660 24256
rect 15344 24216 15350 24228
rect 15654 24216 15660 24228
rect 15712 24256 15718 24268
rect 15841 24259 15899 24265
rect 15841 24256 15853 24259
rect 15712 24228 15853 24256
rect 15712 24216 15718 24228
rect 15841 24225 15853 24228
rect 15887 24225 15899 24259
rect 15841 24219 15899 24225
rect 17589 24259 17647 24265
rect 17589 24225 17601 24259
rect 17635 24256 17647 24259
rect 18046 24256 18052 24268
rect 17635 24228 18052 24256
rect 17635 24225 17647 24228
rect 17589 24219 17647 24225
rect 18046 24216 18052 24228
rect 18104 24256 18110 24268
rect 18417 24259 18475 24265
rect 18417 24256 18429 24259
rect 18104 24228 18429 24256
rect 18104 24216 18110 24228
rect 18417 24225 18429 24228
rect 18463 24225 18475 24259
rect 18417 24219 18475 24225
rect 19334 24216 19340 24268
rect 19392 24256 19398 24268
rect 19705 24259 19763 24265
rect 19705 24256 19717 24259
rect 19392 24228 19717 24256
rect 19392 24216 19398 24228
rect 19705 24225 19717 24228
rect 19751 24225 19763 24259
rect 19705 24219 19763 24225
rect 21082 24216 21088 24268
rect 21140 24256 21146 24268
rect 21269 24259 21327 24265
rect 21269 24256 21281 24259
rect 21140 24228 21281 24256
rect 21140 24216 21146 24228
rect 21269 24225 21281 24228
rect 21315 24225 21327 24259
rect 22830 24256 22836 24268
rect 22791 24228 22836 24256
rect 21269 24219 21327 24225
rect 22830 24216 22836 24228
rect 22888 24216 22894 24268
rect 23934 24216 23940 24268
rect 23992 24256 23998 24268
rect 24029 24259 24087 24265
rect 24029 24256 24041 24259
rect 23992 24228 24041 24256
rect 23992 24216 23998 24228
rect 24029 24225 24041 24228
rect 24075 24256 24087 24259
rect 24854 24256 24860 24268
rect 24075 24228 24860 24256
rect 24075 24225 24087 24228
rect 24029 24219 24087 24225
rect 24854 24216 24860 24228
rect 24912 24216 24918 24268
rect 25317 24259 25375 24265
rect 25317 24225 25329 24259
rect 25363 24256 25375 24259
rect 25774 24256 25780 24268
rect 25363 24228 25780 24256
rect 25363 24225 25375 24228
rect 25317 24219 25375 24225
rect 25774 24216 25780 24228
rect 25832 24216 25838 24268
rect 2774 24148 2780 24200
rect 2832 24188 2838 24200
rect 3053 24191 3111 24197
rect 3053 24188 3065 24191
rect 2832 24160 3065 24188
rect 2832 24148 2838 24160
rect 3053 24157 3065 24160
rect 3099 24157 3111 24191
rect 3053 24151 3111 24157
rect 4338 24148 4344 24200
rect 4396 24188 4402 24200
rect 4798 24188 4804 24200
rect 4396 24160 4804 24188
rect 4396 24148 4402 24160
rect 4798 24148 4804 24160
rect 4856 24148 4862 24200
rect 8389 24191 8447 24197
rect 8389 24188 8401 24191
rect 8128 24160 8401 24188
rect 6914 24080 6920 24132
rect 6972 24120 6978 24132
rect 7285 24123 7343 24129
rect 7285 24120 7297 24123
rect 6972 24092 7297 24120
rect 6972 24080 6978 24092
rect 7285 24089 7297 24092
rect 7331 24089 7343 24123
rect 7285 24083 7343 24089
rect 8128 24064 8156 24160
rect 8389 24157 8401 24160
rect 8435 24157 8447 24191
rect 8389 24151 8447 24157
rect 9490 24148 9496 24200
rect 9548 24188 9554 24200
rect 10229 24191 10287 24197
rect 10229 24188 10241 24191
rect 9548 24160 10241 24188
rect 9548 24148 9554 24160
rect 10229 24157 10241 24160
rect 10275 24188 10287 24191
rect 11422 24188 11428 24200
rect 10275 24160 11428 24188
rect 10275 24157 10287 24160
rect 10229 24151 10287 24157
rect 11422 24148 11428 24160
rect 11480 24148 11486 24200
rect 12161 24191 12219 24197
rect 12161 24157 12173 24191
rect 12207 24157 12219 24191
rect 12161 24151 12219 24157
rect 11054 24080 11060 24132
rect 11112 24120 11118 24132
rect 11517 24123 11575 24129
rect 11517 24120 11529 24123
rect 11112 24092 11529 24120
rect 11112 24080 11118 24092
rect 11517 24089 11529 24092
rect 11563 24120 11575 24123
rect 12176 24120 12204 24151
rect 12250 24148 12256 24200
rect 12308 24188 12314 24200
rect 13909 24191 13967 24197
rect 12308 24160 12353 24188
rect 12308 24148 12314 24160
rect 13909 24157 13921 24191
rect 13955 24157 13967 24191
rect 13909 24151 13967 24157
rect 11563 24092 12204 24120
rect 13924 24120 13952 24151
rect 14182 24148 14188 24200
rect 14240 24188 14246 24200
rect 14369 24191 14427 24197
rect 14369 24188 14381 24191
rect 14240 24160 14381 24188
rect 14240 24148 14246 24160
rect 14369 24157 14381 24160
rect 14415 24188 14427 24191
rect 14642 24188 14648 24200
rect 14415 24160 14648 24188
rect 14415 24157 14427 24160
rect 14369 24151 14427 24157
rect 14642 24148 14648 24160
rect 14700 24148 14706 24200
rect 15930 24188 15936 24200
rect 15891 24160 15936 24188
rect 15930 24148 15936 24160
rect 15988 24148 15994 24200
rect 16025 24191 16083 24197
rect 16025 24157 16037 24191
rect 16071 24157 16083 24191
rect 16025 24151 16083 24157
rect 17037 24191 17095 24197
rect 17037 24157 17049 24191
rect 17083 24188 17095 24191
rect 17862 24188 17868 24200
rect 17083 24160 17868 24188
rect 17083 24157 17095 24160
rect 17037 24151 17095 24157
rect 14734 24120 14740 24132
rect 13924 24092 14740 24120
rect 11563 24089 11575 24092
rect 11517 24083 11575 24089
rect 14734 24080 14740 24092
rect 14792 24080 14798 24132
rect 15838 24080 15844 24132
rect 15896 24120 15902 24132
rect 16040 24120 16068 24151
rect 17862 24148 17868 24160
rect 17920 24148 17926 24200
rect 18506 24188 18512 24200
rect 18467 24160 18512 24188
rect 18506 24148 18512 24160
rect 18564 24148 18570 24200
rect 18690 24188 18696 24200
rect 18651 24160 18696 24188
rect 18690 24148 18696 24160
rect 18748 24148 18754 24200
rect 20806 24148 20812 24200
rect 20864 24188 20870 24200
rect 21361 24191 21419 24197
rect 21361 24188 21373 24191
rect 20864 24160 21373 24188
rect 20864 24148 20870 24160
rect 21361 24157 21373 24160
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 21545 24191 21603 24197
rect 21545 24157 21557 24191
rect 21591 24188 21603 24191
rect 21591 24160 22232 24188
rect 21591 24157 21603 24160
rect 21545 24151 21603 24157
rect 15896 24092 16068 24120
rect 15896 24080 15902 24092
rect 19242 24080 19248 24132
rect 19300 24120 19306 24132
rect 19518 24120 19524 24132
rect 19300 24092 19524 24120
rect 19300 24080 19306 24092
rect 19518 24080 19524 24092
rect 19576 24120 19582 24132
rect 20346 24120 20352 24132
rect 19576 24092 20352 24120
rect 19576 24080 19582 24092
rect 20346 24080 20352 24092
rect 20404 24120 20410 24132
rect 20625 24123 20683 24129
rect 20625 24120 20637 24123
rect 20404 24092 20637 24120
rect 20404 24080 20410 24092
rect 20625 24089 20637 24092
rect 20671 24120 20683 24123
rect 21634 24120 21640 24132
rect 20671 24092 21640 24120
rect 20671 24089 20683 24092
rect 20625 24083 20683 24089
rect 21634 24080 21640 24092
rect 21692 24120 21698 24132
rect 21913 24123 21971 24129
rect 21913 24120 21925 24123
rect 21692 24092 21925 24120
rect 21692 24080 21698 24092
rect 21913 24089 21925 24092
rect 21959 24089 21971 24123
rect 22204 24120 22232 24160
rect 22278 24148 22284 24200
rect 22336 24188 22342 24200
rect 22925 24191 22983 24197
rect 22925 24188 22937 24191
rect 22336 24160 22937 24188
rect 22336 24148 22342 24160
rect 22925 24157 22937 24160
rect 22971 24157 22983 24191
rect 22925 24151 22983 24157
rect 23014 24148 23020 24200
rect 23072 24188 23078 24200
rect 23072 24160 23117 24188
rect 23072 24148 23078 24160
rect 23474 24148 23480 24200
rect 23532 24188 23538 24200
rect 24213 24191 24271 24197
rect 24213 24188 24225 24191
rect 23532 24160 24225 24188
rect 23532 24148 23538 24160
rect 24213 24157 24225 24160
rect 24259 24157 24271 24191
rect 24213 24151 24271 24157
rect 22370 24120 22376 24132
rect 22204 24092 22376 24120
rect 21913 24083 21971 24089
rect 1394 24012 1400 24064
rect 1452 24052 1458 24064
rect 1581 24055 1639 24061
rect 1581 24052 1593 24055
rect 1452 24024 1593 24052
rect 1452 24012 1458 24024
rect 1581 24021 1593 24024
rect 1627 24021 1639 24055
rect 1581 24015 1639 24021
rect 1762 24012 1768 24064
rect 1820 24052 1826 24064
rect 1949 24055 2007 24061
rect 1949 24052 1961 24055
rect 1820 24024 1961 24052
rect 1820 24012 1826 24024
rect 1949 24021 1961 24024
rect 1995 24021 2007 24055
rect 1949 24015 2007 24021
rect 2685 24055 2743 24061
rect 2685 24021 2697 24055
rect 2731 24052 2743 24055
rect 2774 24052 2780 24064
rect 2731 24024 2780 24052
rect 2731 24021 2743 24024
rect 2685 24015 2743 24021
rect 2774 24012 2780 24024
rect 2832 24012 2838 24064
rect 4890 24052 4896 24064
rect 4851 24024 4896 24052
rect 4890 24012 4896 24024
rect 4948 24012 4954 24064
rect 5258 24052 5264 24064
rect 5219 24024 5264 24052
rect 5258 24012 5264 24024
rect 5316 24012 5322 24064
rect 7006 24052 7012 24064
rect 6919 24024 7012 24052
rect 7006 24012 7012 24024
rect 7064 24052 7070 24064
rect 7650 24052 7656 24064
rect 7064 24024 7656 24052
rect 7064 24012 7070 24024
rect 7650 24012 7656 24024
rect 7708 24012 7714 24064
rect 7745 24055 7803 24061
rect 7745 24021 7757 24055
rect 7791 24052 7803 24055
rect 8110 24052 8116 24064
rect 7791 24024 8116 24052
rect 7791 24021 7803 24024
rect 7745 24015 7803 24021
rect 8110 24012 8116 24024
rect 8168 24012 8174 24064
rect 8938 24052 8944 24064
rect 8899 24024 8944 24052
rect 8938 24012 8944 24024
rect 8996 24012 9002 24064
rect 10686 24052 10692 24064
rect 10647 24024 10692 24052
rect 10686 24012 10692 24024
rect 10744 24012 10750 24064
rect 11701 24055 11759 24061
rect 11701 24021 11713 24055
rect 11747 24052 11759 24055
rect 12342 24052 12348 24064
rect 11747 24024 12348 24052
rect 11747 24021 11759 24024
rect 11701 24015 11759 24021
rect 12342 24012 12348 24024
rect 12400 24012 12406 24064
rect 12986 24052 12992 24064
rect 12947 24024 12992 24052
rect 12986 24012 12992 24024
rect 13044 24012 13050 24064
rect 13265 24055 13323 24061
rect 13265 24021 13277 24055
rect 13311 24052 13323 24055
rect 13722 24052 13728 24064
rect 13311 24024 13728 24052
rect 13311 24021 13323 24024
rect 13265 24015 13323 24021
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 15105 24055 15163 24061
rect 15105 24021 15117 24055
rect 15151 24052 15163 24055
rect 15470 24052 15476 24064
rect 15151 24024 15476 24052
rect 15151 24021 15163 24024
rect 15105 24015 15163 24021
rect 15470 24012 15476 24024
rect 15528 24012 15534 24064
rect 17957 24055 18015 24061
rect 17957 24021 17969 24055
rect 18003 24052 18015 24055
rect 18598 24052 18604 24064
rect 18003 24024 18604 24052
rect 18003 24021 18015 24024
rect 17957 24015 18015 24021
rect 18598 24012 18604 24024
rect 18656 24012 18662 24064
rect 19150 24052 19156 24064
rect 19111 24024 19156 24052
rect 19150 24012 19156 24024
rect 19208 24012 19214 24064
rect 20714 24012 20720 24064
rect 20772 24052 20778 24064
rect 20901 24055 20959 24061
rect 20901 24052 20913 24055
rect 20772 24024 20913 24052
rect 20772 24012 20778 24024
rect 20901 24021 20913 24024
rect 20947 24021 20959 24055
rect 21928 24052 21956 24083
rect 22370 24080 22376 24092
rect 22428 24080 22434 24132
rect 22281 24055 22339 24061
rect 22281 24052 22293 24055
rect 21928 24024 22293 24052
rect 20901 24015 20959 24021
rect 22281 24021 22293 24024
rect 22327 24021 22339 24055
rect 22281 24015 22339 24021
rect 22465 24055 22523 24061
rect 22465 24021 22477 24055
rect 22511 24052 22523 24055
rect 23566 24052 23572 24064
rect 22511 24024 23572 24052
rect 22511 24021 22523 24024
rect 22465 24015 22523 24021
rect 23566 24012 23572 24024
rect 23624 24012 23630 24064
rect 23753 24055 23811 24061
rect 23753 24021 23765 24055
rect 23799 24052 23811 24055
rect 24118 24052 24124 24064
rect 23799 24024 24124 24052
rect 23799 24021 23811 24024
rect 23753 24015 23811 24021
rect 24118 24012 24124 24024
rect 24176 24012 24182 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2130 23808 2136 23860
rect 2188 23848 2194 23860
rect 2682 23848 2688 23860
rect 2188 23820 2688 23848
rect 2188 23808 2194 23820
rect 2682 23808 2688 23820
rect 2740 23808 2746 23860
rect 3145 23851 3203 23857
rect 3145 23817 3157 23851
rect 3191 23848 3203 23851
rect 3234 23848 3240 23860
rect 3191 23820 3240 23848
rect 3191 23817 3203 23820
rect 3145 23811 3203 23817
rect 3234 23808 3240 23820
rect 3292 23808 3298 23860
rect 3786 23848 3792 23860
rect 3747 23820 3792 23848
rect 3786 23808 3792 23820
rect 3844 23808 3850 23860
rect 4614 23848 4620 23860
rect 4575 23820 4620 23848
rect 4614 23808 4620 23820
rect 4672 23848 4678 23860
rect 5074 23848 5080 23860
rect 4672 23820 5080 23848
rect 4672 23808 4678 23820
rect 5074 23808 5080 23820
rect 5132 23808 5138 23860
rect 8294 23848 8300 23860
rect 8255 23820 8300 23848
rect 8294 23808 8300 23820
rect 8352 23848 8358 23860
rect 8846 23848 8852 23860
rect 8352 23820 8852 23848
rect 8352 23808 8358 23820
rect 8846 23808 8852 23820
rect 8904 23808 8910 23860
rect 9766 23808 9772 23860
rect 9824 23848 9830 23860
rect 11057 23851 11115 23857
rect 11057 23848 11069 23851
rect 9824 23820 11069 23848
rect 9824 23808 9830 23820
rect 11057 23817 11069 23820
rect 11103 23817 11115 23851
rect 11422 23848 11428 23860
rect 11383 23820 11428 23848
rect 11057 23811 11115 23817
rect 11422 23808 11428 23820
rect 11480 23808 11486 23860
rect 12250 23848 12256 23860
rect 12211 23820 12256 23848
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 15105 23851 15163 23857
rect 15105 23817 15117 23851
rect 15151 23848 15163 23851
rect 15838 23848 15844 23860
rect 15151 23820 15844 23848
rect 15151 23817 15163 23820
rect 15105 23811 15163 23817
rect 15838 23808 15844 23820
rect 15896 23808 15902 23860
rect 15930 23808 15936 23860
rect 15988 23848 15994 23860
rect 16853 23851 16911 23857
rect 16853 23848 16865 23851
rect 15988 23820 16865 23848
rect 15988 23808 15994 23820
rect 16853 23817 16865 23820
rect 16899 23817 16911 23851
rect 16853 23811 16911 23817
rect 17865 23851 17923 23857
rect 17865 23817 17877 23851
rect 17911 23848 17923 23851
rect 18690 23848 18696 23860
rect 17911 23820 18696 23848
rect 17911 23817 17923 23820
rect 17865 23811 17923 23817
rect 18690 23808 18696 23820
rect 18748 23848 18754 23860
rect 19429 23851 19487 23857
rect 19429 23848 19441 23851
rect 18748 23820 19441 23848
rect 18748 23808 18754 23820
rect 19429 23817 19441 23820
rect 19475 23817 19487 23851
rect 19429 23811 19487 23817
rect 22097 23851 22155 23857
rect 22097 23817 22109 23851
rect 22143 23848 22155 23851
rect 22370 23848 22376 23860
rect 22143 23820 22376 23848
rect 22143 23817 22155 23820
rect 22097 23811 22155 23817
rect 22370 23808 22376 23820
rect 22428 23808 22434 23860
rect 24026 23848 24032 23860
rect 23400 23820 24032 23848
rect 6825 23783 6883 23789
rect 6825 23780 6837 23783
rect 5644 23752 6837 23780
rect 5258 23672 5264 23724
rect 5316 23712 5322 23724
rect 5644 23721 5672 23752
rect 6825 23749 6837 23752
rect 6871 23749 6883 23783
rect 8389 23783 8447 23789
rect 8389 23780 8401 23783
rect 6825 23743 6883 23749
rect 7300 23752 8401 23780
rect 7300 23724 7328 23752
rect 8389 23749 8401 23752
rect 8435 23749 8447 23783
rect 8389 23743 8447 23749
rect 10045 23783 10103 23789
rect 10045 23749 10057 23783
rect 10091 23780 10103 23783
rect 10870 23780 10876 23792
rect 10091 23752 10876 23780
rect 10091 23749 10103 23752
rect 10045 23743 10103 23749
rect 10870 23740 10876 23752
rect 10928 23740 10934 23792
rect 5629 23715 5687 23721
rect 5629 23712 5641 23715
rect 5316 23684 5641 23712
rect 5316 23672 5322 23684
rect 5629 23681 5641 23684
rect 5675 23681 5687 23715
rect 5629 23675 5687 23681
rect 5813 23715 5871 23721
rect 5813 23681 5825 23715
rect 5859 23712 5871 23715
rect 7006 23712 7012 23724
rect 5859 23684 7012 23712
rect 5859 23681 5871 23684
rect 5813 23675 5871 23681
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 2409 23647 2467 23653
rect 1443 23616 1992 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 1964 23520 1992 23616
rect 2409 23613 2421 23647
rect 2455 23644 2467 23647
rect 2498 23644 2504 23656
rect 2455 23616 2504 23644
rect 2455 23613 2467 23616
rect 2409 23607 2467 23613
rect 2498 23604 2504 23616
rect 2556 23604 2562 23656
rect 3605 23647 3663 23653
rect 3605 23613 3617 23647
rect 3651 23644 3663 23647
rect 4249 23647 4307 23653
rect 4249 23644 4261 23647
rect 3651 23616 4261 23644
rect 3651 23613 3663 23616
rect 3605 23607 3663 23613
rect 4249 23613 4261 23616
rect 4295 23644 4307 23647
rect 4522 23644 4528 23656
rect 4295 23616 4528 23644
rect 4295 23613 4307 23616
rect 4249 23607 4307 23613
rect 4522 23604 4528 23616
rect 4580 23604 4586 23656
rect 4890 23604 4896 23656
rect 4948 23644 4954 23656
rect 5537 23647 5595 23653
rect 5537 23644 5549 23647
rect 4948 23616 5549 23644
rect 4948 23604 4954 23616
rect 5537 23613 5549 23616
rect 5583 23613 5595 23647
rect 5537 23607 5595 23613
rect 5077 23579 5135 23585
rect 5077 23545 5089 23579
rect 5123 23576 5135 23579
rect 5828 23576 5856 23675
rect 7006 23672 7012 23684
rect 7064 23672 7070 23724
rect 7282 23712 7288 23724
rect 7195 23684 7288 23712
rect 7282 23672 7288 23684
rect 7340 23672 7346 23724
rect 7377 23715 7435 23721
rect 7377 23681 7389 23715
rect 7423 23681 7435 23715
rect 7377 23675 7435 23681
rect 6546 23604 6552 23656
rect 6604 23644 6610 23656
rect 7392 23644 7420 23675
rect 8294 23672 8300 23724
rect 8352 23712 8358 23724
rect 8938 23712 8944 23724
rect 8352 23684 8944 23712
rect 8352 23672 8358 23684
rect 8938 23672 8944 23684
rect 8996 23672 9002 23724
rect 9769 23715 9827 23721
rect 9769 23681 9781 23715
rect 9815 23712 9827 23715
rect 9950 23712 9956 23724
rect 9815 23684 9956 23712
rect 9815 23681 9827 23684
rect 9769 23675 9827 23681
rect 9950 23672 9956 23684
rect 10008 23672 10014 23724
rect 10686 23712 10692 23724
rect 10647 23684 10692 23712
rect 10686 23672 10692 23684
rect 10744 23672 10750 23724
rect 14826 23672 14832 23724
rect 14884 23712 14890 23724
rect 15197 23715 15255 23721
rect 15197 23712 15209 23715
rect 14884 23684 15209 23712
rect 14884 23672 14890 23684
rect 15197 23681 15209 23684
rect 15243 23681 15255 23715
rect 20346 23712 20352 23724
rect 20307 23684 20352 23712
rect 15197 23675 15255 23681
rect 20346 23672 20352 23684
rect 20404 23672 20410 23724
rect 23400 23712 23428 23820
rect 24026 23808 24032 23820
rect 24084 23808 24090 23860
rect 25409 23851 25467 23857
rect 25409 23817 25421 23851
rect 25455 23848 25467 23851
rect 25590 23848 25596 23860
rect 25455 23820 25596 23848
rect 25455 23817 25467 23820
rect 25409 23811 25467 23817
rect 25590 23808 25596 23820
rect 25648 23808 25654 23860
rect 25774 23848 25780 23860
rect 25735 23820 25780 23848
rect 25774 23808 25780 23820
rect 25832 23808 25838 23860
rect 23661 23783 23719 23789
rect 23661 23749 23673 23783
rect 23707 23780 23719 23783
rect 25222 23780 25228 23792
rect 23707 23752 25228 23780
rect 23707 23749 23719 23752
rect 23661 23743 23719 23749
rect 25222 23740 25228 23752
rect 25280 23740 25286 23792
rect 24213 23715 24271 23721
rect 24213 23712 24225 23715
rect 22112 23684 23428 23712
rect 23492 23684 24225 23712
rect 6604 23616 7420 23644
rect 7929 23647 7987 23653
rect 6604 23604 6610 23616
rect 7929 23613 7941 23647
rect 7975 23644 7987 23647
rect 8757 23647 8815 23653
rect 8757 23644 8769 23647
rect 7975 23616 8769 23644
rect 7975 23613 7987 23616
rect 7929 23607 7987 23613
rect 8757 23613 8769 23616
rect 8803 23644 8815 23647
rect 10042 23644 10048 23656
rect 8803 23616 10048 23644
rect 8803 23613 8815 23616
rect 8757 23607 8815 23613
rect 10042 23604 10048 23616
rect 10100 23604 10106 23656
rect 10134 23604 10140 23656
rect 10192 23644 10198 23656
rect 10413 23647 10471 23653
rect 10413 23644 10425 23647
rect 10192 23616 10425 23644
rect 10192 23604 10198 23616
rect 10413 23613 10425 23616
rect 10459 23644 10471 23647
rect 10778 23644 10784 23656
rect 10459 23616 10784 23644
rect 10459 23613 10471 23616
rect 10413 23607 10471 23613
rect 10778 23604 10784 23616
rect 10836 23604 10842 23656
rect 11330 23604 11336 23656
rect 11388 23644 11394 23656
rect 12437 23647 12495 23653
rect 12437 23644 12449 23647
rect 11388 23616 12449 23644
rect 11388 23604 11394 23616
rect 12437 23613 12449 23616
rect 12483 23613 12495 23647
rect 12437 23607 12495 23613
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23644 18107 23647
rect 19242 23644 19248 23656
rect 18095 23616 19248 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 19242 23604 19248 23616
rect 19300 23604 19306 23656
rect 21910 23604 21916 23656
rect 21968 23644 21974 23656
rect 22112 23644 22140 23684
rect 22646 23644 22652 23656
rect 21968 23616 22140 23644
rect 22204 23616 22652 23644
rect 21968 23604 21974 23616
rect 8846 23576 8852 23588
rect 5123 23548 5856 23576
rect 8807 23548 8852 23576
rect 5123 23545 5135 23548
rect 5077 23539 5135 23545
rect 8846 23536 8852 23548
rect 8904 23536 8910 23588
rect 10594 23536 10600 23588
rect 10652 23536 10658 23588
rect 11885 23579 11943 23585
rect 11885 23545 11897 23579
rect 11931 23576 11943 23579
rect 12250 23576 12256 23588
rect 11931 23548 12256 23576
rect 11931 23545 11943 23548
rect 11885 23539 11943 23545
rect 12250 23536 12256 23548
rect 12308 23576 12314 23588
rect 12710 23585 12716 23588
rect 12682 23579 12716 23585
rect 12682 23576 12694 23579
rect 12308 23548 12694 23576
rect 12308 23536 12314 23548
rect 12682 23545 12694 23548
rect 12768 23576 12774 23588
rect 15470 23585 15476 23588
rect 15464 23576 15476 23585
rect 12768 23548 12830 23576
rect 15431 23548 15476 23576
rect 12682 23539 12716 23545
rect 12710 23536 12716 23539
rect 12768 23536 12774 23548
rect 15464 23539 15476 23548
rect 15470 23536 15476 23539
rect 15528 23536 15534 23588
rect 18294 23579 18352 23585
rect 18294 23576 18306 23579
rect 17512 23548 18306 23576
rect 1581 23511 1639 23517
rect 1581 23477 1593 23511
rect 1627 23508 1639 23511
rect 1670 23508 1676 23520
rect 1627 23480 1676 23508
rect 1627 23477 1639 23480
rect 1581 23471 1639 23477
rect 1670 23468 1676 23480
rect 1728 23468 1734 23520
rect 1946 23508 1952 23520
rect 1907 23480 1952 23508
rect 1946 23468 1952 23480
rect 2004 23468 2010 23520
rect 2682 23508 2688 23520
rect 2643 23480 2688 23508
rect 2682 23468 2688 23480
rect 2740 23468 2746 23520
rect 3510 23508 3516 23520
rect 3471 23480 3516 23508
rect 3510 23468 3516 23480
rect 3568 23468 3574 23520
rect 5166 23508 5172 23520
rect 5127 23480 5172 23508
rect 5166 23468 5172 23480
rect 5224 23468 5230 23520
rect 6273 23511 6331 23517
rect 6273 23477 6285 23511
rect 6319 23508 6331 23511
rect 6546 23508 6552 23520
rect 6319 23480 6552 23508
rect 6319 23477 6331 23480
rect 6273 23471 6331 23477
rect 6546 23468 6552 23480
rect 6604 23468 6610 23520
rect 6914 23468 6920 23520
rect 6972 23508 6978 23520
rect 7193 23511 7251 23517
rect 7193 23508 7205 23511
rect 6972 23480 7205 23508
rect 6972 23468 6978 23480
rect 7193 23477 7205 23480
rect 7239 23477 7251 23511
rect 7193 23471 7251 23477
rect 9766 23468 9772 23520
rect 9824 23508 9830 23520
rect 10505 23511 10563 23517
rect 10505 23508 10517 23511
rect 9824 23480 10517 23508
rect 9824 23468 9830 23480
rect 10505 23477 10517 23480
rect 10551 23477 10563 23511
rect 10612 23508 10640 23536
rect 17512 23520 17540 23548
rect 18294 23545 18306 23548
rect 18340 23545 18352 23579
rect 18294 23539 18352 23545
rect 20530 23536 20536 23588
rect 20588 23585 20594 23588
rect 20588 23579 20652 23585
rect 20588 23545 20606 23579
rect 20640 23545 20652 23579
rect 20588 23539 20652 23545
rect 20588 23536 20594 23539
rect 22094 23536 22100 23588
rect 22152 23576 22158 23588
rect 22204 23576 22232 23616
rect 22646 23604 22652 23616
rect 22704 23604 22710 23656
rect 22152 23548 22232 23576
rect 22152 23536 22158 23548
rect 22462 23536 22468 23588
rect 22520 23576 22526 23588
rect 22830 23576 22836 23588
rect 22520 23548 22836 23576
rect 22520 23536 22526 23548
rect 22830 23536 22836 23548
rect 22888 23576 22894 23588
rect 23017 23579 23075 23585
rect 23017 23576 23029 23579
rect 22888 23548 23029 23576
rect 22888 23536 22894 23548
rect 23017 23545 23029 23548
rect 23063 23545 23075 23579
rect 23017 23539 23075 23545
rect 10778 23508 10784 23520
rect 10612 23480 10784 23508
rect 10505 23471 10563 23477
rect 10778 23468 10784 23480
rect 10836 23468 10842 23520
rect 13814 23508 13820 23520
rect 13775 23480 13820 23508
rect 13814 23468 13820 23480
rect 13872 23468 13878 23520
rect 14182 23508 14188 23520
rect 14143 23480 14188 23508
rect 14182 23468 14188 23480
rect 14240 23468 14246 23520
rect 14553 23511 14611 23517
rect 14553 23477 14565 23511
rect 14599 23508 14611 23511
rect 14734 23508 14740 23520
rect 14599 23480 14740 23508
rect 14599 23477 14611 23480
rect 14553 23471 14611 23477
rect 14734 23468 14740 23480
rect 14792 23468 14798 23520
rect 15838 23468 15844 23520
rect 15896 23508 15902 23520
rect 16574 23508 16580 23520
rect 15896 23480 16580 23508
rect 15896 23468 15902 23480
rect 16574 23468 16580 23480
rect 16632 23468 16638 23520
rect 17494 23508 17500 23520
rect 17455 23480 17500 23508
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 19334 23468 19340 23520
rect 19392 23508 19398 23520
rect 19705 23511 19763 23517
rect 19705 23508 19717 23511
rect 19392 23480 19717 23508
rect 19392 23468 19398 23480
rect 19705 23477 19717 23480
rect 19751 23477 19763 23511
rect 19705 23471 19763 23477
rect 20257 23511 20315 23517
rect 20257 23477 20269 23511
rect 20303 23508 20315 23511
rect 20346 23508 20352 23520
rect 20303 23480 20352 23508
rect 20303 23477 20315 23480
rect 20257 23471 20315 23477
rect 20346 23468 20352 23480
rect 20404 23508 20410 23520
rect 20806 23508 20812 23520
rect 20404 23480 20812 23508
rect 20404 23468 20410 23480
rect 20806 23468 20812 23480
rect 20864 23468 20870 23520
rect 21726 23508 21732 23520
rect 21687 23480 21732 23508
rect 21726 23468 21732 23480
rect 21784 23468 21790 23520
rect 22278 23468 22284 23520
rect 22336 23508 22342 23520
rect 22373 23511 22431 23517
rect 22373 23508 22385 23511
rect 22336 23480 22385 23508
rect 22336 23468 22342 23480
rect 22373 23477 22385 23480
rect 22419 23477 22431 23511
rect 22554 23508 22560 23520
rect 22515 23480 22560 23508
rect 22373 23471 22431 23477
rect 22554 23468 22560 23480
rect 22612 23468 22618 23520
rect 23382 23468 23388 23520
rect 23440 23508 23446 23520
rect 23492 23517 23520 23684
rect 24213 23681 24225 23684
rect 24259 23681 24271 23715
rect 24213 23675 24271 23681
rect 25225 23647 25283 23653
rect 25225 23644 25237 23647
rect 25056 23616 25237 23644
rect 24673 23579 24731 23585
rect 24673 23576 24685 23579
rect 24044 23548 24685 23576
rect 24044 23520 24072 23548
rect 24673 23545 24685 23548
rect 24719 23545 24731 23579
rect 24673 23539 24731 23545
rect 23477 23511 23535 23517
rect 23477 23508 23489 23511
rect 23440 23480 23489 23508
rect 23440 23468 23446 23480
rect 23477 23477 23489 23480
rect 23523 23477 23535 23511
rect 24026 23508 24032 23520
rect 23987 23480 24032 23508
rect 23477 23471 23535 23477
rect 24026 23468 24032 23480
rect 24084 23468 24090 23520
rect 24118 23468 24124 23520
rect 24176 23508 24182 23520
rect 24176 23480 24221 23508
rect 24176 23468 24182 23480
rect 24946 23468 24952 23520
rect 25004 23508 25010 23520
rect 25056 23517 25084 23616
rect 25225 23613 25237 23616
rect 25271 23613 25283 23647
rect 25225 23607 25283 23613
rect 25041 23511 25099 23517
rect 25041 23508 25053 23511
rect 25004 23480 25053 23508
rect 25004 23468 25010 23480
rect 25041 23477 25053 23480
rect 25087 23477 25099 23511
rect 25041 23471 25099 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2501 23307 2559 23313
rect 2501 23273 2513 23307
rect 2547 23304 2559 23307
rect 2590 23304 2596 23316
rect 2547 23276 2596 23304
rect 2547 23273 2559 23276
rect 2501 23267 2559 23273
rect 2590 23264 2596 23276
rect 2648 23264 2654 23316
rect 4062 23264 4068 23316
rect 4120 23304 4126 23316
rect 4249 23307 4307 23313
rect 4249 23304 4261 23307
rect 4120 23276 4261 23304
rect 4120 23264 4126 23276
rect 4249 23273 4261 23276
rect 4295 23273 4307 23307
rect 5442 23304 5448 23316
rect 4249 23267 4307 23273
rect 5184 23276 5448 23304
rect 2222 23236 2228 23248
rect 1688 23208 2228 23236
rect 1688 23177 1716 23208
rect 2222 23196 2228 23208
rect 2280 23196 2286 23248
rect 3510 23236 3516 23248
rect 3423 23208 3516 23236
rect 3510 23196 3516 23208
rect 3568 23236 3574 23248
rect 3881 23239 3939 23245
rect 3881 23236 3893 23239
rect 3568 23208 3893 23236
rect 3568 23196 3574 23208
rect 3881 23205 3893 23208
rect 3927 23236 3939 23239
rect 3970 23236 3976 23248
rect 3927 23208 3976 23236
rect 3927 23205 3939 23208
rect 3881 23199 3939 23205
rect 3970 23196 3976 23208
rect 4028 23236 4034 23248
rect 5184 23236 5212 23276
rect 5442 23264 5448 23276
rect 5500 23264 5506 23316
rect 7282 23304 7288 23316
rect 7243 23276 7288 23304
rect 7282 23264 7288 23276
rect 7340 23264 7346 23316
rect 9030 23304 9036 23316
rect 8991 23276 9036 23304
rect 9030 23264 9036 23276
rect 9088 23264 9094 23316
rect 9493 23307 9551 23313
rect 9493 23273 9505 23307
rect 9539 23304 9551 23307
rect 9582 23304 9588 23316
rect 9539 23276 9588 23304
rect 9539 23273 9551 23276
rect 9493 23267 9551 23273
rect 9582 23264 9588 23276
rect 9640 23264 9646 23316
rect 9677 23307 9735 23313
rect 9677 23273 9689 23307
rect 9723 23304 9735 23307
rect 9766 23304 9772 23316
rect 9723 23276 9772 23304
rect 9723 23273 9735 23276
rect 9677 23267 9735 23273
rect 9766 23264 9772 23276
rect 9824 23264 9830 23316
rect 11238 23304 11244 23316
rect 11151 23276 11244 23304
rect 11238 23264 11244 23276
rect 11296 23304 11302 23316
rect 12066 23304 12072 23316
rect 11296 23276 12072 23304
rect 11296 23264 11302 23276
rect 12066 23264 12072 23276
rect 12124 23264 12130 23316
rect 12710 23304 12716 23316
rect 12671 23276 12716 23304
rect 12710 23264 12716 23276
rect 12768 23264 12774 23316
rect 13357 23307 13415 23313
rect 13357 23273 13369 23307
rect 13403 23304 13415 23307
rect 13630 23304 13636 23316
rect 13403 23276 13636 23304
rect 13403 23273 13415 23276
rect 13357 23267 13415 23273
rect 13630 23264 13636 23276
rect 13688 23264 13694 23316
rect 13722 23264 13728 23316
rect 13780 23304 13786 23316
rect 13909 23307 13967 23313
rect 13909 23304 13921 23307
rect 13780 23276 13921 23304
rect 13780 23264 13786 23276
rect 13909 23273 13921 23276
rect 13955 23273 13967 23307
rect 15102 23304 15108 23316
rect 15063 23276 15108 23304
rect 13909 23267 13967 23273
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 15470 23264 15476 23316
rect 15528 23304 15534 23316
rect 15841 23307 15899 23313
rect 15841 23304 15853 23307
rect 15528 23276 15853 23304
rect 15528 23264 15534 23276
rect 15841 23273 15853 23276
rect 15887 23304 15899 23307
rect 16482 23304 16488 23316
rect 15887 23276 16488 23304
rect 15887 23273 15899 23276
rect 15841 23267 15899 23273
rect 16482 23264 16488 23276
rect 16540 23264 16546 23316
rect 17494 23264 17500 23316
rect 17552 23304 17558 23316
rect 17681 23307 17739 23313
rect 17681 23304 17693 23307
rect 17552 23276 17693 23304
rect 17552 23264 17558 23276
rect 17681 23273 17693 23276
rect 17727 23304 17739 23307
rect 18049 23307 18107 23313
rect 18049 23304 18061 23307
rect 17727 23276 18061 23304
rect 17727 23273 17739 23276
rect 17681 23267 17739 23273
rect 18049 23273 18061 23276
rect 18095 23304 18107 23307
rect 18322 23304 18328 23316
rect 18095 23276 18328 23304
rect 18095 23273 18107 23276
rect 18049 23267 18107 23273
rect 18322 23264 18328 23276
rect 18380 23264 18386 23316
rect 18506 23304 18512 23316
rect 18467 23276 18512 23304
rect 18506 23264 18512 23276
rect 18564 23264 18570 23316
rect 19981 23307 20039 23313
rect 19981 23273 19993 23307
rect 20027 23304 20039 23307
rect 20441 23307 20499 23313
rect 20441 23304 20453 23307
rect 20027 23276 20453 23304
rect 20027 23273 20039 23276
rect 19981 23267 20039 23273
rect 20441 23273 20453 23276
rect 20487 23304 20499 23307
rect 20530 23304 20536 23316
rect 20487 23276 20536 23304
rect 20487 23273 20499 23276
rect 20441 23267 20499 23273
rect 20530 23264 20536 23276
rect 20588 23264 20594 23316
rect 22925 23307 22983 23313
rect 22925 23273 22937 23307
rect 22971 23304 22983 23307
rect 23014 23304 23020 23316
rect 22971 23276 23020 23304
rect 22971 23273 22983 23276
rect 22925 23267 22983 23273
rect 23014 23264 23020 23276
rect 23072 23304 23078 23316
rect 23201 23307 23259 23313
rect 23201 23304 23213 23307
rect 23072 23276 23213 23304
rect 23072 23264 23078 23276
rect 23201 23273 23213 23276
rect 23247 23273 23259 23307
rect 23566 23304 23572 23316
rect 23527 23276 23572 23304
rect 23201 23267 23259 23273
rect 23566 23264 23572 23276
rect 23624 23304 23630 23316
rect 24213 23307 24271 23313
rect 24213 23304 24225 23307
rect 23624 23276 24225 23304
rect 23624 23264 23630 23276
rect 24213 23273 24225 23276
rect 24259 23273 24271 23307
rect 24854 23304 24860 23316
rect 24815 23276 24860 23304
rect 24213 23267 24271 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 25498 23304 25504 23316
rect 25459 23276 25504 23304
rect 25498 23264 25504 23276
rect 25556 23264 25562 23316
rect 4028 23208 5212 23236
rect 4028 23196 4034 23208
rect 5184 23177 5212 23208
rect 12434 23196 12440 23248
rect 12492 23236 12498 23248
rect 16114 23236 16120 23248
rect 12492 23208 16120 23236
rect 12492 23196 12498 23208
rect 16114 23196 16120 23208
rect 16172 23196 16178 23248
rect 16574 23245 16580 23248
rect 16568 23236 16580 23245
rect 16535 23208 16580 23236
rect 16568 23199 16580 23208
rect 16574 23196 16580 23199
rect 16632 23196 16638 23248
rect 18690 23196 18696 23248
rect 18748 23236 18754 23248
rect 18846 23239 18904 23245
rect 18846 23236 18858 23239
rect 18748 23208 18858 23236
rect 18748 23196 18754 23208
rect 18846 23205 18858 23208
rect 18892 23205 18904 23239
rect 18846 23199 18904 23205
rect 21726 23196 21732 23248
rect 21784 23245 21790 23248
rect 21784 23239 21848 23245
rect 21784 23205 21802 23239
rect 21836 23205 21848 23239
rect 21784 23199 21848 23205
rect 21784 23196 21790 23199
rect 1673 23171 1731 23177
rect 1673 23137 1685 23171
rect 1719 23137 1731 23171
rect 1673 23131 1731 23137
rect 1949 23171 2007 23177
rect 1949 23137 1961 23171
rect 1995 23168 2007 23171
rect 4065 23171 4123 23177
rect 4065 23168 4077 23171
rect 1995 23140 4077 23168
rect 1995 23137 2007 23140
rect 1949 23131 2007 23137
rect 4065 23137 4077 23140
rect 4111 23168 4123 23171
rect 4617 23171 4675 23177
rect 4617 23168 4629 23171
rect 4111 23140 4629 23168
rect 4111 23137 4123 23140
rect 4065 23131 4123 23137
rect 4617 23137 4629 23140
rect 4663 23137 4675 23171
rect 4617 23131 4675 23137
rect 5169 23171 5227 23177
rect 5169 23137 5181 23171
rect 5215 23137 5227 23171
rect 5169 23131 5227 23137
rect 5436 23171 5494 23177
rect 5436 23137 5448 23171
rect 5482 23168 5494 23171
rect 6178 23168 6184 23180
rect 5482 23140 6184 23168
rect 5482 23137 5494 23140
rect 5436 23131 5494 23137
rect 6178 23128 6184 23140
rect 6236 23128 6242 23180
rect 7650 23177 7656 23180
rect 7644 23168 7656 23177
rect 7611 23140 7656 23168
rect 7644 23131 7656 23140
rect 7650 23128 7656 23131
rect 7708 23128 7714 23180
rect 10042 23168 10048 23180
rect 10003 23140 10048 23168
rect 10042 23128 10048 23140
rect 10100 23128 10106 23180
rect 11606 23177 11612 23180
rect 11600 23168 11612 23177
rect 11567 23140 11612 23168
rect 11600 23131 11612 23140
rect 11606 23128 11612 23131
rect 11664 23128 11670 23180
rect 12618 23128 12624 23180
rect 12676 23168 12682 23180
rect 14001 23171 14059 23177
rect 14001 23168 14013 23171
rect 12676 23140 14013 23168
rect 12676 23128 12682 23140
rect 14001 23137 14013 23140
rect 14047 23137 14059 23171
rect 14001 23131 14059 23137
rect 15930 23128 15936 23180
rect 15988 23168 15994 23180
rect 16301 23171 16359 23177
rect 16301 23168 16313 23171
rect 15988 23140 16313 23168
rect 15988 23128 15994 23140
rect 16301 23137 16313 23140
rect 16347 23168 16359 23171
rect 16390 23168 16396 23180
rect 16347 23140 16396 23168
rect 16347 23137 16359 23140
rect 16301 23131 16359 23137
rect 16390 23128 16396 23140
rect 16448 23128 16454 23180
rect 18601 23171 18659 23177
rect 18601 23137 18613 23171
rect 18647 23168 18659 23171
rect 19242 23168 19248 23180
rect 18647 23140 19248 23168
rect 18647 23137 18659 23140
rect 18601 23131 18659 23137
rect 19242 23128 19248 23140
rect 19300 23128 19306 23180
rect 21545 23171 21603 23177
rect 21545 23137 21557 23171
rect 21591 23168 21603 23171
rect 21634 23168 21640 23180
rect 21591 23140 21640 23168
rect 21591 23137 21603 23140
rect 21545 23131 21603 23137
rect 21634 23128 21640 23140
rect 21692 23128 21698 23180
rect 23842 23128 23848 23180
rect 23900 23168 23906 23180
rect 24121 23171 24179 23177
rect 24121 23168 24133 23171
rect 23900 23140 24133 23168
rect 23900 23128 23906 23140
rect 24121 23137 24133 23140
rect 24167 23137 24179 23171
rect 25314 23168 25320 23180
rect 25275 23140 25320 23168
rect 24121 23131 24179 23137
rect 25314 23128 25320 23140
rect 25372 23128 25378 23180
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23100 3019 23103
rect 4982 23100 4988 23112
rect 3007 23072 4988 23100
rect 3007 23069 3019 23072
rect 2961 23063 3019 23069
rect 4982 23060 4988 23072
rect 5040 23060 5046 23112
rect 7374 23100 7380 23112
rect 7335 23072 7380 23100
rect 7374 23060 7380 23072
rect 7432 23060 7438 23112
rect 9490 23060 9496 23112
rect 9548 23100 9554 23112
rect 10137 23103 10195 23109
rect 10137 23100 10149 23103
rect 9548 23072 10149 23100
rect 9548 23060 9554 23072
rect 10137 23069 10149 23072
rect 10183 23069 10195 23103
rect 10137 23063 10195 23069
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23069 10287 23103
rect 10229 23063 10287 23069
rect 2869 23035 2927 23041
rect 2869 23001 2881 23035
rect 2915 23032 2927 23035
rect 3878 23032 3884 23044
rect 2915 23004 3884 23032
rect 2915 23001 2927 23004
rect 2869 22995 2927 23001
rect 3878 22992 3884 23004
rect 3936 22992 3942 23044
rect 9766 22992 9772 23044
rect 9824 23032 9830 23044
rect 10244 23032 10272 23063
rect 10594 23060 10600 23112
rect 10652 23100 10658 23112
rect 10778 23100 10784 23112
rect 10652 23072 10784 23100
rect 10652 23060 10658 23072
rect 10778 23060 10784 23072
rect 10836 23060 10842 23112
rect 11330 23100 11336 23112
rect 11291 23072 11336 23100
rect 11330 23060 11336 23072
rect 11388 23060 11394 23112
rect 12526 23060 12532 23112
rect 12584 23100 12590 23112
rect 13630 23100 13636 23112
rect 12584 23072 13636 23100
rect 12584 23060 12590 23072
rect 13630 23060 13636 23072
rect 13688 23060 13694 23112
rect 14090 23060 14096 23112
rect 14148 23100 14154 23112
rect 15286 23100 15292 23112
rect 14148 23072 14193 23100
rect 15247 23072 15292 23100
rect 14148 23060 14154 23072
rect 15286 23060 15292 23072
rect 15344 23060 15350 23112
rect 23934 23060 23940 23112
rect 23992 23100 23998 23112
rect 24305 23103 24363 23109
rect 24305 23100 24317 23103
rect 23992 23072 24317 23100
rect 23992 23060 23998 23072
rect 24305 23069 24317 23072
rect 24351 23069 24363 23103
rect 24305 23063 24363 23069
rect 9824 23004 10272 23032
rect 9824 22992 9830 23004
rect 23474 22992 23480 23044
rect 23532 23032 23538 23044
rect 23753 23035 23811 23041
rect 23753 23032 23765 23035
rect 23532 23004 23765 23032
rect 23532 22992 23538 23004
rect 23753 23001 23765 23004
rect 23799 23001 23811 23035
rect 23753 22995 23811 23001
rect 5074 22964 5080 22976
rect 5035 22936 5080 22964
rect 5074 22924 5080 22936
rect 5132 22924 5138 22976
rect 6546 22964 6552 22976
rect 6507 22936 6552 22964
rect 6546 22924 6552 22936
rect 6604 22924 6610 22976
rect 6917 22967 6975 22973
rect 6917 22933 6929 22967
rect 6963 22964 6975 22967
rect 7190 22964 7196 22976
rect 6963 22936 7196 22964
rect 6963 22933 6975 22936
rect 6917 22927 6975 22933
rect 7190 22924 7196 22936
rect 7248 22924 7254 22976
rect 8386 22924 8392 22976
rect 8444 22964 8450 22976
rect 8757 22967 8815 22973
rect 8757 22964 8769 22967
rect 8444 22936 8769 22964
rect 8444 22924 8450 22936
rect 8757 22933 8769 22936
rect 8803 22933 8815 22967
rect 10778 22964 10784 22976
rect 10739 22936 10784 22964
rect 8757 22927 8815 22933
rect 10778 22924 10784 22936
rect 10836 22924 10842 22976
rect 12802 22924 12808 22976
rect 12860 22964 12866 22976
rect 13541 22967 13599 22973
rect 13541 22964 13553 22967
rect 12860 22936 13553 22964
rect 12860 22924 12866 22936
rect 13541 22933 13553 22936
rect 13587 22933 13599 22967
rect 13541 22927 13599 22933
rect 14366 22924 14372 22976
rect 14424 22964 14430 22976
rect 14553 22967 14611 22973
rect 14553 22964 14565 22967
rect 14424 22936 14565 22964
rect 14424 22924 14430 22936
rect 14553 22933 14565 22936
rect 14599 22933 14611 22967
rect 14553 22927 14611 22933
rect 16209 22967 16267 22973
rect 16209 22933 16221 22967
rect 16255 22964 16267 22967
rect 16666 22964 16672 22976
rect 16255 22936 16672 22964
rect 16255 22933 16267 22936
rect 16209 22927 16267 22933
rect 16666 22924 16672 22936
rect 16724 22924 16730 22976
rect 21082 22964 21088 22976
rect 21043 22936 21088 22964
rect 21082 22924 21088 22936
rect 21140 22924 21146 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2222 22760 2228 22772
rect 2183 22732 2228 22760
rect 2222 22720 2228 22732
rect 2280 22720 2286 22772
rect 4890 22720 4896 22772
rect 4948 22760 4954 22772
rect 5169 22763 5227 22769
rect 5169 22760 5181 22763
rect 4948 22732 5181 22760
rect 4948 22720 4954 22732
rect 5169 22729 5181 22732
rect 5215 22729 5227 22763
rect 5169 22723 5227 22729
rect 7006 22720 7012 22772
rect 7064 22760 7070 22772
rect 7837 22763 7895 22769
rect 7837 22760 7849 22763
rect 7064 22732 7849 22760
rect 7064 22720 7070 22732
rect 7837 22729 7849 22732
rect 7883 22760 7895 22763
rect 7883 22732 8892 22760
rect 7883 22729 7895 22732
rect 7837 22723 7895 22729
rect 4982 22692 4988 22704
rect 4943 22664 4988 22692
rect 4982 22652 4988 22664
rect 5040 22652 5046 22704
rect 6825 22695 6883 22701
rect 6825 22692 6837 22695
rect 5644 22664 6837 22692
rect 2590 22624 2596 22636
rect 1412 22596 2596 22624
rect 1412 22565 1440 22596
rect 2590 22584 2596 22596
rect 2648 22584 2654 22636
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22525 1455 22559
rect 1397 22519 1455 22525
rect 1673 22559 1731 22565
rect 1673 22525 1685 22559
rect 1719 22556 1731 22559
rect 2130 22556 2136 22568
rect 1719 22528 2136 22556
rect 1719 22525 1731 22528
rect 1673 22519 1731 22525
rect 2130 22516 2136 22528
rect 2188 22516 2194 22568
rect 2685 22559 2743 22565
rect 2685 22525 2697 22559
rect 2731 22556 2743 22559
rect 3970 22556 3976 22568
rect 2731 22528 3976 22556
rect 2731 22525 2743 22528
rect 2685 22519 2743 22525
rect 3970 22516 3976 22528
rect 4028 22516 4034 22568
rect 5000 22556 5028 22652
rect 5074 22584 5080 22636
rect 5132 22624 5138 22636
rect 5644 22633 5672 22664
rect 6825 22661 6837 22664
rect 6871 22661 6883 22695
rect 6825 22655 6883 22661
rect 8864 22692 8892 22732
rect 8938 22720 8944 22772
rect 8996 22760 9002 22772
rect 9490 22760 9496 22772
rect 8996 22732 9496 22760
rect 8996 22720 9002 22732
rect 9490 22720 9496 22732
rect 9548 22720 9554 22772
rect 9861 22763 9919 22769
rect 9861 22760 9873 22763
rect 9600 22732 9873 22760
rect 9600 22692 9628 22732
rect 9861 22729 9873 22732
rect 9907 22729 9919 22763
rect 9861 22723 9919 22729
rect 10321 22763 10379 22769
rect 10321 22729 10333 22763
rect 10367 22760 10379 22763
rect 10962 22760 10968 22772
rect 10367 22732 10968 22760
rect 10367 22729 10379 22732
rect 10321 22723 10379 22729
rect 10962 22720 10968 22732
rect 11020 22720 11026 22772
rect 12710 22720 12716 22772
rect 12768 22760 12774 22772
rect 13541 22763 13599 22769
rect 13541 22760 13553 22763
rect 12768 22732 13553 22760
rect 12768 22720 12774 22732
rect 13541 22729 13553 22732
rect 13587 22760 13599 22763
rect 14090 22760 14096 22772
rect 13587 22732 14096 22760
rect 13587 22729 13599 22732
rect 13541 22723 13599 22729
rect 14090 22720 14096 22732
rect 14148 22720 14154 22772
rect 15838 22760 15844 22772
rect 15799 22732 15844 22760
rect 15838 22720 15844 22732
rect 15896 22720 15902 22772
rect 18046 22760 18052 22772
rect 18007 22732 18052 22760
rect 18046 22720 18052 22732
rect 18104 22720 18110 22772
rect 18690 22720 18696 22772
rect 18748 22760 18754 22772
rect 19061 22763 19119 22769
rect 19061 22760 19073 22763
rect 18748 22732 19073 22760
rect 18748 22720 18754 22732
rect 19061 22729 19073 22732
rect 19107 22729 19119 22763
rect 19061 22723 19119 22729
rect 19889 22763 19947 22769
rect 19889 22729 19901 22763
rect 19935 22760 19947 22763
rect 19978 22760 19984 22772
rect 19935 22732 19984 22760
rect 19935 22729 19947 22732
rect 19889 22723 19947 22729
rect 19978 22720 19984 22732
rect 20036 22720 20042 22772
rect 20349 22763 20407 22769
rect 20349 22729 20361 22763
rect 20395 22760 20407 22763
rect 20622 22760 20628 22772
rect 20395 22732 20628 22760
rect 20395 22729 20407 22732
rect 20349 22723 20407 22729
rect 20622 22720 20628 22732
rect 20680 22720 20686 22772
rect 21545 22763 21603 22769
rect 21545 22729 21557 22763
rect 21591 22760 21603 22763
rect 21726 22760 21732 22772
rect 21591 22732 21732 22760
rect 21591 22729 21603 22732
rect 21545 22723 21603 22729
rect 8864 22664 9628 22692
rect 5629 22627 5687 22633
rect 5629 22624 5641 22627
rect 5132 22596 5641 22624
rect 5132 22584 5138 22596
rect 5629 22593 5641 22596
rect 5675 22593 5687 22627
rect 5810 22624 5816 22636
rect 5771 22596 5816 22624
rect 5629 22587 5687 22593
rect 5810 22584 5816 22596
rect 5868 22624 5874 22636
rect 6546 22624 6552 22636
rect 5868 22596 6552 22624
rect 5868 22584 5874 22596
rect 6546 22584 6552 22596
rect 6604 22584 6610 22636
rect 7466 22624 7472 22636
rect 7379 22596 7472 22624
rect 7466 22584 7472 22596
rect 7524 22624 7530 22636
rect 8202 22624 8208 22636
rect 7524 22596 8208 22624
rect 7524 22584 7530 22596
rect 8202 22584 8208 22596
rect 8260 22584 8266 22636
rect 8864 22633 8892 22664
rect 8849 22627 8907 22633
rect 8849 22593 8861 22627
rect 8895 22593 8907 22627
rect 9030 22624 9036 22636
rect 8991 22596 9036 22624
rect 8849 22587 8907 22593
rect 9030 22584 9036 22596
rect 9088 22584 9094 22636
rect 9600 22624 9628 22664
rect 9766 22652 9772 22704
rect 9824 22692 9830 22704
rect 11333 22695 11391 22701
rect 11333 22692 11345 22695
rect 9824 22664 11345 22692
rect 9824 22652 9830 22664
rect 11333 22661 11345 22664
rect 11379 22661 11391 22695
rect 11333 22655 11391 22661
rect 12176 22664 13124 22692
rect 10781 22627 10839 22633
rect 10781 22624 10793 22627
rect 9600 22596 10793 22624
rect 10781 22593 10793 22596
rect 10827 22593 10839 22627
rect 10781 22587 10839 22593
rect 10873 22627 10931 22633
rect 10873 22593 10885 22627
rect 10919 22624 10931 22627
rect 11606 22624 11612 22636
rect 10919 22596 11612 22624
rect 10919 22593 10931 22596
rect 10873 22587 10931 22593
rect 5537 22559 5595 22565
rect 5537 22556 5549 22559
rect 5000 22528 5549 22556
rect 5537 22525 5549 22528
rect 5583 22525 5595 22559
rect 5537 22519 5595 22525
rect 6178 22516 6184 22568
rect 6236 22556 6242 22568
rect 6273 22559 6331 22565
rect 6273 22556 6285 22559
rect 6236 22528 6285 22556
rect 6236 22516 6242 22528
rect 6273 22525 6285 22528
rect 6319 22556 6331 22559
rect 7484 22556 7512 22584
rect 6319 22528 7512 22556
rect 8297 22559 8355 22565
rect 6319 22525 6331 22528
rect 6273 22519 6331 22525
rect 8297 22525 8309 22559
rect 8343 22556 8355 22559
rect 8757 22559 8815 22565
rect 8757 22556 8769 22559
rect 8343 22528 8769 22556
rect 8343 22525 8355 22528
rect 8297 22519 8355 22525
rect 8757 22525 8769 22528
rect 8803 22556 8815 22559
rect 10229 22559 10287 22565
rect 10229 22556 10241 22559
rect 8803 22528 10241 22556
rect 8803 22525 8815 22528
rect 8757 22519 8815 22525
rect 10229 22525 10241 22528
rect 10275 22556 10287 22559
rect 10594 22556 10600 22568
rect 10275 22528 10600 22556
rect 10275 22525 10287 22528
rect 10229 22519 10287 22525
rect 10594 22516 10600 22528
rect 10652 22556 10658 22568
rect 10689 22559 10747 22565
rect 10689 22556 10701 22559
rect 10652 22528 10701 22556
rect 10652 22516 10658 22528
rect 10689 22525 10701 22528
rect 10735 22525 10747 22559
rect 10888 22556 10916 22587
rect 11606 22584 11612 22596
rect 11664 22624 11670 22636
rect 11701 22627 11759 22633
rect 11701 22624 11713 22627
rect 11664 22596 11713 22624
rect 11664 22584 11670 22596
rect 11701 22593 11713 22596
rect 11747 22593 11759 22627
rect 11701 22587 11759 22593
rect 10689 22519 10747 22525
rect 10796 22528 10916 22556
rect 2593 22491 2651 22497
rect 2593 22457 2605 22491
rect 2639 22488 2651 22491
rect 2952 22491 3010 22497
rect 2952 22488 2964 22491
rect 2639 22460 2964 22488
rect 2639 22457 2651 22460
rect 2593 22451 2651 22457
rect 2952 22457 2964 22460
rect 2998 22488 3010 22491
rect 4154 22488 4160 22500
rect 2998 22460 4160 22488
rect 2998 22457 3010 22460
rect 2952 22451 3010 22457
rect 4154 22448 4160 22460
rect 4212 22448 4218 22500
rect 4709 22491 4767 22497
rect 4709 22457 4721 22491
rect 4755 22488 4767 22491
rect 6196 22488 6224 22516
rect 10796 22500 10824 22528
rect 11330 22516 11336 22568
rect 11388 22556 11394 22568
rect 12176 22565 12204 22664
rect 12434 22584 12440 22636
rect 12492 22624 12498 22636
rect 13096 22633 13124 22664
rect 15654 22652 15660 22704
rect 15712 22692 15718 22704
rect 16390 22692 16396 22704
rect 15712 22664 16396 22692
rect 15712 22652 15718 22664
rect 16390 22652 16396 22664
rect 16448 22652 16454 22704
rect 12897 22627 12955 22633
rect 12897 22624 12909 22627
rect 12492 22596 12909 22624
rect 12492 22584 12498 22596
rect 12897 22593 12909 22596
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 13081 22627 13139 22633
rect 13081 22593 13093 22627
rect 13127 22624 13139 22627
rect 13814 22624 13820 22636
rect 13127 22596 13820 22624
rect 13127 22593 13139 22596
rect 13081 22587 13139 22593
rect 13814 22584 13820 22596
rect 13872 22584 13878 22636
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 16132 22596 16865 22624
rect 12161 22559 12219 22565
rect 12161 22556 12173 22559
rect 11388 22528 12173 22556
rect 11388 22516 11394 22528
rect 12161 22525 12173 22528
rect 12207 22525 12219 22559
rect 12161 22519 12219 22525
rect 12526 22516 12532 22568
rect 12584 22556 12590 22568
rect 12802 22556 12808 22568
rect 12584 22528 12808 22556
rect 12584 22516 12590 22528
rect 12802 22516 12808 22528
rect 12860 22516 12866 22568
rect 14090 22556 14096 22568
rect 14051 22528 14096 22556
rect 14090 22516 14096 22528
rect 14148 22516 14154 22568
rect 4755 22460 6224 22488
rect 6641 22491 6699 22497
rect 4755 22457 4767 22460
rect 4709 22451 4767 22457
rect 6641 22457 6653 22491
rect 6687 22488 6699 22491
rect 7282 22488 7288 22500
rect 6687 22460 7288 22488
rect 6687 22457 6699 22460
rect 6641 22451 6699 22457
rect 4062 22420 4068 22432
rect 4023 22392 4068 22420
rect 4062 22380 4068 22392
rect 4120 22380 4126 22432
rect 5350 22380 5356 22432
rect 5408 22420 5414 22432
rect 6656 22420 6684 22451
rect 7282 22448 7288 22460
rect 7340 22448 7346 22500
rect 10778 22448 10784 22500
rect 10836 22448 10842 22500
rect 13446 22448 13452 22500
rect 13504 22488 13510 22500
rect 13814 22488 13820 22500
rect 13504 22460 13820 22488
rect 13504 22448 13510 22460
rect 13814 22448 13820 22460
rect 13872 22448 13878 22500
rect 14001 22491 14059 22497
rect 14001 22457 14013 22491
rect 14047 22488 14059 22491
rect 14338 22491 14396 22497
rect 14338 22488 14350 22491
rect 14047 22460 14350 22488
rect 14047 22457 14059 22460
rect 14001 22451 14059 22457
rect 14338 22457 14350 22460
rect 14384 22488 14396 22491
rect 15378 22488 15384 22500
rect 14384 22460 15384 22488
rect 14384 22457 14396 22460
rect 14338 22451 14396 22457
rect 15378 22448 15384 22460
rect 15436 22448 15442 22500
rect 7190 22420 7196 22432
rect 5408 22392 6684 22420
rect 7151 22392 7196 22420
rect 5408 22380 5414 22392
rect 7190 22380 7196 22392
rect 7248 22380 7254 22432
rect 8386 22420 8392 22432
rect 8347 22392 8392 22420
rect 8386 22380 8392 22392
rect 8444 22380 8450 22432
rect 12434 22380 12440 22432
rect 12492 22420 12498 22432
rect 12492 22392 12537 22420
rect 12492 22380 12498 22392
rect 14734 22380 14740 22432
rect 14792 22420 14798 22432
rect 15473 22423 15531 22429
rect 15473 22420 15485 22423
rect 14792 22392 15485 22420
rect 14792 22380 14798 22392
rect 15473 22389 15485 22392
rect 15519 22389 15531 22423
rect 15473 22383 15531 22389
rect 15838 22380 15844 22432
rect 15896 22420 15902 22432
rect 16132 22429 16160 22596
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 18322 22584 18328 22636
rect 18380 22624 18386 22636
rect 18601 22627 18659 22633
rect 18601 22624 18613 22627
rect 18380 22596 18613 22624
rect 18380 22584 18386 22596
rect 18601 22593 18613 22596
rect 18647 22593 18659 22627
rect 18601 22587 18659 22593
rect 18874 22584 18880 22636
rect 18932 22624 18938 22636
rect 19242 22624 19248 22636
rect 18932 22596 19248 22624
rect 18932 22584 18938 22596
rect 19242 22584 19248 22596
rect 19300 22584 19306 22636
rect 20257 22627 20315 22633
rect 20257 22593 20269 22627
rect 20303 22624 20315 22627
rect 20993 22627 21051 22633
rect 20993 22624 21005 22627
rect 20303 22596 21005 22624
rect 20303 22593 20315 22596
rect 20257 22587 20315 22593
rect 20993 22593 21005 22596
rect 21039 22624 21051 22627
rect 21560 22624 21588 22723
rect 21726 22720 21732 22732
rect 21784 22720 21790 22772
rect 22002 22760 22008 22772
rect 21963 22732 22008 22760
rect 22002 22720 22008 22732
rect 22060 22720 22066 22772
rect 22554 22720 22560 22772
rect 22612 22760 22618 22772
rect 23017 22763 23075 22769
rect 23017 22760 23029 22763
rect 22612 22732 23029 22760
rect 22612 22720 22618 22732
rect 23017 22729 23029 22732
rect 23063 22729 23075 22763
rect 23017 22723 23075 22729
rect 21818 22652 21824 22704
rect 21876 22692 21882 22704
rect 21913 22695 21971 22701
rect 21913 22692 21925 22695
rect 21876 22664 21925 22692
rect 21876 22652 21882 22664
rect 21913 22661 21925 22664
rect 21959 22692 21971 22695
rect 21959 22664 22508 22692
rect 21959 22661 21971 22664
rect 21913 22655 21971 22661
rect 21039 22596 21588 22624
rect 21039 22593 21051 22596
rect 20993 22587 21051 22593
rect 17865 22559 17923 22565
rect 17865 22525 17877 22559
rect 17911 22556 17923 22559
rect 18509 22559 18567 22565
rect 18509 22556 18521 22559
rect 17911 22528 18521 22556
rect 17911 22525 17923 22528
rect 17865 22519 17923 22525
rect 18509 22525 18521 22528
rect 18555 22556 18567 22559
rect 18892 22556 18920 22584
rect 18555 22528 18920 22556
rect 18555 22525 18567 22528
rect 18509 22519 18567 22525
rect 19978 22516 19984 22568
rect 20036 22556 20042 22568
rect 20809 22559 20867 22565
rect 20809 22556 20821 22559
rect 20036 22528 20821 22556
rect 20036 22516 20042 22528
rect 20809 22525 20821 22528
rect 20855 22525 20867 22559
rect 20809 22519 20867 22525
rect 21082 22516 21088 22568
rect 21140 22556 21146 22568
rect 21726 22556 21732 22568
rect 21140 22528 21732 22556
rect 21140 22516 21146 22528
rect 21726 22516 21732 22528
rect 21784 22516 21790 22568
rect 22186 22516 22192 22568
rect 22244 22556 22250 22568
rect 22480 22565 22508 22664
rect 22649 22627 22707 22633
rect 22649 22593 22661 22627
rect 22695 22624 22707 22627
rect 22922 22624 22928 22636
rect 22695 22596 22928 22624
rect 22695 22593 22707 22596
rect 22649 22587 22707 22593
rect 22922 22584 22928 22596
rect 22980 22584 22986 22636
rect 22373 22559 22431 22565
rect 22373 22556 22385 22559
rect 22244 22528 22385 22556
rect 22244 22516 22250 22528
rect 22373 22525 22385 22528
rect 22419 22525 22431 22559
rect 22373 22519 22431 22525
rect 22465 22559 22523 22565
rect 22465 22525 22477 22559
rect 22511 22556 22523 22559
rect 22554 22556 22560 22568
rect 22511 22528 22560 22556
rect 22511 22525 22523 22528
rect 22465 22519 22523 22525
rect 22554 22516 22560 22528
rect 22612 22516 22618 22568
rect 23032 22556 23060 22723
rect 25314 22720 25320 22772
rect 25372 22760 25378 22772
rect 26053 22763 26111 22769
rect 26053 22760 26065 22763
rect 25372 22732 26065 22760
rect 25372 22720 25378 22732
rect 26053 22729 26065 22732
rect 26099 22729 26111 22763
rect 26053 22723 26111 22729
rect 24302 22624 24308 22636
rect 24263 22596 24308 22624
rect 24302 22584 24308 22596
rect 24360 22584 24366 22636
rect 24121 22559 24179 22565
rect 24121 22556 24133 22559
rect 23032 22528 24133 22556
rect 24121 22525 24133 22528
rect 24167 22525 24179 22559
rect 25317 22559 25375 22565
rect 25317 22556 25329 22559
rect 24121 22519 24179 22525
rect 25148 22528 25329 22556
rect 16761 22491 16819 22497
rect 16761 22457 16773 22491
rect 16807 22488 16819 22491
rect 17402 22488 17408 22500
rect 16807 22460 17408 22488
rect 16807 22457 16819 22460
rect 16761 22451 16819 22457
rect 17402 22448 17408 22460
rect 17460 22448 17466 22500
rect 19521 22491 19579 22497
rect 19521 22457 19533 22491
rect 19567 22488 19579 22491
rect 20717 22491 20775 22497
rect 20717 22488 20729 22491
rect 19567 22460 20729 22488
rect 19567 22457 19579 22460
rect 19521 22451 19579 22457
rect 20717 22457 20729 22460
rect 20763 22488 20775 22491
rect 20898 22488 20904 22500
rect 20763 22460 20904 22488
rect 20763 22457 20775 22460
rect 20717 22451 20775 22457
rect 20898 22448 20904 22460
rect 20956 22448 20962 22500
rect 23400 22460 23888 22488
rect 16117 22423 16175 22429
rect 16117 22420 16129 22423
rect 15896 22392 16129 22420
rect 15896 22380 15902 22392
rect 16117 22389 16129 22392
rect 16163 22389 16175 22423
rect 16117 22383 16175 22389
rect 16301 22423 16359 22429
rect 16301 22389 16313 22423
rect 16347 22420 16359 22423
rect 16482 22420 16488 22432
rect 16347 22392 16488 22420
rect 16347 22389 16359 22392
rect 16301 22383 16359 22389
rect 16482 22380 16488 22392
rect 16540 22380 16546 22432
rect 16666 22420 16672 22432
rect 16627 22392 16672 22420
rect 16666 22380 16672 22392
rect 16724 22380 16730 22432
rect 18046 22380 18052 22432
rect 18104 22420 18110 22432
rect 18417 22423 18475 22429
rect 18417 22420 18429 22423
rect 18104 22392 18429 22420
rect 18104 22380 18110 22392
rect 18417 22389 18429 22392
rect 18463 22389 18475 22423
rect 18417 22383 18475 22389
rect 22646 22380 22652 22432
rect 22704 22420 22710 22432
rect 23400 22429 23428 22460
rect 23385 22423 23443 22429
rect 23385 22420 23397 22423
rect 22704 22392 23397 22420
rect 22704 22380 22710 22392
rect 23385 22389 23397 22392
rect 23431 22389 23443 22423
rect 23385 22383 23443 22389
rect 23658 22380 23664 22432
rect 23716 22420 23722 22432
rect 23753 22423 23811 22429
rect 23753 22420 23765 22423
rect 23716 22392 23765 22420
rect 23716 22380 23722 22392
rect 23753 22389 23765 22392
rect 23799 22389 23811 22423
rect 23860 22420 23888 22460
rect 23934 22448 23940 22500
rect 23992 22488 23998 22500
rect 24765 22491 24823 22497
rect 24765 22488 24777 22491
rect 23992 22460 24777 22488
rect 23992 22448 23998 22460
rect 24765 22457 24777 22460
rect 24811 22457 24823 22491
rect 24765 22451 24823 22457
rect 25148 22432 25176 22528
rect 25317 22525 25329 22528
rect 25363 22525 25375 22559
rect 25317 22519 25375 22525
rect 25222 22448 25228 22500
rect 25280 22488 25286 22500
rect 25593 22491 25651 22497
rect 25593 22488 25605 22491
rect 25280 22460 25605 22488
rect 25280 22448 25286 22460
rect 25593 22457 25605 22460
rect 25639 22457 25651 22491
rect 25593 22451 25651 22457
rect 24213 22423 24271 22429
rect 24213 22420 24225 22423
rect 23860 22392 24225 22420
rect 23753 22383 23811 22389
rect 24213 22389 24225 22392
rect 24259 22420 24271 22423
rect 24946 22420 24952 22432
rect 24259 22392 24952 22420
rect 24259 22389 24271 22392
rect 24213 22383 24271 22389
rect 24946 22380 24952 22392
rect 25004 22380 25010 22432
rect 25130 22420 25136 22432
rect 25091 22392 25136 22420
rect 25130 22380 25136 22392
rect 25188 22380 25194 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 2774 22176 2780 22228
rect 2832 22216 2838 22228
rect 5445 22219 5503 22225
rect 2832 22188 2877 22216
rect 2832 22176 2838 22188
rect 5445 22185 5457 22219
rect 5491 22185 5503 22219
rect 5810 22216 5816 22228
rect 5771 22188 5816 22216
rect 5445 22179 5503 22185
rect 4062 22108 4068 22160
rect 4120 22108 4126 22160
rect 5460 22148 5488 22179
rect 5810 22176 5816 22188
rect 5868 22176 5874 22228
rect 7009 22219 7067 22225
rect 7009 22185 7021 22219
rect 7055 22216 7067 22219
rect 7098 22216 7104 22228
rect 7055 22188 7104 22216
rect 7055 22185 7067 22188
rect 7009 22179 7067 22185
rect 7098 22176 7104 22188
rect 7156 22176 7162 22228
rect 7650 22216 7656 22228
rect 7611 22188 7656 22216
rect 7650 22176 7656 22188
rect 7708 22176 7714 22228
rect 10778 22176 10784 22228
rect 10836 22216 10842 22228
rect 11790 22216 11796 22228
rect 10836 22188 11796 22216
rect 10836 22176 10842 22188
rect 11790 22176 11796 22188
rect 11848 22176 11854 22228
rect 13262 22216 13268 22228
rect 12912 22188 13268 22216
rect 12912 22160 12940 22188
rect 13262 22176 13268 22188
rect 13320 22176 13326 22228
rect 13814 22216 13820 22228
rect 13372 22188 13820 22216
rect 6178 22148 6184 22160
rect 5460 22120 6184 22148
rect 6178 22108 6184 22120
rect 6236 22108 6242 22160
rect 11330 22157 11336 22160
rect 11324 22148 11336 22157
rect 11291 22120 11336 22148
rect 11324 22111 11336 22120
rect 11330 22108 11336 22111
rect 11388 22108 11394 22160
rect 12894 22108 12900 22160
rect 12952 22108 12958 22160
rect 13078 22108 13084 22160
rect 13136 22148 13142 22160
rect 13372 22148 13400 22188
rect 13814 22176 13820 22188
rect 13872 22176 13878 22228
rect 18046 22216 18052 22228
rect 18007 22188 18052 22216
rect 18046 22176 18052 22188
rect 18104 22176 18110 22228
rect 18322 22176 18328 22228
rect 18380 22216 18386 22228
rect 18417 22219 18475 22225
rect 18417 22216 18429 22219
rect 18380 22188 18429 22216
rect 18380 22176 18386 22188
rect 18417 22185 18429 22188
rect 18463 22185 18475 22219
rect 18417 22179 18475 22185
rect 13538 22148 13544 22160
rect 13136 22120 13400 22148
rect 13464 22120 13544 22148
rect 13136 22108 13142 22120
rect 4080 22080 4108 22108
rect 4321 22083 4379 22089
rect 4321 22080 4333 22083
rect 4080 22052 4333 22080
rect 4321 22049 4333 22052
rect 4367 22049 4379 22083
rect 4321 22043 4379 22049
rect 8297 22083 8355 22089
rect 8297 22049 8309 22083
rect 8343 22080 8355 22083
rect 9122 22080 9128 22092
rect 8343 22052 9128 22080
rect 8343 22049 8355 22052
rect 8297 22043 8355 22049
rect 9122 22040 9128 22052
rect 9180 22040 9186 22092
rect 9582 22040 9588 22092
rect 9640 22080 9646 22092
rect 9677 22083 9735 22089
rect 9677 22080 9689 22083
rect 9640 22052 9689 22080
rect 9640 22040 9646 22052
rect 9677 22049 9689 22052
rect 9723 22049 9735 22083
rect 9677 22043 9735 22049
rect 9953 22083 10011 22089
rect 9953 22049 9965 22083
rect 9999 22080 10011 22083
rect 10962 22080 10968 22092
rect 9999 22052 10968 22080
rect 9999 22049 10011 22052
rect 9953 22043 10011 22049
rect 10962 22040 10968 22052
rect 11020 22040 11026 22092
rect 11057 22083 11115 22089
rect 11057 22049 11069 22083
rect 11103 22080 11115 22083
rect 11606 22080 11612 22092
rect 11103 22052 11612 22080
rect 11103 22049 11115 22052
rect 11057 22043 11115 22049
rect 11606 22040 11612 22052
rect 11664 22040 11670 22092
rect 12805 22083 12863 22089
rect 12805 22049 12817 22083
rect 12851 22080 12863 22083
rect 13464 22080 13492 22120
rect 13538 22108 13544 22120
rect 13596 22108 13602 22160
rect 18432 22148 18460 22179
rect 18506 22176 18512 22228
rect 18564 22216 18570 22228
rect 18601 22219 18659 22225
rect 18601 22216 18613 22219
rect 18564 22188 18613 22216
rect 18564 22176 18570 22188
rect 18601 22185 18613 22188
rect 18647 22185 18659 22219
rect 18601 22179 18659 22185
rect 20070 22176 20076 22228
rect 20128 22216 20134 22228
rect 20898 22216 20904 22228
rect 20128 22188 20760 22216
rect 20859 22188 20904 22216
rect 20128 22176 20134 22188
rect 18432 22120 19104 22148
rect 12851 22052 13492 22080
rect 13633 22083 13691 22089
rect 12851 22049 12863 22052
rect 12805 22043 12863 22049
rect 13633 22049 13645 22083
rect 13679 22049 13691 22083
rect 13633 22043 13691 22049
rect 13725 22083 13783 22089
rect 13725 22049 13737 22083
rect 13771 22080 13783 22083
rect 14366 22080 14372 22092
rect 13771 22052 14044 22080
rect 13771 22049 13783 22052
rect 13725 22043 13783 22049
rect 2590 21972 2596 22024
rect 2648 22012 2654 22024
rect 2869 22015 2927 22021
rect 2869 22012 2881 22015
rect 2648 21984 2881 22012
rect 2648 21972 2654 21984
rect 2869 21981 2881 21984
rect 2915 21981 2927 22015
rect 2869 21975 2927 21981
rect 3053 22015 3111 22021
rect 3053 21981 3065 22015
rect 3099 22012 3111 22015
rect 3510 22012 3516 22024
rect 3099 21984 3516 22012
rect 3099 21981 3111 21984
rect 3053 21975 3111 21981
rect 2317 21947 2375 21953
rect 2317 21913 2329 21947
rect 2363 21944 2375 21947
rect 3068 21944 3096 21975
rect 3510 21972 3516 21984
rect 3568 21972 3574 22024
rect 3970 21972 3976 22024
rect 4028 22012 4034 22024
rect 4065 22015 4123 22021
rect 4065 22012 4077 22015
rect 4028 21984 4077 22012
rect 4028 21972 4034 21984
rect 4065 21981 4077 21984
rect 4111 21981 4123 22015
rect 4065 21975 4123 21981
rect 6730 21972 6736 22024
rect 6788 22012 6794 22024
rect 7101 22015 7159 22021
rect 7101 22012 7113 22015
rect 6788 21984 7113 22012
rect 6788 21972 6794 21984
rect 7101 21981 7113 21984
rect 7147 21981 7159 22015
rect 7101 21975 7159 21981
rect 7285 22015 7343 22021
rect 7285 21981 7297 22015
rect 7331 22012 7343 22015
rect 7466 22012 7472 22024
rect 7331 21984 7472 22012
rect 7331 21981 7343 21984
rect 7285 21975 7343 21981
rect 7466 21972 7472 21984
rect 7524 21972 7530 22024
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 9490 22012 9496 22024
rect 8619 21984 9496 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 9490 21972 9496 21984
rect 9548 21972 9554 22024
rect 12618 21972 12624 22024
rect 12676 22012 12682 22024
rect 13081 22015 13139 22021
rect 13081 22012 13093 22015
rect 12676 21984 13093 22012
rect 12676 21972 12682 21984
rect 13081 21981 13093 21984
rect 13127 21981 13139 22015
rect 13081 21975 13139 21981
rect 6086 21944 6092 21956
rect 2363 21916 3096 21944
rect 6047 21916 6092 21944
rect 2363 21913 2375 21916
rect 2317 21907 2375 21913
rect 6086 21904 6092 21916
rect 6144 21904 6150 21956
rect 6641 21947 6699 21953
rect 6641 21913 6653 21947
rect 6687 21944 6699 21947
rect 6822 21944 6828 21956
rect 6687 21916 6828 21944
rect 6687 21913 6699 21916
rect 6641 21907 6699 21913
rect 6822 21904 6828 21916
rect 6880 21904 6886 21956
rect 9030 21944 9036 21956
rect 8991 21916 9036 21944
rect 9030 21904 9036 21916
rect 9088 21904 9094 21956
rect 13096 21944 13124 21975
rect 13170 21972 13176 22024
rect 13228 22012 13234 22024
rect 13648 22012 13676 22043
rect 14016 22024 14044 22052
rect 14200 22052 14372 22080
rect 13906 22012 13912 22024
rect 13228 21984 13676 22012
rect 13867 21984 13912 22012
rect 13228 21972 13234 21984
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 13998 21972 14004 22024
rect 14056 21972 14062 22024
rect 13265 21947 13323 21953
rect 13265 21944 13277 21947
rect 13096 21916 13277 21944
rect 13265 21913 13277 21916
rect 13311 21913 13323 21947
rect 13265 21907 13323 21913
rect 1486 21836 1492 21888
rect 1544 21876 1550 21888
rect 1581 21879 1639 21885
rect 1581 21876 1593 21879
rect 1544 21848 1593 21876
rect 1544 21836 1550 21848
rect 1581 21845 1593 21848
rect 1627 21845 1639 21879
rect 2406 21876 2412 21888
rect 2367 21848 2412 21876
rect 1581 21839 1639 21845
rect 2406 21836 2412 21848
rect 2464 21836 2470 21888
rect 3418 21876 3424 21888
rect 3379 21848 3424 21876
rect 3418 21836 3424 21848
rect 3476 21836 3482 21888
rect 3786 21876 3792 21888
rect 3747 21848 3792 21876
rect 3786 21836 3792 21848
rect 3844 21836 3850 21888
rect 6270 21836 6276 21888
rect 6328 21876 6334 21888
rect 6549 21879 6607 21885
rect 6549 21876 6561 21879
rect 6328 21848 6561 21876
rect 6328 21836 6334 21848
rect 6549 21845 6561 21848
rect 6595 21876 6607 21879
rect 7374 21876 7380 21888
rect 6595 21848 7380 21876
rect 6595 21845 6607 21848
rect 6549 21839 6607 21845
rect 7374 21836 7380 21848
rect 7432 21876 7438 21888
rect 8021 21879 8079 21885
rect 8021 21876 8033 21879
rect 7432 21848 8033 21876
rect 7432 21836 7438 21848
rect 8021 21845 8033 21848
rect 8067 21876 8079 21879
rect 9401 21879 9459 21885
rect 9401 21876 9413 21879
rect 8067 21848 9413 21876
rect 8067 21845 8079 21848
rect 8021 21839 8079 21845
rect 9401 21845 9413 21848
rect 9447 21845 9459 21879
rect 9401 21839 9459 21845
rect 9766 21836 9772 21888
rect 9824 21876 9830 21888
rect 10042 21876 10048 21888
rect 9824 21848 10048 21876
rect 9824 21836 9830 21848
rect 10042 21836 10048 21848
rect 10100 21876 10106 21888
rect 10413 21879 10471 21885
rect 10413 21876 10425 21879
rect 10100 21848 10425 21876
rect 10100 21836 10106 21848
rect 10413 21845 10425 21848
rect 10459 21845 10471 21879
rect 10413 21839 10471 21845
rect 10873 21879 10931 21885
rect 10873 21845 10885 21879
rect 10919 21876 10931 21879
rect 10962 21876 10968 21888
rect 10919 21848 10968 21876
rect 10919 21845 10931 21848
rect 10873 21839 10931 21845
rect 10962 21836 10968 21848
rect 11020 21836 11026 21888
rect 12437 21879 12495 21885
rect 12437 21845 12449 21879
rect 12483 21876 12495 21879
rect 12986 21876 12992 21888
rect 12483 21848 12992 21876
rect 12483 21845 12495 21848
rect 12437 21839 12495 21845
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 13906 21836 13912 21888
rect 13964 21876 13970 21888
rect 14200 21876 14228 22052
rect 14366 22040 14372 22052
rect 14424 22040 14430 22092
rect 15289 22083 15347 22089
rect 15289 22080 15301 22083
rect 15028 22052 15301 22080
rect 14274 21904 14280 21956
rect 14332 21944 14338 21956
rect 14369 21947 14427 21953
rect 14369 21944 14381 21947
rect 14332 21916 14381 21944
rect 14332 21904 14338 21916
rect 14369 21913 14381 21916
rect 14415 21944 14427 21947
rect 14826 21944 14832 21956
rect 14415 21916 14832 21944
rect 14415 21913 14427 21916
rect 14369 21907 14427 21913
rect 14826 21904 14832 21916
rect 14884 21904 14890 21956
rect 14645 21879 14703 21885
rect 14645 21876 14657 21879
rect 13964 21848 14657 21876
rect 13964 21836 13970 21848
rect 14645 21845 14657 21848
rect 14691 21845 14703 21879
rect 14645 21839 14703 21845
rect 14734 21836 14740 21888
rect 14792 21876 14798 21888
rect 15028 21885 15056 22052
rect 15289 22049 15301 22052
rect 15335 22049 15347 22083
rect 15289 22043 15347 22049
rect 16660 22083 16718 22089
rect 16660 22049 16672 22083
rect 16706 22080 16718 22083
rect 17034 22080 17040 22092
rect 16706 22052 17040 22080
rect 16706 22049 16718 22052
rect 16660 22043 16718 22049
rect 17034 22040 17040 22052
rect 17092 22040 17098 22092
rect 18966 22080 18972 22092
rect 18927 22052 18972 22080
rect 18966 22040 18972 22052
rect 19024 22040 19030 22092
rect 19076 22080 19104 22120
rect 20530 22108 20536 22160
rect 20588 22148 20594 22160
rect 20732 22148 20760 22188
rect 20898 22176 20904 22188
rect 20956 22176 20962 22228
rect 21266 22216 21272 22228
rect 21227 22188 21272 22216
rect 21266 22176 21272 22188
rect 21324 22176 21330 22228
rect 22097 22219 22155 22225
rect 22097 22185 22109 22219
rect 22143 22216 22155 22219
rect 22186 22216 22192 22228
rect 22143 22188 22192 22216
rect 22143 22185 22155 22188
rect 22097 22179 22155 22185
rect 22186 22176 22192 22188
rect 22244 22176 22250 22228
rect 23842 22176 23848 22228
rect 23900 22176 23906 22228
rect 23934 22176 23940 22228
rect 23992 22216 23998 22228
rect 24121 22219 24179 22225
rect 24121 22216 24133 22219
rect 23992 22188 24133 22216
rect 23992 22176 23998 22188
rect 24121 22185 24133 22188
rect 24167 22185 24179 22219
rect 24121 22179 24179 22185
rect 21634 22148 21640 22160
rect 20588 22120 20668 22148
rect 20732 22120 21640 22148
rect 20588 22108 20594 22120
rect 20640 22080 20668 22120
rect 21634 22108 21640 22120
rect 21692 22148 21698 22160
rect 22465 22151 22523 22157
rect 21692 22120 22416 22148
rect 21692 22108 21698 22120
rect 19076 22052 19196 22080
rect 20640 22052 21496 22080
rect 15654 21972 15660 22024
rect 15712 22012 15718 22024
rect 15930 22012 15936 22024
rect 15712 21984 15936 22012
rect 15712 21972 15718 21984
rect 15930 21972 15936 21984
rect 15988 22012 15994 22024
rect 16393 22015 16451 22021
rect 16393 22012 16405 22015
rect 15988 21984 16405 22012
rect 15988 21972 15994 21984
rect 16393 21981 16405 21984
rect 16439 21981 16451 22015
rect 16393 21975 16451 21981
rect 17770 21972 17776 22024
rect 17828 22012 17834 22024
rect 19168 22021 19196 22052
rect 19061 22015 19119 22021
rect 19061 22012 19073 22015
rect 17828 21984 19073 22012
rect 17828 21972 17834 21984
rect 19061 21981 19073 21984
rect 19107 21981 19119 22015
rect 19061 21975 19119 21981
rect 19153 22015 19211 22021
rect 19153 21981 19165 22015
rect 19199 21981 19211 22015
rect 21358 22012 21364 22024
rect 21319 21984 21364 22012
rect 19153 21975 19211 21981
rect 21358 21972 21364 21984
rect 21416 21972 21422 22024
rect 21468 22021 21496 22052
rect 21542 22040 21548 22092
rect 21600 22080 21606 22092
rect 21818 22080 21824 22092
rect 21600 22052 21824 22080
rect 21600 22040 21606 22052
rect 21818 22040 21824 22052
rect 21876 22040 21882 22092
rect 22388 22080 22416 22120
rect 22465 22117 22477 22151
rect 22511 22148 22523 22151
rect 22922 22148 22928 22160
rect 22511 22120 22928 22148
rect 22511 22117 22523 22120
rect 22465 22111 22523 22117
rect 22922 22108 22928 22120
rect 22980 22157 22986 22160
rect 22980 22151 23044 22157
rect 22980 22117 22998 22151
rect 23032 22117 23044 22151
rect 23860 22148 23888 22176
rect 23860 22120 24808 22148
rect 22980 22111 23044 22117
rect 22980 22108 22986 22111
rect 22738 22080 22744 22092
rect 22388 22052 22744 22080
rect 22738 22040 22744 22052
rect 22796 22040 22802 22092
rect 24302 22040 24308 22092
rect 24360 22080 24366 22092
rect 24780 22080 24808 22120
rect 24857 22083 24915 22089
rect 24857 22080 24869 22083
rect 24360 22052 24532 22080
rect 24780 22052 24869 22080
rect 24360 22040 24366 22052
rect 21453 22015 21511 22021
rect 21453 21981 21465 22015
rect 21499 22012 21511 22015
rect 22186 22012 22192 22024
rect 21499 21984 22192 22012
rect 21499 21981 21511 21984
rect 21453 21975 21511 21981
rect 22186 21972 22192 21984
rect 22244 21972 22250 22024
rect 24394 21972 24400 22024
rect 24452 21972 24458 22024
rect 15473 21947 15531 21953
rect 15473 21913 15485 21947
rect 15519 21944 15531 21947
rect 16298 21944 16304 21956
rect 15519 21916 16304 21944
rect 15519 21913 15531 21916
rect 15473 21907 15531 21913
rect 16298 21904 16304 21916
rect 16356 21904 16362 21956
rect 19705 21947 19763 21953
rect 19705 21913 19717 21947
rect 19751 21944 19763 21947
rect 20530 21944 20536 21956
rect 19751 21916 20536 21944
rect 19751 21913 19763 21916
rect 19705 21907 19763 21913
rect 20530 21904 20536 21916
rect 20588 21904 20594 21956
rect 21376 21944 21404 21972
rect 21910 21944 21916 21956
rect 21376 21916 21916 21944
rect 21910 21904 21916 21916
rect 21968 21904 21974 21956
rect 24412 21944 24440 21972
rect 23860 21916 24440 21944
rect 23860 21888 23888 21916
rect 15013 21879 15071 21885
rect 15013 21876 15025 21879
rect 14792 21848 15025 21876
rect 14792 21836 14798 21848
rect 15013 21845 15025 21848
rect 15059 21845 15071 21879
rect 15013 21839 15071 21845
rect 15930 21836 15936 21888
rect 15988 21876 15994 21888
rect 16117 21879 16175 21885
rect 16117 21876 16129 21879
rect 15988 21848 16129 21876
rect 15988 21836 15994 21848
rect 16117 21845 16129 21848
rect 16163 21845 16175 21879
rect 16117 21839 16175 21845
rect 16574 21836 16580 21888
rect 16632 21876 16638 21888
rect 17773 21879 17831 21885
rect 17773 21876 17785 21879
rect 16632 21848 17785 21876
rect 16632 21836 16638 21848
rect 17773 21845 17785 21848
rect 17819 21845 17831 21879
rect 19978 21876 19984 21888
rect 19939 21848 19984 21876
rect 17773 21839 17831 21845
rect 19978 21836 19984 21848
rect 20036 21836 20042 21888
rect 20717 21879 20775 21885
rect 20717 21845 20729 21879
rect 20763 21876 20775 21879
rect 21542 21876 21548 21888
rect 20763 21848 21548 21876
rect 20763 21845 20775 21848
rect 20717 21839 20775 21845
rect 21542 21836 21548 21848
rect 21600 21836 21606 21888
rect 23842 21836 23848 21888
rect 23900 21836 23906 21888
rect 24504 21885 24532 22052
rect 24857 22049 24869 22052
rect 24903 22049 24915 22083
rect 24857 22043 24915 22049
rect 24949 22083 25007 22089
rect 24949 22049 24961 22083
rect 24995 22049 25007 22083
rect 24949 22043 25007 22049
rect 24964 22012 24992 22043
rect 24872 21984 24992 22012
rect 25225 22015 25283 22021
rect 24872 21956 24900 21984
rect 25225 21981 25237 22015
rect 25271 22012 25283 22015
rect 26142 22012 26148 22024
rect 25271 21984 26148 22012
rect 25271 21981 25283 21984
rect 25225 21975 25283 21981
rect 26142 21972 26148 21984
rect 26200 21972 26206 22024
rect 24854 21904 24860 21956
rect 24912 21904 24918 21956
rect 24489 21879 24547 21885
rect 24489 21845 24501 21879
rect 24535 21876 24547 21879
rect 24946 21876 24952 21888
rect 24535 21848 24952 21876
rect 24535 21845 24547 21848
rect 24489 21839 24547 21845
rect 24946 21836 24952 21848
rect 25004 21836 25010 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2498 21672 2504 21684
rect 2459 21644 2504 21672
rect 2498 21632 2504 21644
rect 2556 21632 2562 21684
rect 4154 21672 4160 21684
rect 4115 21644 4160 21672
rect 4154 21632 4160 21644
rect 4212 21672 4218 21684
rect 4614 21672 4620 21684
rect 4212 21644 4620 21672
rect 4212 21632 4218 21644
rect 4614 21632 4620 21644
rect 4672 21672 4678 21684
rect 4801 21675 4859 21681
rect 4801 21672 4813 21675
rect 4672 21644 4813 21672
rect 4672 21632 4678 21644
rect 4801 21641 4813 21644
rect 4847 21641 4859 21675
rect 6178 21672 6184 21684
rect 6139 21644 6184 21672
rect 4801 21635 4859 21641
rect 4062 21564 4068 21616
rect 4120 21604 4126 21616
rect 4433 21607 4491 21613
rect 4433 21604 4445 21607
rect 4120 21576 4445 21604
rect 4120 21564 4126 21576
rect 4433 21573 4445 21576
rect 4479 21573 4491 21607
rect 4816 21604 4844 21635
rect 6178 21632 6184 21644
rect 6236 21632 6242 21684
rect 8754 21672 8760 21684
rect 8715 21644 8760 21672
rect 8754 21632 8760 21644
rect 8812 21632 8818 21684
rect 9122 21672 9128 21684
rect 9083 21644 9128 21672
rect 9122 21632 9128 21644
rect 9180 21632 9186 21684
rect 9674 21632 9680 21684
rect 9732 21672 9738 21684
rect 10229 21675 10287 21681
rect 10229 21672 10241 21675
rect 9732 21644 10241 21672
rect 9732 21632 9738 21644
rect 10229 21641 10241 21644
rect 10275 21641 10287 21675
rect 11330 21672 11336 21684
rect 11291 21644 11336 21672
rect 10229 21635 10287 21641
rect 11330 21632 11336 21644
rect 11388 21632 11394 21684
rect 12253 21675 12311 21681
rect 12253 21641 12265 21675
rect 12299 21672 12311 21675
rect 12342 21672 12348 21684
rect 12299 21644 12348 21672
rect 12299 21641 12311 21644
rect 12253 21635 12311 21641
rect 12342 21632 12348 21644
rect 12400 21632 12406 21684
rect 14826 21632 14832 21684
rect 14884 21672 14890 21684
rect 15381 21675 15439 21681
rect 15381 21672 15393 21675
rect 14884 21644 15393 21672
rect 14884 21632 14890 21644
rect 15381 21641 15393 21644
rect 15427 21641 15439 21675
rect 15381 21635 15439 21641
rect 15930 21632 15936 21684
rect 15988 21672 15994 21684
rect 16298 21672 16304 21684
rect 15988 21644 16304 21672
rect 15988 21632 15994 21644
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 19334 21632 19340 21684
rect 19392 21672 19398 21684
rect 19613 21675 19671 21681
rect 19613 21672 19625 21675
rect 19392 21644 19625 21672
rect 19392 21632 19398 21644
rect 19613 21641 19625 21644
rect 19659 21641 19671 21675
rect 21174 21672 21180 21684
rect 21135 21644 21180 21672
rect 19613 21635 19671 21641
rect 21174 21632 21180 21644
rect 21232 21632 21238 21684
rect 22186 21672 22192 21684
rect 22147 21644 22192 21672
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 22833 21675 22891 21681
rect 22833 21641 22845 21675
rect 22879 21672 22891 21675
rect 22922 21672 22928 21684
rect 22879 21644 22928 21672
rect 22879 21641 22891 21644
rect 22833 21635 22891 21641
rect 22922 21632 22928 21644
rect 22980 21632 22986 21684
rect 15289 21607 15347 21613
rect 4816 21576 5580 21604
rect 4433 21567 4491 21573
rect 1762 21536 1768 21548
rect 1723 21508 1768 21536
rect 1762 21496 1768 21508
rect 1820 21496 1826 21548
rect 5442 21536 5448 21548
rect 5403 21508 5448 21536
rect 5442 21496 5448 21508
rect 5500 21496 5506 21548
rect 5552 21545 5580 21576
rect 15289 21573 15301 21607
rect 15335 21604 15347 21607
rect 15838 21604 15844 21616
rect 15335 21576 15844 21604
rect 15335 21573 15347 21576
rect 15289 21567 15347 21573
rect 5537 21539 5595 21545
rect 5537 21505 5549 21539
rect 5583 21505 5595 21539
rect 5537 21499 5595 21505
rect 9122 21496 9128 21548
rect 9180 21536 9186 21548
rect 9398 21536 9404 21548
rect 9180 21508 9404 21536
rect 9180 21496 9186 21508
rect 9398 21496 9404 21508
rect 9456 21496 9462 21548
rect 10042 21496 10048 21548
rect 10100 21536 10106 21548
rect 10781 21539 10839 21545
rect 10781 21536 10793 21539
rect 10100 21508 10793 21536
rect 10100 21496 10106 21508
rect 10781 21505 10793 21508
rect 10827 21505 10839 21539
rect 10781 21499 10839 21505
rect 11885 21539 11943 21545
rect 11885 21505 11897 21539
rect 11931 21536 11943 21539
rect 12342 21536 12348 21548
rect 11931 21508 12348 21536
rect 11931 21505 11943 21508
rect 11885 21499 11943 21505
rect 12342 21496 12348 21508
rect 12400 21496 12406 21548
rect 12713 21539 12771 21545
rect 12713 21505 12725 21539
rect 12759 21536 12771 21539
rect 13722 21536 13728 21548
rect 12759 21508 13728 21536
rect 12759 21505 12771 21508
rect 12713 21499 12771 21505
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 1486 21468 1492 21480
rect 1447 21440 1492 21468
rect 1486 21428 1492 21440
rect 1544 21428 1550 21480
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21468 2835 21471
rect 3970 21468 3976 21480
rect 2823 21440 3976 21468
rect 2823 21437 2835 21440
rect 2777 21431 2835 21437
rect 3970 21428 3976 21440
rect 4028 21428 4034 21480
rect 5258 21428 5264 21480
rect 5316 21468 5322 21480
rect 5353 21471 5411 21477
rect 5353 21468 5365 21471
rect 5316 21440 5365 21468
rect 5316 21428 5322 21440
rect 5353 21437 5365 21440
rect 5399 21437 5411 21471
rect 7374 21468 7380 21480
rect 7335 21440 7380 21468
rect 5353 21431 5411 21437
rect 7374 21428 7380 21440
rect 7432 21428 7438 21480
rect 7650 21477 7656 21480
rect 7644 21468 7656 21477
rect 7563 21440 7656 21468
rect 7644 21431 7656 21440
rect 7708 21468 7714 21480
rect 8202 21468 8208 21480
rect 7708 21440 8208 21468
rect 7650 21428 7656 21431
rect 7708 21428 7714 21440
rect 8202 21428 8208 21440
rect 8260 21428 8266 21480
rect 11054 21428 11060 21480
rect 11112 21468 11118 21480
rect 12158 21468 12164 21480
rect 11112 21440 12164 21468
rect 11112 21428 11118 21440
rect 12158 21428 12164 21440
rect 12216 21468 12222 21480
rect 12437 21471 12495 21477
rect 12437 21468 12449 21471
rect 12216 21440 12449 21468
rect 12216 21428 12222 21440
rect 12437 21437 12449 21440
rect 12483 21437 12495 21471
rect 12437 21431 12495 21437
rect 13909 21471 13967 21477
rect 13909 21437 13921 21471
rect 13955 21468 13967 21471
rect 13955 21440 14136 21468
rect 13955 21437 13967 21440
rect 13909 21431 13967 21437
rect 3044 21403 3102 21409
rect 3044 21369 3056 21403
rect 3090 21400 3102 21403
rect 3510 21400 3516 21412
rect 3090 21372 3516 21400
rect 3090 21369 3102 21372
rect 3044 21363 3102 21369
rect 3510 21360 3516 21372
rect 3568 21360 3574 21412
rect 10689 21403 10747 21409
rect 10689 21400 10701 21403
rect 9692 21372 10701 21400
rect 9692 21344 9720 21372
rect 10689 21369 10701 21372
rect 10735 21369 10747 21403
rect 10689 21363 10747 21369
rect 14108 21344 14136 21440
rect 14642 21428 14648 21480
rect 14700 21468 14706 21480
rect 15304 21468 15332 21567
rect 15838 21564 15844 21576
rect 15896 21604 15902 21616
rect 17770 21604 17776 21616
rect 15896 21576 17540 21604
rect 17731 21576 17776 21604
rect 15896 21564 15902 21576
rect 17512 21545 17540 21576
rect 17770 21564 17776 21576
rect 17828 21564 17834 21616
rect 18506 21564 18512 21616
rect 18564 21604 18570 21616
rect 18966 21604 18972 21616
rect 18564 21576 18972 21604
rect 18564 21564 18570 21576
rect 18966 21564 18972 21576
rect 19024 21604 19030 21616
rect 19061 21607 19119 21613
rect 19061 21604 19073 21607
rect 19024 21576 19073 21604
rect 19024 21564 19030 21576
rect 19061 21573 19073 21576
rect 19107 21573 19119 21607
rect 19061 21567 19119 21573
rect 16761 21539 16819 21545
rect 16761 21505 16773 21539
rect 16807 21505 16819 21539
rect 16761 21499 16819 21505
rect 17497 21539 17555 21545
rect 17497 21505 17509 21539
rect 17543 21536 17555 21539
rect 18601 21539 18659 21545
rect 18601 21536 18613 21539
rect 17543 21508 18613 21536
rect 17543 21505 17555 21508
rect 17497 21499 17555 21505
rect 18601 21505 18613 21508
rect 18647 21505 18659 21539
rect 20257 21539 20315 21545
rect 20257 21536 20269 21539
rect 18601 21499 18659 21505
rect 19352 21508 20269 21536
rect 14700 21440 15332 21468
rect 15381 21471 15439 21477
rect 14700 21428 14706 21440
rect 15381 21437 15393 21471
rect 15427 21468 15439 21471
rect 15657 21471 15715 21477
rect 15657 21468 15669 21471
rect 15427 21440 15669 21468
rect 15427 21437 15439 21440
rect 15381 21431 15439 21437
rect 15657 21437 15669 21440
rect 15703 21468 15715 21471
rect 16666 21468 16672 21480
rect 15703 21440 16672 21468
rect 15703 21437 15715 21440
rect 15657 21431 15715 21437
rect 16666 21428 16672 21440
rect 16724 21468 16730 21480
rect 16776 21468 16804 21499
rect 19352 21468 19380 21508
rect 20257 21505 20269 21508
rect 20303 21536 20315 21539
rect 20530 21536 20536 21548
rect 20303 21508 20536 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 20530 21496 20536 21508
rect 20588 21496 20594 21548
rect 21726 21536 21732 21548
rect 21687 21508 21732 21536
rect 21726 21496 21732 21508
rect 21784 21496 21790 21548
rect 22462 21496 22468 21548
rect 22520 21536 22526 21548
rect 22830 21536 22836 21548
rect 22520 21508 22836 21536
rect 22520 21496 22526 21508
rect 22830 21496 22836 21508
rect 22888 21496 22894 21548
rect 23477 21539 23535 21545
rect 23477 21505 23489 21539
rect 23523 21536 23535 21539
rect 23523 21508 23796 21536
rect 23523 21505 23535 21508
rect 23477 21499 23535 21505
rect 16724 21440 19380 21468
rect 16724 21428 16730 21440
rect 19426 21428 19432 21480
rect 19484 21468 19490 21480
rect 19981 21471 20039 21477
rect 19981 21468 19993 21471
rect 19484 21440 19993 21468
rect 19484 21428 19490 21440
rect 19981 21437 19993 21440
rect 20027 21437 20039 21471
rect 19981 21431 20039 21437
rect 22738 21428 22744 21480
rect 22796 21468 22802 21480
rect 23661 21471 23719 21477
rect 23661 21468 23673 21471
rect 22796 21440 23673 21468
rect 22796 21428 22802 21440
rect 23661 21437 23673 21440
rect 23707 21437 23719 21471
rect 23768 21468 23796 21508
rect 23934 21477 23940 21480
rect 23928 21468 23940 21477
rect 23768 21440 23940 21468
rect 23661 21431 23719 21437
rect 23928 21431 23940 21440
rect 23934 21428 23940 21431
rect 23992 21428 23998 21480
rect 14176 21403 14234 21409
rect 14176 21369 14188 21403
rect 14222 21400 14234 21403
rect 14274 21400 14280 21412
rect 14222 21372 14280 21400
rect 14222 21369 14234 21372
rect 14176 21363 14234 21369
rect 14274 21360 14280 21372
rect 14332 21360 14338 21412
rect 15286 21360 15292 21412
rect 15344 21400 15350 21412
rect 15470 21400 15476 21412
rect 15344 21372 15476 21400
rect 15344 21360 15350 21372
rect 15470 21360 15476 21372
rect 15528 21360 15534 21412
rect 16577 21403 16635 21409
rect 16577 21400 16589 21403
rect 15948 21372 16589 21400
rect 2866 21292 2872 21344
rect 2924 21332 2930 21344
rect 4985 21335 5043 21341
rect 4985 21332 4997 21335
rect 2924 21304 4997 21332
rect 2924 21292 2930 21304
rect 4985 21301 4997 21304
rect 5031 21301 5043 21335
rect 6638 21332 6644 21344
rect 6599 21304 6644 21332
rect 4985 21295 5043 21301
rect 6638 21292 6644 21304
rect 6696 21292 6702 21344
rect 7098 21332 7104 21344
rect 7059 21304 7104 21332
rect 7098 21292 7104 21304
rect 7156 21292 7162 21344
rect 9674 21332 9680 21344
rect 9635 21304 9680 21332
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 10042 21332 10048 21344
rect 10003 21304 10048 21332
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 10597 21335 10655 21341
rect 10597 21301 10609 21335
rect 10643 21332 10655 21335
rect 10962 21332 10968 21344
rect 10643 21304 10968 21332
rect 10643 21301 10655 21304
rect 10597 21295 10655 21301
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 13170 21292 13176 21344
rect 13228 21332 13234 21344
rect 13265 21335 13323 21341
rect 13265 21332 13277 21335
rect 13228 21304 13277 21332
rect 13228 21292 13234 21304
rect 13265 21301 13277 21304
rect 13311 21301 13323 21335
rect 13265 21295 13323 21301
rect 13725 21335 13783 21341
rect 13725 21301 13737 21335
rect 13771 21332 13783 21335
rect 13998 21332 14004 21344
rect 13771 21304 14004 21332
rect 13771 21301 13783 21304
rect 13725 21295 13783 21301
rect 13998 21292 14004 21304
rect 14056 21292 14062 21344
rect 14090 21292 14096 21344
rect 14148 21292 14154 21344
rect 15838 21292 15844 21344
rect 15896 21332 15902 21344
rect 15948 21341 15976 21372
rect 16577 21369 16589 21372
rect 16623 21369 16635 21403
rect 16577 21363 16635 21369
rect 17586 21360 17592 21412
rect 17644 21400 17650 21412
rect 18509 21403 18567 21409
rect 18509 21400 18521 21403
rect 17644 21372 18521 21400
rect 17644 21360 17650 21372
rect 18509 21369 18521 21372
rect 18555 21369 18567 21403
rect 18509 21363 18567 21369
rect 20714 21360 20720 21412
rect 20772 21400 20778 21412
rect 21637 21403 21695 21409
rect 21637 21400 21649 21403
rect 20772 21372 21649 21400
rect 20772 21360 20778 21372
rect 21637 21369 21649 21372
rect 21683 21369 21695 21403
rect 21637 21363 21695 21369
rect 24854 21360 24860 21412
rect 24912 21400 24918 21412
rect 25317 21403 25375 21409
rect 25317 21400 25329 21403
rect 24912 21372 25329 21400
rect 24912 21360 24918 21372
rect 25317 21369 25329 21372
rect 25363 21369 25375 21403
rect 25317 21363 25375 21369
rect 15933 21335 15991 21341
rect 15933 21332 15945 21335
rect 15896 21304 15945 21332
rect 15896 21292 15902 21304
rect 15933 21301 15945 21304
rect 15979 21301 15991 21335
rect 16114 21332 16120 21344
rect 16075 21304 16120 21332
rect 15933 21295 15991 21301
rect 16114 21292 16120 21304
rect 16172 21292 16178 21344
rect 16298 21292 16304 21344
rect 16356 21332 16362 21344
rect 16485 21335 16543 21341
rect 16485 21332 16497 21335
rect 16356 21304 16497 21332
rect 16356 21292 16362 21304
rect 16485 21301 16497 21304
rect 16531 21301 16543 21335
rect 16485 21295 16543 21301
rect 16942 21292 16948 21344
rect 17000 21332 17006 21344
rect 18049 21335 18107 21341
rect 18049 21332 18061 21335
rect 17000 21304 18061 21332
rect 17000 21292 17006 21304
rect 18049 21301 18061 21304
rect 18095 21301 18107 21335
rect 18414 21332 18420 21344
rect 18375 21304 18420 21332
rect 18049 21295 18107 21301
rect 18414 21292 18420 21304
rect 18472 21292 18478 21344
rect 19058 21292 19064 21344
rect 19116 21332 19122 21344
rect 19429 21335 19487 21341
rect 19429 21332 19441 21335
rect 19116 21304 19441 21332
rect 19116 21292 19122 21304
rect 19429 21301 19441 21304
rect 19475 21332 19487 21335
rect 20073 21335 20131 21341
rect 20073 21332 20085 21335
rect 19475 21304 20085 21332
rect 19475 21301 19487 21304
rect 19429 21295 19487 21301
rect 20073 21301 20085 21304
rect 20119 21332 20131 21335
rect 20901 21335 20959 21341
rect 20901 21332 20913 21335
rect 20119 21304 20913 21332
rect 20119 21301 20131 21304
rect 20073 21295 20131 21301
rect 20901 21301 20913 21304
rect 20947 21332 20959 21335
rect 21358 21332 21364 21344
rect 20947 21304 21364 21332
rect 20947 21301 20959 21304
rect 20901 21295 20959 21301
rect 21358 21292 21364 21304
rect 21416 21292 21422 21344
rect 21542 21332 21548 21344
rect 21503 21304 21548 21332
rect 21542 21292 21548 21304
rect 21600 21292 21606 21344
rect 24946 21292 24952 21344
rect 25004 21332 25010 21344
rect 25041 21335 25099 21341
rect 25041 21332 25053 21335
rect 25004 21304 25053 21332
rect 25004 21292 25010 21304
rect 25041 21301 25053 21304
rect 25087 21301 25099 21335
rect 25682 21332 25688 21344
rect 25643 21304 25688 21332
rect 25041 21295 25099 21301
rect 25682 21292 25688 21304
rect 25740 21292 25746 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1486 21088 1492 21140
rect 1544 21128 1550 21140
rect 2409 21131 2467 21137
rect 2409 21128 2421 21131
rect 1544 21100 2421 21128
rect 1544 21088 1550 21100
rect 2409 21097 2421 21100
rect 2455 21097 2467 21131
rect 2409 21091 2467 21097
rect 5169 21131 5227 21137
rect 5169 21097 5181 21131
rect 5215 21128 5227 21131
rect 5442 21128 5448 21140
rect 5215 21100 5448 21128
rect 5215 21097 5227 21100
rect 5169 21091 5227 21097
rect 5442 21088 5448 21100
rect 5500 21088 5506 21140
rect 6181 21131 6239 21137
rect 6181 21097 6193 21131
rect 6227 21128 6239 21131
rect 6270 21128 6276 21140
rect 6227 21100 6276 21128
rect 6227 21097 6239 21100
rect 6181 21091 6239 21097
rect 6270 21088 6276 21100
rect 6328 21088 6334 21140
rect 7561 21131 7619 21137
rect 7561 21097 7573 21131
rect 7607 21128 7619 21131
rect 7650 21128 7656 21140
rect 7607 21100 7656 21128
rect 7607 21097 7619 21100
rect 7561 21091 7619 21097
rect 7650 21088 7656 21100
rect 7708 21088 7714 21140
rect 8018 21128 8024 21140
rect 7979 21100 8024 21128
rect 8018 21088 8024 21100
rect 8076 21088 8082 21140
rect 8294 21088 8300 21140
rect 8352 21128 8358 21140
rect 8389 21131 8447 21137
rect 8389 21128 8401 21131
rect 8352 21100 8401 21128
rect 8352 21088 8358 21100
rect 8389 21097 8401 21100
rect 8435 21128 8447 21131
rect 8570 21128 8576 21140
rect 8435 21100 8576 21128
rect 8435 21097 8447 21100
rect 8389 21091 8447 21097
rect 8570 21088 8576 21100
rect 8628 21088 8634 21140
rect 11238 21088 11244 21140
rect 11296 21128 11302 21140
rect 12345 21131 12403 21137
rect 12345 21128 12357 21131
rect 11296 21100 12357 21128
rect 11296 21088 11302 21100
rect 12345 21097 12357 21100
rect 12391 21097 12403 21131
rect 12345 21091 12403 21097
rect 12618 21088 12624 21140
rect 12676 21128 12682 21140
rect 12805 21131 12863 21137
rect 12805 21128 12817 21131
rect 12676 21100 12817 21128
rect 12676 21088 12682 21100
rect 12805 21097 12817 21100
rect 12851 21097 12863 21131
rect 13446 21128 13452 21140
rect 13407 21100 13452 21128
rect 12805 21091 12863 21097
rect 13446 21088 13452 21100
rect 13504 21088 13510 21140
rect 16114 21088 16120 21140
rect 16172 21128 16178 21140
rect 17221 21131 17279 21137
rect 17221 21128 17233 21131
rect 16172 21100 17233 21128
rect 16172 21088 16178 21100
rect 17221 21097 17233 21100
rect 17267 21128 17279 21131
rect 18414 21128 18420 21140
rect 17267 21100 18420 21128
rect 17267 21097 17279 21100
rect 17221 21091 17279 21097
rect 18414 21088 18420 21100
rect 18472 21088 18478 21140
rect 19334 21088 19340 21140
rect 19392 21128 19398 21140
rect 19981 21131 20039 21137
rect 19981 21128 19993 21131
rect 19392 21100 19993 21128
rect 19392 21088 19398 21100
rect 19981 21097 19993 21100
rect 20027 21128 20039 21131
rect 20070 21128 20076 21140
rect 20027 21100 20076 21128
rect 20027 21097 20039 21100
rect 19981 21091 20039 21097
rect 20070 21088 20076 21100
rect 20128 21088 20134 21140
rect 20714 21128 20720 21140
rect 20675 21100 20720 21128
rect 20714 21088 20720 21100
rect 20772 21088 20778 21140
rect 21177 21131 21235 21137
rect 21177 21097 21189 21131
rect 21223 21128 21235 21131
rect 21266 21128 21272 21140
rect 21223 21100 21272 21128
rect 21223 21097 21235 21100
rect 21177 21091 21235 21097
rect 21266 21088 21272 21100
rect 21324 21088 21330 21140
rect 21545 21131 21603 21137
rect 21545 21097 21557 21131
rect 21591 21128 21603 21131
rect 21726 21128 21732 21140
rect 21591 21100 21732 21128
rect 21591 21097 21603 21100
rect 21545 21091 21603 21097
rect 2866 21060 2872 21072
rect 2827 21032 2872 21060
rect 2866 21020 2872 21032
rect 2924 21020 2930 21072
rect 3513 21063 3571 21069
rect 3513 21029 3525 21063
rect 3559 21060 3571 21063
rect 3602 21060 3608 21072
rect 3559 21032 3608 21060
rect 3559 21029 3571 21032
rect 3513 21023 3571 21029
rect 3602 21020 3608 21032
rect 3660 21020 3666 21072
rect 4154 21020 4160 21072
rect 4212 21060 4218 21072
rect 4525 21063 4583 21069
rect 4525 21060 4537 21063
rect 4212 21032 4537 21060
rect 4212 21020 4218 21032
rect 4525 21029 4537 21032
rect 4571 21029 4583 21063
rect 4525 21023 4583 21029
rect 7929 21063 7987 21069
rect 7929 21029 7941 21063
rect 7975 21060 7987 21063
rect 8110 21060 8116 21072
rect 7975 21032 8116 21060
rect 7975 21029 7987 21032
rect 7929 21023 7987 21029
rect 8110 21020 8116 21032
rect 8168 21020 8174 21072
rect 11606 21060 11612 21072
rect 10060 21032 11612 21060
rect 2317 20995 2375 21001
rect 2317 20961 2329 20995
rect 2363 20992 2375 20995
rect 2590 20992 2596 21004
rect 2363 20964 2596 20992
rect 2363 20961 2375 20964
rect 2317 20955 2375 20961
rect 2590 20952 2596 20964
rect 2648 20952 2654 21004
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20992 2835 20995
rect 3697 20995 3755 21001
rect 3697 20992 3709 20995
rect 2823 20964 3709 20992
rect 2823 20961 2835 20964
rect 2777 20955 2835 20961
rect 3697 20961 3709 20964
rect 3743 20961 3755 20995
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 3697 20955 3755 20961
rect 4172 20964 4445 20992
rect 1394 20924 1400 20936
rect 1355 20896 1400 20924
rect 1394 20884 1400 20896
rect 1452 20884 1458 20936
rect 1949 20927 2007 20933
rect 1949 20893 1961 20927
rect 1995 20924 2007 20927
rect 2866 20924 2872 20936
rect 1995 20896 2872 20924
rect 1995 20893 2007 20896
rect 1949 20887 2007 20893
rect 2866 20884 2872 20896
rect 2924 20884 2930 20936
rect 3053 20927 3111 20933
rect 3053 20893 3065 20927
rect 3099 20924 3111 20927
rect 4062 20924 4068 20936
rect 3099 20896 4068 20924
rect 3099 20893 3111 20896
rect 3053 20887 3111 20893
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 2498 20816 2504 20868
rect 2556 20856 2562 20868
rect 3789 20859 3847 20865
rect 3789 20856 3801 20859
rect 2556 20828 3801 20856
rect 2556 20816 2562 20828
rect 3789 20825 3801 20828
rect 3835 20856 3847 20859
rect 4172 20856 4200 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 5258 20952 5264 21004
rect 5316 20992 5322 21004
rect 5445 20995 5503 21001
rect 5445 20992 5457 20995
rect 5316 20964 5457 20992
rect 5316 20952 5322 20964
rect 5445 20961 5457 20964
rect 5491 20961 5503 20995
rect 5445 20955 5503 20961
rect 6086 20952 6092 21004
rect 6144 20992 6150 21004
rect 6365 20995 6423 21001
rect 6365 20992 6377 20995
rect 6144 20964 6377 20992
rect 6144 20952 6150 20964
rect 6365 20961 6377 20964
rect 6411 20961 6423 20995
rect 6365 20955 6423 20961
rect 6546 20952 6552 21004
rect 6604 20992 6610 21004
rect 6825 20995 6883 21001
rect 6825 20992 6837 20995
rect 6604 20964 6837 20992
rect 6604 20952 6610 20964
rect 6825 20961 6837 20964
rect 6871 20992 6883 20995
rect 8294 20992 8300 21004
rect 6871 20964 8300 20992
rect 6871 20961 6883 20964
rect 6825 20955 6883 20961
rect 8294 20952 8300 20964
rect 8352 20952 8358 21004
rect 9766 20952 9772 21004
rect 9824 20992 9830 21004
rect 10060 21001 10088 21032
rect 11606 21020 11612 21032
rect 11664 21020 11670 21072
rect 12158 21060 12164 21072
rect 12119 21032 12164 21060
rect 12158 21020 12164 21032
rect 12216 21020 12222 21072
rect 13814 21020 13820 21072
rect 13872 21060 13878 21072
rect 15013 21063 15071 21069
rect 15013 21060 15025 21063
rect 13872 21032 15025 21060
rect 13872 21020 13878 21032
rect 15013 21029 15025 21032
rect 15059 21060 15071 21063
rect 15657 21063 15715 21069
rect 15657 21060 15669 21063
rect 15059 21032 15669 21060
rect 15059 21029 15071 21032
rect 15013 21023 15071 21029
rect 15657 21029 15669 21032
rect 15703 21029 15715 21063
rect 15657 21023 15715 21029
rect 16853 21063 16911 21069
rect 16853 21029 16865 21063
rect 16899 21060 16911 21063
rect 16942 21060 16948 21072
rect 16899 21032 16948 21060
rect 16899 21029 16911 21032
rect 16853 21023 16911 21029
rect 16942 21020 16948 21032
rect 17000 21020 17006 21072
rect 17586 21060 17592 21072
rect 17547 21032 17592 21060
rect 17586 21020 17592 21032
rect 17644 21020 17650 21072
rect 18040 21063 18098 21069
rect 18040 21029 18052 21063
rect 18086 21060 18098 21063
rect 19150 21060 19156 21072
rect 18086 21032 19156 21060
rect 18086 21029 18098 21032
rect 18040 21023 18098 21029
rect 19150 21020 19156 21032
rect 19208 21020 19214 21072
rect 20806 21020 20812 21072
rect 20864 21060 20870 21072
rect 21560 21060 21588 21091
rect 21726 21088 21732 21100
rect 21784 21088 21790 21140
rect 22002 21088 22008 21140
rect 22060 21128 22066 21140
rect 22189 21131 22247 21137
rect 22189 21128 22201 21131
rect 22060 21100 22201 21128
rect 22060 21088 22066 21100
rect 22189 21097 22201 21100
rect 22235 21097 22247 21131
rect 22189 21091 22247 21097
rect 22738 21088 22744 21140
rect 22796 21128 22802 21140
rect 22833 21131 22891 21137
rect 22833 21128 22845 21131
rect 22796 21100 22845 21128
rect 22796 21088 22802 21100
rect 22833 21097 22845 21100
rect 22879 21128 22891 21131
rect 23109 21131 23167 21137
rect 23109 21128 23121 21131
rect 22879 21100 23121 21128
rect 22879 21097 22891 21100
rect 22833 21091 22891 21097
rect 23109 21097 23121 21100
rect 23155 21128 23167 21131
rect 23201 21131 23259 21137
rect 23201 21128 23213 21131
rect 23155 21100 23213 21128
rect 23155 21097 23167 21100
rect 23109 21091 23167 21097
rect 23201 21097 23213 21100
rect 23247 21097 23259 21131
rect 23201 21091 23259 21097
rect 23934 21088 23940 21140
rect 23992 21128 23998 21140
rect 24765 21131 24823 21137
rect 24765 21128 24777 21131
rect 23992 21100 24777 21128
rect 23992 21088 23998 21100
rect 24765 21097 24777 21100
rect 24811 21097 24823 21131
rect 24765 21091 24823 21097
rect 20864 21032 21588 21060
rect 20864 21020 20870 21032
rect 10318 21001 10324 21004
rect 10045 20995 10103 21001
rect 10045 20992 10057 20995
rect 9824 20964 10057 20992
rect 9824 20952 9830 20964
rect 10045 20961 10057 20964
rect 10091 20961 10103 20995
rect 10312 20992 10324 21001
rect 10045 20955 10103 20961
rect 10152 20964 10324 20992
rect 4614 20924 4620 20936
rect 4575 20896 4620 20924
rect 4614 20884 4620 20896
rect 4672 20884 4678 20936
rect 6914 20924 6920 20936
rect 6875 20896 6920 20924
rect 6914 20884 6920 20896
rect 6972 20884 6978 20936
rect 7009 20927 7067 20933
rect 7009 20893 7021 20927
rect 7055 20893 7067 20927
rect 7009 20887 7067 20893
rect 3835 20828 4200 20856
rect 3835 20825 3847 20828
rect 3789 20819 3847 20825
rect 6730 20816 6736 20868
rect 6788 20856 6794 20868
rect 7024 20856 7052 20887
rect 7558 20884 7564 20936
rect 7616 20924 7622 20936
rect 8481 20927 8539 20933
rect 8481 20924 8493 20927
rect 7616 20896 8493 20924
rect 7616 20884 7622 20896
rect 8481 20893 8493 20896
rect 8527 20893 8539 20927
rect 8481 20887 8539 20893
rect 8662 20884 8668 20936
rect 8720 20924 8726 20936
rect 10152 20924 10180 20964
rect 10312 20955 10324 20964
rect 10318 20952 10324 20955
rect 10376 20952 10382 21004
rect 12713 20995 12771 21001
rect 12713 20961 12725 20995
rect 12759 20992 12771 20995
rect 13354 20992 13360 21004
rect 12759 20964 13360 20992
rect 12759 20961 12771 20964
rect 12713 20955 12771 20961
rect 13354 20952 13360 20964
rect 13412 20952 13418 21004
rect 13909 20995 13967 21001
rect 13909 20961 13921 20995
rect 13955 20992 13967 20995
rect 16485 20995 16543 21001
rect 13955 20964 14780 20992
rect 13955 20961 13967 20964
rect 13909 20955 13967 20961
rect 8720 20896 10180 20924
rect 12989 20927 13047 20933
rect 8720 20884 8726 20896
rect 12989 20893 13001 20927
rect 13035 20924 13047 20927
rect 13446 20924 13452 20936
rect 13035 20896 13452 20924
rect 13035 20893 13047 20896
rect 12989 20887 13047 20893
rect 13446 20884 13452 20896
rect 13504 20924 13510 20936
rect 13814 20924 13820 20936
rect 13504 20896 13820 20924
rect 13504 20884 13510 20896
rect 13814 20884 13820 20896
rect 13872 20884 13878 20936
rect 14185 20927 14243 20933
rect 14185 20893 14197 20927
rect 14231 20924 14243 20927
rect 14274 20924 14280 20936
rect 14231 20896 14280 20924
rect 14231 20893 14243 20896
rect 14185 20887 14243 20893
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 6788 20828 7052 20856
rect 6788 20816 6794 20828
rect 3510 20748 3516 20800
rect 3568 20788 3574 20800
rect 3697 20791 3755 20797
rect 3697 20788 3709 20791
rect 3568 20760 3709 20788
rect 3568 20748 3574 20760
rect 3697 20757 3709 20760
rect 3743 20788 3755 20791
rect 4065 20791 4123 20797
rect 4065 20788 4077 20791
rect 3743 20760 4077 20788
rect 3743 20757 3755 20760
rect 3697 20751 3755 20757
rect 4065 20757 4077 20760
rect 4111 20757 4123 20791
rect 6086 20788 6092 20800
rect 6047 20760 6092 20788
rect 4065 20751 4123 20757
rect 6086 20748 6092 20760
rect 6144 20748 6150 20800
rect 6457 20791 6515 20797
rect 6457 20757 6469 20791
rect 6503 20788 6515 20791
rect 6914 20788 6920 20800
rect 6503 20760 6920 20788
rect 6503 20757 6515 20760
rect 6457 20751 6515 20757
rect 6914 20748 6920 20760
rect 6972 20748 6978 20800
rect 9125 20791 9183 20797
rect 9125 20757 9137 20791
rect 9171 20788 9183 20791
rect 9398 20788 9404 20800
rect 9171 20760 9404 20788
rect 9171 20757 9183 20760
rect 9125 20751 9183 20757
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 9493 20791 9551 20797
rect 9493 20757 9505 20791
rect 9539 20788 9551 20791
rect 9674 20788 9680 20800
rect 9539 20760 9680 20788
rect 9539 20757 9551 20760
rect 9493 20751 9551 20757
rect 9674 20748 9680 20760
rect 9732 20748 9738 20800
rect 9953 20791 10011 20797
rect 9953 20757 9965 20791
rect 9999 20788 10011 20791
rect 10042 20788 10048 20800
rect 9999 20760 10048 20788
rect 9999 20757 10011 20760
rect 9953 20751 10011 20757
rect 10042 20748 10048 20760
rect 10100 20788 10106 20800
rect 11425 20791 11483 20797
rect 11425 20788 11437 20791
rect 10100 20760 11437 20788
rect 10100 20748 10106 20760
rect 11425 20757 11437 20760
rect 11471 20757 11483 20791
rect 11425 20751 11483 20757
rect 11885 20791 11943 20797
rect 11885 20757 11897 20791
rect 11931 20788 11943 20791
rect 12342 20788 12348 20800
rect 11931 20760 12348 20788
rect 11931 20757 11943 20760
rect 11885 20751 11943 20757
rect 12342 20748 12348 20760
rect 12400 20748 12406 20800
rect 13725 20791 13783 20797
rect 13725 20757 13737 20791
rect 13771 20788 13783 20791
rect 13906 20788 13912 20800
rect 13771 20760 13912 20788
rect 13771 20757 13783 20760
rect 13725 20751 13783 20757
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 14752 20797 14780 20964
rect 16485 20961 16497 20995
rect 16531 20992 16543 20995
rect 17034 20992 17040 21004
rect 16531 20964 17040 20992
rect 16531 20961 16543 20964
rect 16485 20955 16543 20961
rect 17034 20952 17040 20964
rect 17092 20992 17098 21004
rect 20162 20992 20168 21004
rect 17092 20964 19196 20992
rect 20123 20964 20168 20992
rect 17092 20952 17098 20964
rect 15470 20884 15476 20936
rect 15528 20924 15534 20936
rect 15749 20927 15807 20933
rect 15749 20924 15761 20927
rect 15528 20896 15761 20924
rect 15528 20884 15534 20896
rect 15749 20893 15761 20896
rect 15795 20893 15807 20927
rect 15749 20887 15807 20893
rect 15933 20927 15991 20933
rect 15933 20893 15945 20927
rect 15979 20924 15991 20927
rect 16114 20924 16120 20936
rect 15979 20896 16120 20924
rect 15979 20893 15991 20896
rect 15933 20887 15991 20893
rect 16114 20884 16120 20896
rect 16172 20884 16178 20936
rect 17773 20927 17831 20933
rect 17773 20893 17785 20927
rect 17819 20893 17831 20927
rect 17773 20887 17831 20893
rect 15289 20859 15347 20865
rect 15289 20825 15301 20859
rect 15335 20856 15347 20859
rect 15838 20856 15844 20868
rect 15335 20828 15844 20856
rect 15335 20825 15347 20828
rect 15289 20819 15347 20825
rect 15838 20816 15844 20828
rect 15896 20816 15902 20868
rect 14737 20791 14795 20797
rect 14737 20757 14749 20791
rect 14783 20788 14795 20791
rect 14826 20788 14832 20800
rect 14783 20760 14832 20788
rect 14783 20757 14795 20760
rect 14737 20751 14795 20757
rect 14826 20748 14832 20760
rect 14884 20748 14890 20800
rect 17788 20788 17816 20887
rect 19168 20865 19196 20964
rect 20162 20952 20168 20964
rect 20220 20952 20226 21004
rect 23641 20995 23699 21001
rect 23641 20992 23653 20995
rect 23032 20964 23653 20992
rect 23032 20936 23060 20964
rect 23641 20961 23653 20964
rect 23687 20992 23699 20995
rect 24946 20992 24952 21004
rect 23687 20964 24952 20992
rect 23687 20961 23699 20964
rect 23641 20955 23699 20961
rect 24946 20952 24952 20964
rect 25004 20952 25010 21004
rect 22186 20884 22192 20936
rect 22244 20924 22250 20936
rect 22281 20927 22339 20933
rect 22281 20924 22293 20927
rect 22244 20896 22293 20924
rect 22244 20884 22250 20896
rect 22281 20893 22293 20896
rect 22327 20893 22339 20927
rect 22281 20887 22339 20893
rect 22465 20927 22523 20933
rect 22465 20893 22477 20927
rect 22511 20924 22523 20927
rect 23014 20924 23020 20936
rect 22511 20896 23020 20924
rect 22511 20893 22523 20896
rect 22465 20887 22523 20893
rect 23014 20884 23020 20896
rect 23072 20884 23078 20936
rect 23109 20927 23167 20933
rect 23109 20893 23121 20927
rect 23155 20924 23167 20927
rect 23385 20927 23443 20933
rect 23385 20924 23397 20927
rect 23155 20896 23397 20924
rect 23155 20893 23167 20896
rect 23109 20887 23167 20893
rect 23385 20893 23397 20896
rect 23431 20893 23443 20927
rect 23385 20887 23443 20893
rect 19153 20859 19211 20865
rect 19153 20825 19165 20859
rect 19199 20825 19211 20859
rect 19153 20819 19211 20825
rect 17954 20788 17960 20800
rect 17788 20760 17960 20788
rect 17954 20748 17960 20760
rect 18012 20748 18018 20800
rect 19426 20748 19432 20800
rect 19484 20788 19490 20800
rect 19613 20791 19671 20797
rect 19613 20788 19625 20791
rect 19484 20760 19625 20788
rect 19484 20748 19490 20760
rect 19613 20757 19625 20760
rect 19659 20757 19671 20791
rect 21818 20788 21824 20800
rect 21779 20760 21824 20788
rect 19613 20751 19671 20757
rect 21818 20748 21824 20760
rect 21876 20748 21882 20800
rect 25038 20788 25044 20800
rect 24999 20760 25044 20788
rect 25038 20748 25044 20760
rect 25096 20788 25102 20800
rect 25409 20791 25467 20797
rect 25409 20788 25421 20791
rect 25096 20760 25421 20788
rect 25096 20748 25102 20760
rect 25409 20757 25421 20760
rect 25455 20788 25467 20791
rect 25682 20788 25688 20800
rect 25455 20760 25688 20788
rect 25455 20757 25467 20760
rect 25409 20751 25467 20757
rect 25682 20748 25688 20760
rect 25740 20748 25746 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2498 20584 2504 20596
rect 2459 20556 2504 20584
rect 2498 20544 2504 20556
rect 2556 20544 2562 20596
rect 3973 20587 4031 20593
rect 3973 20553 3985 20587
rect 4019 20584 4031 20587
rect 4062 20584 4068 20596
rect 4019 20556 4068 20584
rect 4019 20553 4031 20556
rect 3973 20547 4031 20553
rect 4062 20544 4068 20556
rect 4120 20544 4126 20596
rect 5905 20587 5963 20593
rect 5905 20553 5917 20587
rect 5951 20584 5963 20587
rect 5994 20584 6000 20596
rect 5951 20556 6000 20584
rect 5951 20553 5963 20556
rect 5905 20547 5963 20553
rect 5994 20544 6000 20556
rect 6052 20544 6058 20596
rect 6546 20584 6552 20596
rect 6507 20556 6552 20584
rect 6546 20544 6552 20556
rect 6604 20544 6610 20596
rect 7006 20544 7012 20596
rect 7064 20584 7070 20596
rect 7101 20587 7159 20593
rect 7101 20584 7113 20587
rect 7064 20556 7113 20584
rect 7064 20544 7070 20556
rect 7101 20553 7113 20556
rect 7147 20584 7159 20587
rect 7558 20584 7564 20596
rect 7147 20556 7564 20584
rect 7147 20553 7159 20556
rect 7101 20547 7159 20553
rect 7558 20544 7564 20556
rect 7616 20544 7622 20596
rect 10778 20544 10784 20596
rect 10836 20584 10842 20596
rect 11241 20587 11299 20593
rect 11241 20584 11253 20587
rect 10836 20556 11253 20584
rect 10836 20544 10842 20556
rect 11241 20553 11253 20556
rect 11287 20553 11299 20587
rect 11241 20547 11299 20553
rect 11790 20544 11796 20596
rect 11848 20584 11854 20596
rect 11977 20587 12035 20593
rect 11977 20584 11989 20587
rect 11848 20556 11989 20584
rect 11848 20544 11854 20556
rect 11977 20553 11989 20556
rect 12023 20584 12035 20587
rect 13814 20584 13820 20596
rect 12023 20556 12848 20584
rect 13775 20556 13820 20584
rect 12023 20553 12035 20556
rect 11977 20547 12035 20553
rect 12820 20528 12848 20556
rect 13814 20544 13820 20556
rect 13872 20544 13878 20596
rect 14826 20544 14832 20596
rect 14884 20584 14890 20596
rect 16301 20587 16359 20593
rect 16301 20584 16313 20587
rect 14884 20556 16313 20584
rect 14884 20544 14890 20556
rect 16301 20553 16313 20556
rect 16347 20553 16359 20587
rect 19242 20584 19248 20596
rect 16301 20547 16359 20553
rect 19076 20556 19248 20584
rect 12802 20476 12808 20528
rect 12860 20476 12866 20528
rect 15378 20476 15384 20528
rect 15436 20516 15442 20528
rect 15473 20519 15531 20525
rect 15473 20516 15485 20519
rect 15436 20488 15485 20516
rect 15436 20476 15442 20488
rect 15473 20485 15485 20488
rect 15519 20516 15531 20519
rect 16117 20519 16175 20525
rect 16117 20516 16129 20519
rect 15519 20488 16129 20516
rect 15519 20485 15531 20488
rect 15473 20479 15531 20485
rect 16117 20485 16129 20488
rect 16163 20516 16175 20519
rect 16163 20488 16896 20516
rect 16163 20485 16175 20488
rect 16117 20479 16175 20485
rect 3142 20448 3148 20460
rect 3055 20420 3148 20448
rect 3142 20408 3148 20420
rect 3200 20448 3206 20460
rect 3602 20448 3608 20460
rect 3200 20420 3608 20448
rect 3200 20408 3206 20420
rect 3602 20408 3608 20420
rect 3660 20408 3666 20460
rect 3970 20408 3976 20460
rect 4028 20448 4034 20460
rect 4522 20448 4528 20460
rect 4028 20420 4528 20448
rect 4028 20408 4034 20420
rect 4522 20408 4528 20420
rect 4580 20408 4586 20460
rect 9766 20408 9772 20460
rect 9824 20448 9830 20460
rect 9861 20451 9919 20457
rect 9861 20448 9873 20451
rect 9824 20420 9873 20448
rect 9824 20408 9830 20420
rect 9861 20417 9873 20420
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 11609 20451 11667 20457
rect 11609 20417 11621 20451
rect 11655 20448 11667 20451
rect 11698 20448 11704 20460
rect 11655 20420 11704 20448
rect 11655 20417 11667 20420
rect 11609 20411 11667 20417
rect 11698 20408 11704 20420
rect 11756 20448 11762 20460
rect 12986 20448 12992 20460
rect 11756 20420 12204 20448
rect 12947 20420 12992 20448
rect 11756 20408 11762 20420
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 2406 20380 2412 20392
rect 1443 20352 2084 20380
rect 2367 20352 2412 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 2056 20256 2084 20352
rect 2406 20340 2412 20352
rect 2464 20380 2470 20392
rect 2961 20383 3019 20389
rect 2961 20380 2973 20383
rect 2464 20352 2973 20380
rect 2464 20340 2470 20352
rect 2961 20349 2973 20352
rect 3007 20349 3019 20383
rect 2961 20343 3019 20349
rect 7374 20340 7380 20392
rect 7432 20380 7438 20392
rect 7653 20383 7711 20389
rect 7653 20380 7665 20383
rect 7432 20352 7665 20380
rect 7432 20340 7438 20352
rect 7653 20349 7665 20352
rect 7699 20380 7711 20383
rect 9398 20380 9404 20392
rect 7699 20352 9404 20380
rect 7699 20349 7711 20352
rect 7653 20343 7711 20349
rect 9398 20340 9404 20352
rect 9456 20340 9462 20392
rect 9677 20383 9735 20389
rect 9677 20349 9689 20383
rect 9723 20380 9735 20383
rect 11974 20380 11980 20392
rect 9723 20352 11980 20380
rect 9723 20349 9735 20352
rect 9677 20343 9735 20349
rect 10336 20324 10364 20352
rect 11974 20340 11980 20352
rect 12032 20340 12038 20392
rect 4770 20315 4828 20321
rect 4770 20312 4782 20315
rect 4356 20284 4782 20312
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 2038 20244 2044 20256
rect 1999 20216 2044 20244
rect 2038 20204 2044 20216
rect 2096 20204 2102 20256
rect 2866 20204 2872 20256
rect 2924 20244 2930 20256
rect 3513 20247 3571 20253
rect 3513 20244 3525 20247
rect 2924 20216 3525 20244
rect 2924 20204 2930 20216
rect 3513 20213 3525 20216
rect 3559 20213 3571 20247
rect 3513 20207 3571 20213
rect 3602 20204 3608 20256
rect 3660 20244 3666 20256
rect 4356 20253 4384 20284
rect 4770 20281 4782 20284
rect 4816 20312 4828 20315
rect 5534 20312 5540 20324
rect 4816 20284 5540 20312
rect 4816 20281 4828 20284
rect 4770 20275 4828 20281
rect 5534 20272 5540 20284
rect 5592 20272 5598 20324
rect 7920 20315 7978 20321
rect 7920 20281 7932 20315
rect 7966 20312 7978 20315
rect 8110 20312 8116 20324
rect 7966 20284 8116 20312
rect 7966 20281 7978 20284
rect 7920 20275 7978 20281
rect 8110 20272 8116 20284
rect 8168 20272 8174 20324
rect 10042 20272 10048 20324
rect 10100 20321 10106 20324
rect 10100 20315 10164 20321
rect 10100 20281 10118 20315
rect 10152 20281 10164 20315
rect 10100 20275 10164 20281
rect 10100 20272 10106 20275
rect 10318 20272 10324 20324
rect 10376 20272 10382 20324
rect 11606 20272 11612 20324
rect 11664 20312 11670 20324
rect 12176 20312 12204 20420
rect 12986 20408 12992 20420
rect 13044 20408 13050 20460
rect 16868 20457 16896 20488
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 17954 20408 17960 20460
rect 18012 20448 18018 20460
rect 19076 20457 19104 20556
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 23661 20587 23719 20593
rect 23661 20553 23673 20587
rect 23707 20584 23719 20587
rect 24762 20584 24768 20596
rect 23707 20556 24768 20584
rect 23707 20553 23719 20556
rect 23661 20547 23719 20553
rect 24762 20544 24768 20556
rect 24820 20544 24826 20596
rect 19061 20451 19119 20457
rect 19061 20448 19073 20451
rect 18012 20420 19073 20448
rect 18012 20408 18018 20420
rect 19061 20417 19073 20420
rect 19107 20417 19119 20451
rect 19061 20411 19119 20417
rect 20070 20408 20076 20460
rect 20128 20448 20134 20460
rect 21269 20451 21327 20457
rect 21269 20448 21281 20451
rect 20128 20420 21281 20448
rect 20128 20408 20134 20420
rect 21269 20417 21281 20420
rect 21315 20417 21327 20451
rect 24118 20448 24124 20460
rect 24079 20420 24124 20448
rect 21269 20411 21327 20417
rect 24118 20408 24124 20420
rect 24176 20408 24182 20460
rect 24302 20448 24308 20460
rect 24263 20420 24308 20448
rect 24302 20408 24308 20420
rect 24360 20408 24366 20460
rect 25130 20408 25136 20460
rect 25188 20448 25194 20460
rect 25409 20451 25467 20457
rect 25409 20448 25421 20451
rect 25188 20420 25421 20448
rect 25188 20408 25194 20420
rect 25409 20417 25421 20420
rect 25455 20417 25467 20451
rect 25409 20411 25467 20417
rect 12253 20383 12311 20389
rect 12253 20349 12265 20383
rect 12299 20380 12311 20383
rect 12342 20380 12348 20392
rect 12299 20352 12348 20380
rect 12299 20349 12311 20352
rect 12253 20343 12311 20349
rect 12342 20340 12348 20352
rect 12400 20340 12406 20392
rect 12802 20380 12808 20392
rect 12763 20352 12808 20380
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 14090 20380 14096 20392
rect 14003 20352 14096 20380
rect 14090 20340 14096 20352
rect 14148 20340 14154 20392
rect 14360 20383 14418 20389
rect 14360 20349 14372 20383
rect 14406 20380 14418 20383
rect 14642 20380 14648 20392
rect 14406 20352 14648 20380
rect 14406 20349 14418 20352
rect 14360 20343 14418 20349
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 16574 20340 16580 20392
rect 16632 20380 16638 20392
rect 16669 20383 16727 20389
rect 16669 20380 16681 20383
rect 16632 20352 16681 20380
rect 16632 20340 16638 20352
rect 16669 20349 16681 20352
rect 16715 20380 16727 20383
rect 17313 20383 17371 20389
rect 17313 20380 17325 20383
rect 16715 20352 17325 20380
rect 16715 20349 16727 20352
rect 16669 20343 16727 20349
rect 17313 20349 17325 20352
rect 17359 20349 17371 20383
rect 17313 20343 17371 20349
rect 18969 20383 19027 20389
rect 18969 20349 18981 20383
rect 19015 20380 19027 20383
rect 19328 20383 19386 20389
rect 19328 20380 19340 20383
rect 19015 20352 19340 20380
rect 19015 20349 19027 20352
rect 18969 20343 19027 20349
rect 19328 20349 19340 20352
rect 19374 20380 19386 20383
rect 20622 20380 20628 20392
rect 19374 20352 20628 20380
rect 19374 20349 19386 20352
rect 19328 20343 19386 20349
rect 20622 20340 20628 20352
rect 20680 20340 20686 20392
rect 23382 20380 23388 20392
rect 21560 20352 23388 20380
rect 12897 20315 12955 20321
rect 12897 20312 12909 20315
rect 11664 20284 12112 20312
rect 12176 20284 12909 20312
rect 11664 20272 11670 20284
rect 4341 20247 4399 20253
rect 4341 20244 4353 20247
rect 3660 20216 4353 20244
rect 3660 20204 3666 20216
rect 4341 20213 4353 20216
rect 4387 20213 4399 20247
rect 4341 20207 4399 20213
rect 8018 20204 8024 20256
rect 8076 20244 8082 20256
rect 8846 20244 8852 20256
rect 8076 20216 8852 20244
rect 8076 20204 8082 20216
rect 8846 20204 8852 20216
rect 8904 20244 8910 20256
rect 9033 20247 9091 20253
rect 9033 20244 9045 20247
rect 8904 20216 9045 20244
rect 8904 20204 8910 20216
rect 9033 20213 9045 20216
rect 9079 20213 9091 20247
rect 9398 20244 9404 20256
rect 9359 20216 9404 20244
rect 9033 20207 9091 20213
rect 9398 20204 9404 20216
rect 9456 20204 9462 20256
rect 12084 20253 12112 20284
rect 12897 20281 12909 20284
rect 12943 20281 12955 20315
rect 12897 20275 12955 20281
rect 13814 20272 13820 20324
rect 13872 20312 13878 20324
rect 14108 20312 14136 20340
rect 15378 20312 15384 20324
rect 13872 20284 15384 20312
rect 13872 20272 13878 20284
rect 15378 20272 15384 20284
rect 15436 20312 15442 20324
rect 15654 20312 15660 20324
rect 15436 20284 15660 20312
rect 15436 20272 15442 20284
rect 15654 20272 15660 20284
rect 15712 20272 15718 20324
rect 16761 20315 16819 20321
rect 16761 20281 16773 20315
rect 16807 20312 16819 20315
rect 16942 20312 16948 20324
rect 16807 20284 16948 20312
rect 16807 20281 16819 20284
rect 16761 20275 16819 20281
rect 16942 20272 16948 20284
rect 17000 20272 17006 20324
rect 17865 20315 17923 20321
rect 17865 20281 17877 20315
rect 17911 20312 17923 20315
rect 19150 20312 19156 20324
rect 17911 20284 19156 20312
rect 17911 20281 17923 20284
rect 17865 20275 17923 20281
rect 19150 20272 19156 20284
rect 19208 20312 19214 20324
rect 21560 20321 21588 20352
rect 23382 20340 23388 20352
rect 23440 20380 23446 20392
rect 23658 20380 23664 20392
rect 23440 20352 23664 20380
rect 23440 20340 23446 20352
rect 23658 20340 23664 20352
rect 23716 20340 23722 20392
rect 23750 20340 23756 20392
rect 23808 20380 23814 20392
rect 24029 20383 24087 20389
rect 24029 20380 24041 20383
rect 23808 20352 24041 20380
rect 23808 20340 23814 20352
rect 24029 20349 24041 20352
rect 24075 20349 24087 20383
rect 24136 20380 24164 20408
rect 24673 20383 24731 20389
rect 24673 20380 24685 20383
rect 24136 20352 24685 20380
rect 24029 20343 24087 20349
rect 24673 20349 24685 20352
rect 24719 20349 24731 20383
rect 24673 20343 24731 20349
rect 25225 20383 25283 20389
rect 25225 20349 25237 20383
rect 25271 20380 25283 20383
rect 25314 20380 25320 20392
rect 25271 20352 25320 20380
rect 25271 20349 25283 20352
rect 25225 20343 25283 20349
rect 25314 20340 25320 20352
rect 25372 20380 25378 20392
rect 25961 20383 26019 20389
rect 25961 20380 25973 20383
rect 25372 20352 25973 20380
rect 25372 20340 25378 20352
rect 25961 20349 25973 20352
rect 26007 20349 26019 20383
rect 25961 20343 26019 20349
rect 20809 20315 20867 20321
rect 19208 20284 20484 20312
rect 19208 20272 19214 20284
rect 20456 20256 20484 20284
rect 20809 20281 20821 20315
rect 20855 20312 20867 20315
rect 21514 20315 21588 20321
rect 21514 20312 21526 20315
rect 20855 20284 21526 20312
rect 20855 20281 20867 20284
rect 20809 20275 20867 20281
rect 21514 20281 21526 20284
rect 21560 20284 21588 20315
rect 21560 20281 21572 20284
rect 21514 20275 21572 20281
rect 25130 20272 25136 20324
rect 25188 20312 25194 20324
rect 26234 20312 26240 20324
rect 25188 20284 26240 20312
rect 25188 20272 25194 20284
rect 26234 20272 26240 20284
rect 26292 20272 26298 20324
rect 12069 20247 12127 20253
rect 12069 20213 12081 20247
rect 12115 20244 12127 20247
rect 12158 20244 12164 20256
rect 12115 20216 12164 20244
rect 12115 20213 12127 20216
rect 12069 20207 12127 20213
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 12434 20204 12440 20256
rect 12492 20244 12498 20256
rect 13446 20244 13452 20256
rect 12492 20216 12537 20244
rect 13407 20216 13452 20244
rect 12492 20204 12498 20216
rect 13446 20204 13452 20216
rect 13504 20204 13510 20256
rect 15841 20247 15899 20253
rect 15841 20213 15853 20247
rect 15887 20244 15899 20247
rect 16114 20244 16120 20256
rect 15887 20216 16120 20244
rect 15887 20213 15899 20216
rect 15841 20207 15899 20213
rect 16114 20204 16120 20216
rect 16172 20204 16178 20256
rect 18046 20244 18052 20256
rect 18007 20216 18052 20244
rect 18046 20204 18052 20216
rect 18104 20204 18110 20256
rect 18414 20204 18420 20256
rect 18472 20244 18478 20256
rect 18509 20247 18567 20253
rect 18509 20244 18521 20247
rect 18472 20216 18521 20244
rect 18472 20204 18478 20216
rect 18509 20213 18521 20216
rect 18555 20213 18567 20247
rect 20438 20244 20444 20256
rect 20399 20216 20444 20244
rect 18509 20207 18567 20213
rect 20438 20204 20444 20216
rect 20496 20204 20502 20256
rect 21082 20244 21088 20256
rect 21043 20216 21088 20244
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 21818 20204 21824 20256
rect 21876 20244 21882 20256
rect 22186 20244 22192 20256
rect 21876 20216 22192 20244
rect 21876 20204 21882 20216
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 22370 20204 22376 20256
rect 22428 20244 22434 20256
rect 22646 20244 22652 20256
rect 22428 20216 22652 20244
rect 22428 20204 22434 20216
rect 22646 20204 22652 20216
rect 22704 20204 22710 20256
rect 23014 20244 23020 20256
rect 22975 20216 23020 20244
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 23477 20247 23535 20253
rect 23477 20213 23489 20247
rect 23523 20244 23535 20247
rect 23566 20244 23572 20256
rect 23523 20216 23572 20244
rect 23523 20213 23535 20216
rect 23477 20207 23535 20213
rect 23566 20204 23572 20216
rect 23624 20244 23630 20256
rect 23934 20244 23940 20256
rect 23624 20216 23940 20244
rect 23624 20204 23630 20216
rect 23934 20204 23940 20216
rect 23992 20244 23998 20256
rect 24302 20244 24308 20256
rect 23992 20216 24308 20244
rect 23992 20204 23998 20216
rect 24302 20204 24308 20216
rect 24360 20204 24366 20256
rect 25038 20244 25044 20256
rect 24999 20216 25044 20244
rect 25038 20204 25044 20216
rect 25096 20204 25102 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1397 20043 1455 20049
rect 1397 20009 1409 20043
rect 1443 20040 1455 20043
rect 2866 20040 2872 20052
rect 1443 20012 2872 20040
rect 1443 20009 1455 20012
rect 1397 20003 1455 20009
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 3510 20040 3516 20052
rect 3471 20012 3516 20040
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 3881 20043 3939 20049
rect 3881 20009 3893 20043
rect 3927 20040 3939 20043
rect 4062 20040 4068 20052
rect 3927 20012 4068 20040
rect 3927 20009 3939 20012
rect 3881 20003 3939 20009
rect 2317 19975 2375 19981
rect 2317 19941 2329 19975
rect 2363 19972 2375 19975
rect 3142 19972 3148 19984
rect 2363 19944 3148 19972
rect 2363 19941 2375 19944
rect 2317 19935 2375 19941
rect 2774 19864 2780 19916
rect 2832 19904 2838 19916
rect 2832 19876 2877 19904
rect 2832 19864 2838 19876
rect 2866 19836 2872 19848
rect 2827 19808 2872 19836
rect 2866 19796 2872 19808
rect 2924 19796 2930 19848
rect 3068 19845 3096 19944
rect 3142 19932 3148 19944
rect 3200 19932 3206 19984
rect 3053 19839 3111 19845
rect 3053 19805 3065 19839
rect 3099 19805 3111 19839
rect 3053 19799 3111 19805
rect 2409 19771 2467 19777
rect 2409 19737 2421 19771
rect 2455 19768 2467 19771
rect 3896 19768 3924 20003
rect 4062 20000 4068 20012
rect 4120 20000 4126 20052
rect 4341 20043 4399 20049
rect 4341 20009 4353 20043
rect 4387 20040 4399 20043
rect 4614 20040 4620 20052
rect 4387 20012 4620 20040
rect 4387 20009 4399 20012
rect 4341 20003 4399 20009
rect 4614 20000 4620 20012
rect 4672 20000 4678 20052
rect 6549 20043 6607 20049
rect 6549 20009 6561 20043
rect 6595 20040 6607 20043
rect 6730 20040 6736 20052
rect 6595 20012 6736 20040
rect 6595 20009 6607 20012
rect 6549 20003 6607 20009
rect 4430 19932 4436 19984
rect 4488 19972 4494 19984
rect 4976 19975 5034 19981
rect 4976 19972 4988 19975
rect 4488 19944 4988 19972
rect 4488 19932 4494 19944
rect 4976 19941 4988 19944
rect 5022 19972 5034 19975
rect 6564 19972 6592 20003
rect 6730 20000 6736 20012
rect 6788 20000 6794 20052
rect 6914 20000 6920 20052
rect 6972 20040 6978 20052
rect 7377 20043 7435 20049
rect 7377 20040 7389 20043
rect 6972 20012 7389 20040
rect 6972 20000 6978 20012
rect 7377 20009 7389 20012
rect 7423 20040 7435 20043
rect 7834 20040 7840 20052
rect 7423 20012 7840 20040
rect 7423 20009 7435 20012
rect 7377 20003 7435 20009
rect 7834 20000 7840 20012
rect 7892 20000 7898 20052
rect 8113 20043 8171 20049
rect 8113 20009 8125 20043
rect 8159 20040 8171 20043
rect 8202 20040 8208 20052
rect 8159 20012 8208 20040
rect 8159 20009 8171 20012
rect 8113 20003 8171 20009
rect 8202 20000 8208 20012
rect 8260 20000 8266 20052
rect 8481 20043 8539 20049
rect 8481 20009 8493 20043
rect 8527 20040 8539 20043
rect 8662 20040 8668 20052
rect 8527 20012 8668 20040
rect 8527 20009 8539 20012
rect 8481 20003 8539 20009
rect 8662 20000 8668 20012
rect 8720 20000 8726 20052
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 10321 20043 10379 20049
rect 10321 20040 10333 20043
rect 10192 20012 10333 20040
rect 10192 20000 10198 20012
rect 10321 20009 10333 20012
rect 10367 20009 10379 20043
rect 10778 20040 10784 20052
rect 10739 20012 10784 20040
rect 10321 20003 10379 20009
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 11054 20000 11060 20052
rect 11112 20040 11118 20052
rect 11885 20043 11943 20049
rect 11885 20040 11897 20043
rect 11112 20012 11897 20040
rect 11112 20000 11118 20012
rect 11885 20009 11897 20012
rect 11931 20009 11943 20043
rect 11885 20003 11943 20009
rect 12250 20000 12256 20052
rect 12308 20040 12314 20052
rect 12345 20043 12403 20049
rect 12345 20040 12357 20043
rect 12308 20012 12357 20040
rect 12308 20000 12314 20012
rect 12345 20009 12357 20012
rect 12391 20009 12403 20043
rect 12345 20003 12403 20009
rect 12618 20000 12624 20052
rect 12676 20040 12682 20052
rect 12897 20043 12955 20049
rect 12897 20040 12909 20043
rect 12676 20012 12909 20040
rect 12676 20000 12682 20012
rect 12897 20009 12909 20012
rect 12943 20009 12955 20043
rect 12897 20003 12955 20009
rect 13449 20043 13507 20049
rect 13449 20009 13461 20043
rect 13495 20040 13507 20043
rect 13722 20040 13728 20052
rect 13495 20012 13728 20040
rect 13495 20009 13507 20012
rect 13449 20003 13507 20009
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 14553 20043 14611 20049
rect 14553 20009 14565 20043
rect 14599 20040 14611 20043
rect 14642 20040 14648 20052
rect 14599 20012 14648 20040
rect 14599 20009 14611 20012
rect 14553 20003 14611 20009
rect 14642 20000 14648 20012
rect 14700 20000 14706 20052
rect 16666 20040 16672 20052
rect 16627 20012 16672 20040
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 17770 20000 17776 20052
rect 17828 20040 17834 20052
rect 17865 20043 17923 20049
rect 17865 20040 17877 20043
rect 17828 20012 17877 20040
rect 17828 20000 17834 20012
rect 17865 20009 17877 20012
rect 17911 20040 17923 20043
rect 18230 20040 18236 20052
rect 17911 20012 18236 20040
rect 17911 20009 17923 20012
rect 17865 20003 17923 20009
rect 18230 20000 18236 20012
rect 18288 20000 18294 20052
rect 19518 20000 19524 20052
rect 19576 20040 19582 20052
rect 20901 20043 20959 20049
rect 20901 20040 20913 20043
rect 19576 20012 20913 20040
rect 19576 20000 19582 20012
rect 20901 20009 20913 20012
rect 20947 20009 20959 20043
rect 20901 20003 20959 20009
rect 21082 20000 21088 20052
rect 21140 20040 21146 20052
rect 21818 20040 21824 20052
rect 21140 20012 21824 20040
rect 21140 20000 21146 20012
rect 21818 20000 21824 20012
rect 21876 20000 21882 20052
rect 22373 20043 22431 20049
rect 22373 20009 22385 20043
rect 22419 20040 22431 20043
rect 23014 20040 23020 20052
rect 22419 20012 23020 20040
rect 22419 20009 22431 20012
rect 22373 20003 22431 20009
rect 23014 20000 23020 20012
rect 23072 20000 23078 20052
rect 23750 20000 23756 20052
rect 23808 20040 23814 20052
rect 24305 20043 24363 20049
rect 24305 20040 24317 20043
rect 23808 20012 24317 20040
rect 23808 20000 23814 20012
rect 24305 20009 24317 20012
rect 24351 20009 24363 20043
rect 24854 20040 24860 20052
rect 24815 20012 24860 20040
rect 24305 20003 24363 20009
rect 24854 20000 24860 20012
rect 24912 20000 24918 20052
rect 5022 19944 6592 19972
rect 9493 19975 9551 19981
rect 5022 19941 5034 19944
rect 4976 19935 5034 19941
rect 9493 19941 9505 19975
rect 9539 19972 9551 19975
rect 10796 19972 10824 20000
rect 9539 19944 10824 19972
rect 9539 19941 9551 19944
rect 9493 19935 9551 19941
rect 13354 19932 13360 19984
rect 13412 19972 13418 19984
rect 13909 19975 13967 19981
rect 13909 19972 13921 19975
rect 13412 19944 13921 19972
rect 13412 19932 13418 19944
rect 13909 19941 13921 19944
rect 13955 19941 13967 19975
rect 16298 19972 16304 19984
rect 13909 19935 13967 19941
rect 14108 19944 16304 19972
rect 14108 19916 14136 19944
rect 16298 19932 16304 19944
rect 16356 19932 16362 19984
rect 18414 19932 18420 19984
rect 18472 19972 18478 19984
rect 20162 19972 20168 19984
rect 18472 19944 20168 19972
rect 18472 19932 18478 19944
rect 20162 19932 20168 19944
rect 20220 19972 20226 19984
rect 20257 19975 20315 19981
rect 20257 19972 20269 19975
rect 20220 19944 20269 19972
rect 20220 19932 20226 19944
rect 20257 19941 20269 19944
rect 20303 19941 20315 19975
rect 22002 19972 22008 19984
rect 21963 19944 22008 19972
rect 20257 19935 20315 19941
rect 22002 19932 22008 19944
rect 22060 19932 22066 19984
rect 24673 19975 24731 19981
rect 24673 19972 24685 19975
rect 22756 19944 24685 19972
rect 22756 19916 22784 19944
rect 24673 19941 24685 19944
rect 24719 19972 24731 19975
rect 24762 19972 24768 19984
rect 24719 19944 24768 19972
rect 24719 19941 24731 19944
rect 24673 19935 24731 19941
rect 24762 19932 24768 19944
rect 24820 19972 24826 19984
rect 25038 19972 25044 19984
rect 24820 19944 25044 19972
rect 24820 19932 24826 19944
rect 25038 19932 25044 19944
rect 25096 19932 25102 19984
rect 4522 19864 4528 19916
rect 4580 19904 4586 19916
rect 4709 19907 4767 19913
rect 4709 19904 4721 19907
rect 4580 19876 4721 19904
rect 4580 19864 4586 19876
rect 4709 19873 4721 19876
rect 4755 19873 4767 19907
rect 7282 19904 7288 19916
rect 7243 19876 7288 19904
rect 4709 19867 4767 19873
rect 7282 19864 7288 19876
rect 7340 19864 7346 19916
rect 9858 19864 9864 19916
rect 9916 19904 9922 19916
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 9916 19876 10149 19904
rect 9916 19864 9922 19876
rect 10137 19873 10149 19876
rect 10183 19873 10195 19907
rect 10137 19867 10195 19873
rect 10689 19907 10747 19913
rect 10689 19873 10701 19907
rect 10735 19904 10747 19907
rect 10962 19904 10968 19916
rect 10735 19876 10968 19904
rect 10735 19873 10747 19876
rect 10689 19867 10747 19873
rect 10962 19864 10968 19876
rect 11020 19864 11026 19916
rect 12250 19904 12256 19916
rect 12211 19876 12256 19904
rect 12250 19864 12256 19876
rect 12308 19864 12314 19916
rect 13817 19907 13875 19913
rect 13817 19873 13829 19907
rect 13863 19904 13875 19907
rect 14090 19904 14096 19916
rect 13863 19876 14096 19904
rect 13863 19873 13875 19876
rect 13817 19867 13875 19873
rect 14090 19864 14096 19876
rect 14148 19864 14154 19916
rect 15289 19907 15347 19913
rect 15289 19873 15301 19907
rect 15335 19904 15347 19907
rect 15378 19904 15384 19916
rect 15335 19876 15384 19904
rect 15335 19873 15347 19876
rect 15289 19867 15347 19873
rect 15378 19864 15384 19876
rect 15436 19864 15442 19916
rect 15556 19907 15614 19913
rect 15556 19873 15568 19907
rect 15602 19904 15614 19907
rect 15838 19904 15844 19916
rect 15602 19876 15844 19904
rect 15602 19873 15614 19876
rect 15556 19867 15614 19873
rect 15838 19864 15844 19876
rect 15896 19864 15902 19916
rect 17862 19864 17868 19916
rect 17920 19904 17926 19916
rect 17957 19907 18015 19913
rect 17957 19904 17969 19907
rect 17920 19876 17969 19904
rect 17920 19864 17926 19876
rect 17957 19873 17969 19876
rect 18003 19873 18015 19907
rect 17957 19867 18015 19873
rect 19518 19864 19524 19916
rect 19576 19904 19582 19916
rect 19613 19907 19671 19913
rect 19613 19904 19625 19907
rect 19576 19876 19625 19904
rect 19576 19864 19582 19876
rect 19613 19873 19625 19876
rect 19659 19873 19671 19907
rect 21266 19904 21272 19916
rect 21227 19876 21272 19904
rect 19613 19867 19671 19873
rect 21266 19864 21272 19876
rect 21324 19864 21330 19916
rect 21361 19907 21419 19913
rect 21361 19873 21373 19907
rect 21407 19904 21419 19907
rect 22370 19904 22376 19916
rect 21407 19876 22376 19904
rect 21407 19873 21419 19876
rect 21361 19867 21419 19873
rect 22370 19864 22376 19876
rect 22428 19864 22434 19916
rect 22649 19907 22707 19913
rect 22649 19873 22661 19907
rect 22695 19904 22707 19907
rect 22738 19904 22744 19916
rect 22695 19876 22744 19904
rect 22695 19873 22707 19876
rect 22649 19867 22707 19873
rect 22738 19864 22744 19876
rect 22796 19864 22802 19916
rect 22922 19913 22928 19916
rect 22916 19867 22928 19913
rect 22980 19904 22986 19916
rect 25225 19907 25283 19913
rect 22980 19876 23016 19904
rect 22922 19864 22928 19867
rect 22980 19864 22986 19876
rect 25225 19873 25237 19907
rect 25271 19904 25283 19907
rect 25682 19904 25688 19916
rect 25271 19876 25688 19904
rect 25271 19873 25283 19876
rect 25225 19867 25283 19873
rect 25682 19864 25688 19876
rect 25740 19864 25746 19916
rect 6270 19836 6276 19848
rect 6104 19808 6276 19836
rect 6104 19777 6132 19808
rect 6270 19796 6276 19808
rect 6328 19836 6334 19848
rect 7469 19839 7527 19845
rect 7469 19836 7481 19839
rect 6328 19808 7481 19836
rect 6328 19796 6334 19808
rect 7469 19805 7481 19808
rect 7515 19805 7527 19839
rect 8570 19836 8576 19848
rect 8531 19808 8576 19836
rect 7469 19799 7527 19805
rect 8570 19796 8576 19808
rect 8628 19796 8634 19848
rect 10042 19796 10048 19848
rect 10100 19836 10106 19848
rect 10873 19839 10931 19845
rect 10873 19836 10885 19839
rect 10100 19808 10885 19836
rect 10100 19796 10106 19808
rect 10873 19805 10885 19808
rect 10919 19805 10931 19839
rect 10873 19799 10931 19805
rect 11974 19796 11980 19848
rect 12032 19836 12038 19848
rect 12529 19839 12587 19845
rect 12529 19836 12541 19839
rect 12032 19808 12541 19836
rect 12032 19796 12038 19808
rect 12529 19805 12541 19808
rect 12575 19836 12587 19839
rect 12986 19836 12992 19848
rect 12575 19808 12992 19836
rect 12575 19805 12587 19808
rect 12529 19799 12587 19805
rect 12986 19796 12992 19808
rect 13044 19836 13050 19848
rect 13265 19839 13323 19845
rect 13265 19836 13277 19839
rect 13044 19808 13277 19836
rect 13044 19796 13050 19808
rect 13265 19805 13277 19808
rect 13311 19805 13323 19839
rect 13998 19836 14004 19848
rect 13959 19808 14004 19836
rect 13265 19799 13323 19805
rect 13998 19796 14004 19808
rect 14056 19796 14062 19848
rect 18049 19839 18107 19845
rect 18049 19805 18061 19839
rect 18095 19805 18107 19839
rect 18049 19799 18107 19805
rect 2455 19740 3924 19768
rect 6089 19771 6147 19777
rect 2455 19737 2467 19740
rect 2409 19731 2467 19737
rect 6089 19737 6101 19771
rect 6135 19737 6147 19771
rect 6914 19768 6920 19780
rect 6875 19740 6920 19768
rect 6089 19731 6147 19737
rect 6914 19728 6920 19740
rect 6972 19728 6978 19780
rect 16758 19728 16764 19780
rect 16816 19768 16822 19780
rect 17037 19771 17095 19777
rect 17037 19768 17049 19771
rect 16816 19740 17049 19768
rect 16816 19728 16822 19740
rect 17037 19737 17049 19740
rect 17083 19768 17095 19771
rect 17497 19771 17555 19777
rect 17497 19768 17509 19771
rect 17083 19740 17509 19768
rect 17083 19737 17095 19740
rect 17037 19731 17095 19737
rect 17497 19737 17509 19740
rect 17543 19737 17555 19771
rect 18064 19768 18092 19799
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 19705 19839 19763 19845
rect 19705 19836 19717 19839
rect 19392 19808 19717 19836
rect 19392 19796 19398 19808
rect 19705 19805 19717 19808
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 19797 19839 19855 19845
rect 19797 19805 19809 19839
rect 19843 19805 19855 19839
rect 19797 19799 19855 19805
rect 17497 19731 17555 19737
rect 17880 19740 18092 19768
rect 19153 19771 19211 19777
rect 1854 19700 1860 19712
rect 1815 19672 1860 19700
rect 1854 19660 1860 19672
rect 1912 19660 1918 19712
rect 2866 19660 2872 19712
rect 2924 19700 2930 19712
rect 3694 19700 3700 19712
rect 2924 19672 3700 19700
rect 2924 19660 2930 19672
rect 3694 19660 3700 19672
rect 3752 19700 3758 19712
rect 7190 19700 7196 19712
rect 3752 19672 7196 19700
rect 3752 19660 3758 19672
rect 7190 19660 7196 19672
rect 7248 19660 7254 19712
rect 8938 19660 8944 19712
rect 8996 19700 9002 19712
rect 9125 19703 9183 19709
rect 9125 19700 9137 19703
rect 8996 19672 9137 19700
rect 8996 19660 9002 19672
rect 9125 19669 9137 19672
rect 9171 19700 9183 19703
rect 9398 19700 9404 19712
rect 9171 19672 9404 19700
rect 9171 19669 9183 19672
rect 9125 19663 9183 19669
rect 9398 19660 9404 19672
rect 9456 19700 9462 19712
rect 11422 19700 11428 19712
rect 9456 19672 11428 19700
rect 9456 19660 9462 19672
rect 11422 19660 11428 19672
rect 11480 19700 11486 19712
rect 11701 19703 11759 19709
rect 11701 19700 11713 19703
rect 11480 19672 11713 19700
rect 11480 19660 11486 19672
rect 11701 19669 11713 19672
rect 11747 19669 11759 19703
rect 11701 19663 11759 19669
rect 14642 19660 14648 19712
rect 14700 19700 14706 19712
rect 15013 19703 15071 19709
rect 15013 19700 15025 19703
rect 14700 19672 15025 19700
rect 14700 19660 14706 19672
rect 15013 19669 15025 19672
rect 15059 19700 15071 19703
rect 15470 19700 15476 19712
rect 15059 19672 15476 19700
rect 15059 19669 15071 19672
rect 15013 19663 15071 19669
rect 15470 19660 15476 19672
rect 15528 19660 15534 19712
rect 17405 19703 17463 19709
rect 17405 19669 17417 19703
rect 17451 19700 17463 19703
rect 17770 19700 17776 19712
rect 17451 19672 17776 19700
rect 17451 19669 17463 19672
rect 17405 19663 17463 19669
rect 17770 19660 17776 19672
rect 17828 19700 17834 19712
rect 17880 19700 17908 19740
rect 19153 19737 19165 19771
rect 19199 19768 19211 19771
rect 19812 19768 19840 19799
rect 20530 19796 20536 19848
rect 20588 19836 20594 19848
rect 20898 19836 20904 19848
rect 20588 19808 20904 19836
rect 20588 19796 20594 19808
rect 20898 19796 20904 19808
rect 20956 19836 20962 19848
rect 21453 19839 21511 19845
rect 21453 19836 21465 19839
rect 20956 19808 21465 19836
rect 20956 19796 20962 19808
rect 21453 19805 21465 19808
rect 21499 19805 21511 19839
rect 25314 19836 25320 19848
rect 25275 19808 25320 19836
rect 21453 19799 21511 19805
rect 25314 19796 25320 19808
rect 25372 19796 25378 19848
rect 25501 19839 25559 19845
rect 25501 19805 25513 19839
rect 25547 19836 25559 19839
rect 25590 19836 25596 19848
rect 25547 19808 25596 19836
rect 25547 19805 25559 19808
rect 25501 19799 25559 19805
rect 25590 19796 25596 19808
rect 25648 19796 25654 19848
rect 19978 19768 19984 19780
rect 19199 19740 19984 19768
rect 19199 19737 19211 19740
rect 19153 19731 19211 19737
rect 19978 19728 19984 19740
rect 20036 19728 20042 19780
rect 23658 19728 23664 19780
rect 23716 19768 23722 19780
rect 24029 19771 24087 19777
rect 24029 19768 24041 19771
rect 23716 19740 24041 19768
rect 23716 19728 23722 19740
rect 24029 19737 24041 19740
rect 24075 19737 24087 19771
rect 24029 19731 24087 19737
rect 17828 19672 17908 19700
rect 17828 19660 17834 19672
rect 18322 19660 18328 19712
rect 18380 19700 18386 19712
rect 18509 19703 18567 19709
rect 18509 19700 18521 19703
rect 18380 19672 18521 19700
rect 18380 19660 18386 19672
rect 18509 19669 18521 19672
rect 18555 19669 18567 19703
rect 19242 19700 19248 19712
rect 19203 19672 19248 19700
rect 18509 19663 18567 19669
rect 19242 19660 19248 19672
rect 19300 19660 19306 19712
rect 20438 19660 20444 19712
rect 20496 19700 20502 19712
rect 20717 19703 20775 19709
rect 20717 19700 20729 19703
rect 20496 19672 20729 19700
rect 20496 19660 20502 19672
rect 20717 19669 20729 19672
rect 20763 19700 20775 19703
rect 21910 19700 21916 19712
rect 20763 19672 21916 19700
rect 20763 19669 20775 19672
rect 20717 19663 20775 19669
rect 21910 19660 21916 19672
rect 21968 19660 21974 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2774 19456 2780 19508
rect 2832 19496 2838 19508
rect 3970 19496 3976 19508
rect 2832 19468 3976 19496
rect 2832 19456 2838 19468
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 4430 19496 4436 19508
rect 4391 19468 4436 19496
rect 4430 19456 4436 19468
rect 4488 19456 4494 19508
rect 6822 19496 6828 19508
rect 6735 19468 6828 19496
rect 6822 19456 6828 19468
rect 6880 19496 6886 19508
rect 7282 19496 7288 19508
rect 6880 19468 7288 19496
rect 6880 19456 6886 19468
rect 7282 19456 7288 19468
rect 7340 19456 7346 19508
rect 9122 19456 9128 19508
rect 9180 19496 9186 19508
rect 9677 19499 9735 19505
rect 9180 19468 9352 19496
rect 9180 19456 9186 19468
rect 9324 19440 9352 19468
rect 9677 19465 9689 19499
rect 9723 19496 9735 19499
rect 10042 19496 10048 19508
rect 9723 19468 10048 19496
rect 9723 19465 9735 19468
rect 9677 19459 9735 19465
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 11609 19499 11667 19505
rect 11609 19465 11621 19499
rect 11655 19496 11667 19499
rect 12250 19496 12256 19508
rect 11655 19468 12256 19496
rect 11655 19465 11667 19468
rect 11609 19459 11667 19465
rect 12250 19456 12256 19468
rect 12308 19456 12314 19508
rect 13814 19496 13820 19508
rect 13556 19468 13820 19496
rect 2501 19431 2559 19437
rect 2501 19397 2513 19431
rect 2547 19428 2559 19431
rect 2866 19428 2872 19440
rect 2547 19400 2872 19428
rect 2547 19397 2559 19400
rect 2501 19391 2559 19397
rect 2866 19388 2872 19400
rect 2924 19388 2930 19440
rect 3142 19388 3148 19440
rect 3200 19428 3206 19440
rect 4065 19431 4123 19437
rect 4065 19428 4077 19431
rect 3200 19400 4077 19428
rect 3200 19388 3206 19400
rect 4065 19397 4077 19400
rect 4111 19397 4123 19431
rect 4065 19391 4123 19397
rect 9306 19388 9312 19440
rect 9364 19388 9370 19440
rect 11977 19431 12035 19437
rect 11977 19397 11989 19431
rect 12023 19428 12035 19431
rect 12158 19428 12164 19440
rect 12023 19400 12164 19428
rect 12023 19397 12035 19400
rect 11977 19391 12035 19397
rect 12158 19388 12164 19400
rect 12216 19388 12222 19440
rect 1854 19320 1860 19372
rect 1912 19360 1918 19372
rect 1949 19363 2007 19369
rect 1949 19360 1961 19363
rect 1912 19332 1961 19360
rect 1912 19320 1918 19332
rect 1949 19329 1961 19332
rect 1995 19329 2007 19363
rect 3510 19360 3516 19372
rect 3471 19332 3516 19360
rect 1949 19323 2007 19329
rect 3510 19320 3516 19332
rect 3568 19320 3574 19372
rect 4522 19360 4528 19372
rect 4483 19332 4528 19360
rect 4522 19320 4528 19332
rect 4580 19320 4586 19372
rect 6730 19320 6736 19372
rect 6788 19360 6794 19372
rect 7377 19363 7435 19369
rect 7377 19360 7389 19363
rect 6788 19332 7389 19360
rect 6788 19320 6794 19332
rect 7377 19329 7389 19332
rect 7423 19360 7435 19363
rect 7466 19360 7472 19372
rect 7423 19332 7472 19360
rect 7423 19329 7435 19332
rect 7377 19323 7435 19329
rect 7466 19320 7472 19332
rect 7524 19320 7530 19372
rect 9122 19360 9128 19372
rect 9083 19332 9128 19360
rect 9122 19320 9128 19332
rect 9180 19320 9186 19372
rect 9674 19320 9680 19372
rect 9732 19360 9738 19372
rect 10689 19363 10747 19369
rect 10689 19360 10701 19363
rect 9732 19332 10701 19360
rect 9732 19320 9738 19332
rect 10689 19329 10701 19332
rect 10735 19360 10747 19363
rect 10735 19332 11008 19360
rect 10735 19329 10747 19332
rect 10689 19323 10747 19329
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 2222 19292 2228 19304
rect 1811 19264 2228 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 3329 19295 3387 19301
rect 3329 19261 3341 19295
rect 3375 19292 3387 19295
rect 3786 19292 3792 19304
rect 3375 19264 3792 19292
rect 3375 19261 3387 19264
rect 3329 19255 3387 19261
rect 3786 19252 3792 19264
rect 3844 19252 3850 19304
rect 8113 19295 8171 19301
rect 8113 19261 8125 19295
rect 8159 19292 8171 19295
rect 8662 19292 8668 19304
rect 8159 19264 8668 19292
rect 8159 19261 8171 19264
rect 8113 19255 8171 19261
rect 8662 19252 8668 19264
rect 8720 19252 8726 19304
rect 9950 19292 9956 19304
rect 9911 19264 9956 19292
rect 9950 19252 9956 19264
rect 10008 19292 10014 19304
rect 10597 19295 10655 19301
rect 10597 19292 10609 19295
rect 10008 19264 10609 19292
rect 10008 19252 10014 19264
rect 10597 19261 10609 19264
rect 10643 19261 10655 19295
rect 10980 19292 11008 19332
rect 11330 19292 11336 19304
rect 10980 19264 11336 19292
rect 10597 19255 10655 19261
rect 11330 19252 11336 19264
rect 11388 19252 11394 19304
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 12526 19292 12532 19304
rect 12483 19264 12532 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12526 19252 12532 19264
rect 12584 19292 12590 19304
rect 13078 19292 13084 19304
rect 12584 19264 13084 19292
rect 12584 19252 12590 19264
rect 13078 19252 13084 19264
rect 13136 19252 13142 19304
rect 13354 19292 13360 19304
rect 13315 19264 13360 19292
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 13556 19301 13584 19468
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 17586 19496 17592 19508
rect 17499 19468 17592 19496
rect 17586 19456 17592 19468
rect 17644 19496 17650 19508
rect 17862 19496 17868 19508
rect 17644 19468 17868 19496
rect 17644 19456 17650 19468
rect 17862 19456 17868 19468
rect 17920 19456 17926 19508
rect 19061 19499 19119 19505
rect 19061 19465 19073 19499
rect 19107 19496 19119 19499
rect 19334 19496 19340 19508
rect 19107 19468 19340 19496
rect 19107 19465 19119 19468
rect 19061 19459 19119 19465
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 20533 19499 20591 19505
rect 20533 19465 20545 19499
rect 20579 19496 20591 19499
rect 20622 19496 20628 19508
rect 20579 19468 20628 19496
rect 20579 19465 20591 19468
rect 20533 19459 20591 19465
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 20901 19499 20959 19505
rect 20901 19465 20913 19499
rect 20947 19496 20959 19499
rect 21266 19496 21272 19508
rect 20947 19468 21272 19496
rect 20947 19465 20959 19468
rect 20901 19459 20959 19465
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 22833 19499 22891 19505
rect 22833 19465 22845 19499
rect 22879 19496 22891 19499
rect 22922 19496 22928 19508
rect 22879 19468 22928 19496
rect 22879 19465 22891 19468
rect 22833 19459 22891 19465
rect 22922 19456 22928 19468
rect 22980 19456 22986 19508
rect 17494 19388 17500 19440
rect 17552 19428 17558 19440
rect 17954 19428 17960 19440
rect 17552 19400 17960 19428
rect 17552 19388 17558 19400
rect 17954 19388 17960 19400
rect 18012 19388 18018 19440
rect 16942 19360 16948 19372
rect 16903 19332 16948 19360
rect 16942 19320 16948 19332
rect 17000 19320 17006 19372
rect 21082 19360 21088 19372
rect 20548 19332 21088 19360
rect 20548 19304 20576 19332
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 21910 19360 21916 19372
rect 21871 19332 21916 19360
rect 21910 19320 21916 19332
rect 21968 19320 21974 19372
rect 13541 19295 13599 19301
rect 13541 19261 13553 19295
rect 13587 19261 13599 19295
rect 13541 19255 13599 19261
rect 15381 19295 15439 19301
rect 15381 19261 15393 19295
rect 15427 19292 15439 19295
rect 15838 19292 15844 19304
rect 15427 19264 15844 19292
rect 15427 19261 15439 19264
rect 15381 19255 15439 19261
rect 2866 19224 2872 19236
rect 1412 19196 2872 19224
rect 1412 19165 1440 19196
rect 2866 19184 2872 19196
rect 2924 19184 2930 19236
rect 3418 19224 3424 19236
rect 3379 19196 3424 19224
rect 3418 19184 3424 19196
rect 3476 19184 3482 19236
rect 4798 19233 4804 19236
rect 4792 19224 4804 19233
rect 4759 19196 4804 19224
rect 4792 19187 4804 19196
rect 4798 19184 4804 19187
rect 4856 19184 4862 19236
rect 6273 19227 6331 19233
rect 6273 19193 6285 19227
rect 6319 19224 6331 19227
rect 8481 19227 8539 19233
rect 6319 19196 7328 19224
rect 6319 19193 6331 19196
rect 6273 19187 6331 19193
rect 7300 19168 7328 19196
rect 8481 19193 8493 19227
rect 8527 19224 8539 19227
rect 8527 19196 9076 19224
rect 8527 19193 8539 19196
rect 8481 19187 8539 19193
rect 1397 19159 1455 19165
rect 1397 19125 1409 19159
rect 1443 19125 1455 19159
rect 1397 19119 1455 19125
rect 1670 19116 1676 19168
rect 1728 19156 1734 19168
rect 1857 19159 1915 19165
rect 1857 19156 1869 19159
rect 1728 19128 1869 19156
rect 1728 19116 1734 19128
rect 1857 19125 1869 19128
rect 1903 19125 1915 19159
rect 2958 19156 2964 19168
rect 2919 19128 2964 19156
rect 1857 19119 1915 19125
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 5534 19116 5540 19168
rect 5592 19156 5598 19168
rect 5905 19159 5963 19165
rect 5905 19156 5917 19159
rect 5592 19128 5917 19156
rect 5592 19116 5598 19128
rect 5905 19125 5917 19128
rect 5951 19125 5963 19159
rect 5905 19119 5963 19125
rect 5994 19116 6000 19168
rect 6052 19156 6058 19168
rect 6641 19159 6699 19165
rect 6641 19156 6653 19159
rect 6052 19128 6653 19156
rect 6052 19116 6058 19128
rect 6641 19125 6653 19128
rect 6687 19156 6699 19159
rect 7190 19156 7196 19168
rect 6687 19128 7196 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 7190 19116 7196 19128
rect 7248 19116 7254 19168
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 8570 19156 8576 19168
rect 7340 19128 7385 19156
rect 8531 19128 8576 19156
rect 7340 19116 7346 19128
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 8662 19116 8668 19168
rect 8720 19156 8726 19168
rect 9048 19165 9076 19196
rect 9858 19184 9864 19236
rect 9916 19224 9922 19236
rect 13814 19233 13820 19236
rect 10505 19227 10563 19233
rect 10505 19224 10517 19227
rect 9916 19196 10517 19224
rect 9916 19184 9922 19196
rect 10505 19193 10517 19196
rect 10551 19193 10563 19227
rect 13808 19224 13820 19233
rect 13775 19196 13820 19224
rect 10505 19187 10563 19193
rect 13808 19187 13820 19196
rect 13814 19184 13820 19187
rect 13872 19184 13878 19236
rect 8941 19159 8999 19165
rect 8941 19156 8953 19159
rect 8720 19128 8953 19156
rect 8720 19116 8726 19128
rect 8941 19125 8953 19128
rect 8987 19125 8999 19159
rect 8941 19119 8999 19125
rect 9033 19159 9091 19165
rect 9033 19125 9045 19159
rect 9079 19156 9091 19159
rect 9214 19156 9220 19168
rect 9079 19128 9220 19156
rect 9079 19125 9091 19128
rect 9033 19119 9091 19125
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 10134 19156 10140 19168
rect 10095 19128 10140 19156
rect 10134 19116 10140 19128
rect 10192 19116 10198 19168
rect 10962 19116 10968 19168
rect 11020 19156 11026 19168
rect 11238 19156 11244 19168
rect 11020 19128 11244 19156
rect 11020 19116 11026 19128
rect 11238 19116 11244 19128
rect 11296 19116 11302 19168
rect 12621 19159 12679 19165
rect 12621 19125 12633 19159
rect 12667 19156 12679 19159
rect 12894 19156 12900 19168
rect 12667 19128 12900 19156
rect 12667 19125 12679 19128
rect 12621 19119 12679 19125
rect 12894 19116 12900 19128
rect 12952 19116 12958 19168
rect 13078 19156 13084 19168
rect 13039 19128 13084 19156
rect 13078 19116 13084 19128
rect 13136 19116 13142 19168
rect 14921 19159 14979 19165
rect 14921 19125 14933 19159
rect 14967 19156 14979 19159
rect 15396 19156 15424 19255
rect 15838 19252 15844 19264
rect 15896 19252 15902 19304
rect 16025 19295 16083 19301
rect 16025 19261 16037 19295
rect 16071 19292 16083 19295
rect 16298 19292 16304 19304
rect 16071 19264 16304 19292
rect 16071 19261 16083 19264
rect 16025 19255 16083 19261
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 16758 19292 16764 19304
rect 16719 19264 16764 19292
rect 16758 19252 16764 19264
rect 16816 19252 16822 19304
rect 18049 19295 18107 19301
rect 18049 19261 18061 19295
rect 18095 19292 18107 19295
rect 18322 19292 18328 19304
rect 18095 19264 18328 19292
rect 18095 19261 18107 19264
rect 18049 19255 18107 19261
rect 18322 19252 18328 19264
rect 18380 19252 18386 19304
rect 18966 19252 18972 19304
rect 19024 19292 19030 19304
rect 19153 19295 19211 19301
rect 19153 19292 19165 19295
rect 19024 19264 19165 19292
rect 19024 19252 19030 19264
rect 19153 19261 19165 19264
rect 19199 19292 19211 19295
rect 19886 19292 19892 19304
rect 19199 19264 19892 19292
rect 19199 19261 19211 19264
rect 19153 19255 19211 19261
rect 19886 19252 19892 19264
rect 19944 19252 19950 19304
rect 20530 19252 20536 19304
rect 20588 19252 20594 19304
rect 21726 19292 21732 19304
rect 21687 19264 21732 19292
rect 21726 19252 21732 19264
rect 21784 19252 21790 19304
rect 23661 19295 23719 19301
rect 23661 19261 23673 19295
rect 23707 19292 23719 19295
rect 24762 19292 24768 19304
rect 23707 19264 24768 19292
rect 23707 19261 23719 19264
rect 23661 19255 23719 19261
rect 24762 19252 24768 19264
rect 24820 19252 24826 19304
rect 15749 19227 15807 19233
rect 15749 19193 15761 19227
rect 15795 19224 15807 19227
rect 15795 19196 16896 19224
rect 15795 19193 15807 19196
rect 15749 19187 15807 19193
rect 16868 19168 16896 19196
rect 18138 19184 18144 19236
rect 18196 19224 18202 19236
rect 18601 19227 18659 19233
rect 18601 19224 18613 19227
rect 18196 19196 18613 19224
rect 18196 19184 18202 19196
rect 18601 19193 18613 19196
rect 18647 19224 18659 19227
rect 19058 19224 19064 19236
rect 18647 19196 19064 19224
rect 18647 19193 18659 19196
rect 18601 19187 18659 19193
rect 19058 19184 19064 19196
rect 19116 19184 19122 19236
rect 19420 19227 19478 19233
rect 19420 19193 19432 19227
rect 19466 19224 19478 19227
rect 20070 19224 20076 19236
rect 19466 19196 20076 19224
rect 19466 19193 19478 19196
rect 19420 19187 19478 19193
rect 20070 19184 20076 19196
rect 20128 19184 20134 19236
rect 21821 19227 21879 19233
rect 21821 19224 21833 19227
rect 21192 19196 21833 19224
rect 14967 19128 15424 19156
rect 14967 19125 14979 19128
rect 14921 19119 14979 19125
rect 15470 19116 15476 19168
rect 15528 19156 15534 19168
rect 15654 19156 15660 19168
rect 15528 19128 15660 19156
rect 15528 19116 15534 19128
rect 15654 19116 15660 19128
rect 15712 19156 15718 19168
rect 15841 19159 15899 19165
rect 15841 19156 15853 19159
rect 15712 19128 15853 19156
rect 15712 19116 15718 19128
rect 15841 19125 15853 19128
rect 15887 19125 15899 19159
rect 16390 19156 16396 19168
rect 16351 19128 16396 19156
rect 15841 19119 15899 19125
rect 16390 19116 16396 19128
rect 16448 19116 16454 19168
rect 16850 19156 16856 19168
rect 16811 19128 16856 19156
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 17954 19116 17960 19168
rect 18012 19156 18018 19168
rect 18233 19159 18291 19165
rect 18233 19156 18245 19159
rect 18012 19128 18245 19156
rect 18012 19116 18018 19128
rect 18233 19125 18245 19128
rect 18279 19125 18291 19159
rect 18233 19119 18291 19125
rect 20714 19116 20720 19168
rect 20772 19156 20778 19168
rect 21192 19165 21220 19196
rect 21821 19193 21833 19196
rect 21867 19193 21879 19227
rect 23906 19227 23964 19233
rect 23906 19224 23918 19227
rect 21821 19187 21879 19193
rect 23492 19196 23918 19224
rect 23492 19168 23520 19196
rect 23906 19193 23918 19196
rect 23952 19193 23964 19227
rect 23906 19187 23964 19193
rect 25314 19184 25320 19236
rect 25372 19224 25378 19236
rect 25409 19227 25467 19233
rect 25409 19224 25421 19227
rect 25372 19196 25421 19224
rect 25372 19184 25378 19196
rect 25409 19193 25421 19196
rect 25455 19224 25467 19227
rect 25774 19224 25780 19236
rect 25455 19196 25780 19224
rect 25455 19193 25467 19196
rect 25409 19187 25467 19193
rect 25774 19184 25780 19196
rect 25832 19184 25838 19236
rect 21177 19159 21235 19165
rect 21177 19156 21189 19159
rect 20772 19128 21189 19156
rect 20772 19116 20778 19128
rect 21177 19125 21189 19128
rect 21223 19125 21235 19159
rect 21358 19156 21364 19168
rect 21319 19128 21364 19156
rect 21177 19119 21235 19125
rect 21358 19116 21364 19128
rect 21416 19116 21422 19168
rect 22370 19156 22376 19168
rect 22331 19128 22376 19156
rect 22370 19116 22376 19128
rect 22428 19116 22434 19168
rect 23474 19156 23480 19168
rect 23435 19128 23480 19156
rect 23474 19116 23480 19128
rect 23532 19116 23538 19168
rect 25038 19156 25044 19168
rect 24999 19128 25044 19156
rect 25038 19116 25044 19128
rect 25096 19156 25102 19168
rect 25222 19156 25228 19168
rect 25096 19128 25228 19156
rect 25096 19116 25102 19128
rect 25222 19116 25228 19128
rect 25280 19116 25286 19168
rect 25682 19156 25688 19168
rect 25643 19128 25688 19156
rect 25682 19116 25688 19128
rect 25740 19116 25746 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1394 18912 1400 18964
rect 1452 18952 1458 18964
rect 2317 18955 2375 18961
rect 2317 18952 2329 18955
rect 1452 18924 2329 18952
rect 1452 18912 1458 18924
rect 2317 18921 2329 18924
rect 2363 18921 2375 18955
rect 2317 18915 2375 18921
rect 3053 18955 3111 18961
rect 3053 18921 3065 18955
rect 3099 18952 3111 18955
rect 3510 18952 3516 18964
rect 3099 18924 3516 18952
rect 3099 18921 3111 18924
rect 3053 18915 3111 18921
rect 3510 18912 3516 18924
rect 3568 18912 3574 18964
rect 3786 18912 3792 18964
rect 3844 18952 3850 18964
rect 4893 18955 4951 18961
rect 4893 18952 4905 18955
rect 3844 18924 4905 18952
rect 3844 18912 3850 18924
rect 4893 18921 4905 18924
rect 4939 18921 4951 18955
rect 4893 18915 4951 18921
rect 5997 18955 6055 18961
rect 5997 18921 6009 18955
rect 6043 18952 6055 18955
rect 6822 18952 6828 18964
rect 6043 18924 6828 18952
rect 6043 18921 6055 18924
rect 5997 18915 6055 18921
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 7466 18952 7472 18964
rect 7427 18924 7472 18952
rect 7466 18912 7472 18924
rect 7524 18912 7530 18964
rect 7834 18952 7840 18964
rect 7795 18924 7840 18952
rect 7834 18912 7840 18924
rect 7892 18912 7898 18964
rect 9493 18955 9551 18961
rect 9493 18921 9505 18955
rect 9539 18952 9551 18955
rect 9674 18952 9680 18964
rect 9539 18924 9680 18952
rect 9539 18921 9551 18924
rect 9493 18915 9551 18921
rect 9674 18912 9680 18924
rect 9732 18912 9738 18964
rect 11974 18952 11980 18964
rect 11935 18924 11980 18952
rect 11974 18912 11980 18924
rect 12032 18912 12038 18964
rect 12345 18955 12403 18961
rect 12345 18921 12357 18955
rect 12391 18952 12403 18955
rect 12526 18952 12532 18964
rect 12391 18924 12532 18952
rect 12391 18921 12403 18924
rect 12345 18915 12403 18921
rect 12526 18912 12532 18924
rect 12584 18912 12590 18964
rect 13814 18952 13820 18964
rect 13727 18924 13820 18952
rect 13814 18912 13820 18924
rect 13872 18952 13878 18964
rect 14642 18952 14648 18964
rect 13872 18924 14648 18952
rect 13872 18912 13878 18924
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 16850 18912 16856 18964
rect 16908 18952 16914 18964
rect 18877 18955 18935 18961
rect 18877 18952 18889 18955
rect 16908 18924 18889 18952
rect 16908 18912 16914 18924
rect 18877 18921 18889 18924
rect 18923 18921 18935 18955
rect 18877 18915 18935 18921
rect 19058 18912 19064 18964
rect 19116 18952 19122 18964
rect 19245 18955 19303 18961
rect 19245 18952 19257 18955
rect 19116 18924 19257 18952
rect 19116 18912 19122 18924
rect 19245 18921 19257 18924
rect 19291 18952 19303 18955
rect 19518 18952 19524 18964
rect 19291 18924 19524 18952
rect 19291 18921 19303 18924
rect 19245 18915 19303 18921
rect 19518 18912 19524 18924
rect 19576 18912 19582 18964
rect 19981 18955 20039 18961
rect 19981 18921 19993 18955
rect 20027 18952 20039 18955
rect 20070 18952 20076 18964
rect 20027 18924 20076 18952
rect 20027 18921 20039 18924
rect 19981 18915 20039 18921
rect 20070 18912 20076 18924
rect 20128 18912 20134 18964
rect 20717 18955 20775 18961
rect 20717 18921 20729 18955
rect 20763 18952 20775 18955
rect 20898 18952 20904 18964
rect 20763 18924 20904 18952
rect 20763 18921 20775 18924
rect 20717 18915 20775 18921
rect 20898 18912 20904 18924
rect 20956 18912 20962 18964
rect 21082 18912 21088 18964
rect 21140 18952 21146 18964
rect 21269 18955 21327 18961
rect 21269 18952 21281 18955
rect 21140 18924 21281 18952
rect 21140 18912 21146 18924
rect 21269 18921 21281 18924
rect 21315 18952 21327 18955
rect 21315 18924 21588 18952
rect 21315 18921 21327 18924
rect 21269 18915 21327 18921
rect 21560 18896 21588 18924
rect 21726 18912 21732 18964
rect 21784 18952 21790 18964
rect 21913 18955 21971 18961
rect 21913 18952 21925 18955
rect 21784 18924 21925 18952
rect 21784 18912 21790 18924
rect 21913 18921 21925 18924
rect 21959 18921 21971 18955
rect 21913 18915 21971 18921
rect 23290 18912 23296 18964
rect 23348 18952 23354 18964
rect 23385 18955 23443 18961
rect 23385 18952 23397 18955
rect 23348 18924 23397 18952
rect 23348 18912 23354 18924
rect 23385 18921 23397 18924
rect 23431 18921 23443 18955
rect 23385 18915 23443 18921
rect 24857 18955 24915 18961
rect 24857 18921 24869 18955
rect 24903 18952 24915 18955
rect 25317 18955 25375 18961
rect 25317 18952 25329 18955
rect 24903 18924 25329 18952
rect 24903 18921 24915 18924
rect 24857 18915 24915 18921
rect 25317 18921 25329 18924
rect 25363 18921 25375 18955
rect 25317 18915 25375 18921
rect 4617 18887 4675 18893
rect 4617 18853 4629 18887
rect 4663 18884 4675 18887
rect 4798 18884 4804 18896
rect 4663 18856 4804 18884
rect 4663 18853 4675 18856
rect 4617 18847 4675 18853
rect 4798 18844 4804 18856
rect 4856 18884 4862 18896
rect 6270 18884 6276 18896
rect 4856 18856 5580 18884
rect 6231 18856 6276 18884
rect 4856 18844 4862 18856
rect 5258 18816 5264 18828
rect 5219 18788 5264 18816
rect 5258 18776 5264 18788
rect 5316 18776 5322 18828
rect 5552 18816 5580 18856
rect 6270 18844 6276 18856
rect 6328 18844 6334 18896
rect 9398 18844 9404 18896
rect 9456 18884 9462 18896
rect 9944 18887 10002 18893
rect 9944 18884 9956 18887
rect 9456 18856 9956 18884
rect 9456 18844 9462 18856
rect 9944 18853 9956 18856
rect 9990 18884 10002 18887
rect 10686 18884 10692 18896
rect 9990 18856 10692 18884
rect 9990 18853 10002 18856
rect 9944 18847 10002 18853
rect 10686 18844 10692 18856
rect 10744 18844 10750 18896
rect 12802 18884 12808 18896
rect 12452 18856 12808 18884
rect 6288 18816 6316 18844
rect 5552 18788 6316 18816
rect 2038 18708 2044 18760
rect 2096 18748 2102 18760
rect 2406 18748 2412 18760
rect 2096 18720 2412 18748
rect 2096 18708 2102 18720
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 2501 18751 2559 18757
rect 2501 18717 2513 18751
rect 2547 18717 2559 18751
rect 2501 18711 2559 18717
rect 3881 18751 3939 18757
rect 3881 18717 3893 18751
rect 3927 18748 3939 18751
rect 5166 18748 5172 18760
rect 3927 18720 5172 18748
rect 3927 18717 3939 18720
rect 3881 18711 3939 18717
rect 2516 18680 2544 18711
rect 5166 18708 5172 18720
rect 5224 18748 5230 18760
rect 5552 18757 5580 18788
rect 6362 18776 6368 18828
rect 6420 18816 6426 18828
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 6420 18788 6837 18816
rect 6420 18776 6426 18788
rect 6825 18785 6837 18788
rect 6871 18785 6883 18819
rect 8386 18816 8392 18828
rect 8347 18788 8392 18816
rect 6825 18779 6883 18785
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 12452 18825 12480 18856
rect 12802 18844 12808 18856
rect 12860 18884 12866 18896
rect 12986 18884 12992 18896
rect 12860 18856 12992 18884
rect 12860 18844 12866 18856
rect 12986 18844 12992 18856
rect 13044 18844 13050 18896
rect 15657 18887 15715 18893
rect 15657 18853 15669 18887
rect 15703 18884 15715 18887
rect 16022 18884 16028 18896
rect 15703 18856 16028 18884
rect 15703 18853 15715 18856
rect 15657 18847 15715 18853
rect 16022 18844 16028 18856
rect 16080 18844 16086 18896
rect 18230 18844 18236 18896
rect 18288 18884 18294 18896
rect 18325 18887 18383 18893
rect 18325 18884 18337 18887
rect 18288 18856 18337 18884
rect 18288 18844 18294 18856
rect 18325 18853 18337 18856
rect 18371 18853 18383 18887
rect 18690 18884 18696 18896
rect 18651 18856 18696 18884
rect 18325 18847 18383 18853
rect 18690 18844 18696 18856
rect 18748 18844 18754 18896
rect 19334 18884 19340 18896
rect 19295 18856 19340 18884
rect 19334 18844 19340 18856
rect 19392 18844 19398 18896
rect 19996 18856 21496 18884
rect 19996 18828 20024 18856
rect 9677 18819 9735 18825
rect 9677 18785 9689 18819
rect 9723 18816 9735 18819
rect 12437 18819 12495 18825
rect 9723 18788 10732 18816
rect 9723 18785 9735 18788
rect 9677 18779 9735 18785
rect 10704 18760 10732 18788
rect 12437 18785 12449 18819
rect 12483 18785 12495 18819
rect 12437 18779 12495 18785
rect 12526 18776 12532 18828
rect 12584 18816 12590 18828
rect 12704 18819 12762 18825
rect 12704 18816 12716 18819
rect 12584 18788 12716 18816
rect 12584 18776 12590 18788
rect 12704 18785 12716 18788
rect 12750 18816 12762 18819
rect 13722 18816 13728 18828
rect 12750 18788 13728 18816
rect 12750 18785 12762 18788
rect 12704 18779 12762 18785
rect 13722 18776 13728 18788
rect 13780 18776 13786 18828
rect 14458 18816 14464 18828
rect 14419 18788 14464 18816
rect 14458 18776 14464 18788
rect 14516 18776 14522 18828
rect 15105 18819 15163 18825
rect 15105 18785 15117 18819
rect 15151 18816 15163 18819
rect 15378 18816 15384 18828
rect 15151 18788 15384 18816
rect 15151 18785 15163 18788
rect 15105 18779 15163 18785
rect 15378 18776 15384 18788
rect 15436 18776 15442 18828
rect 16942 18825 16948 18828
rect 16485 18819 16543 18825
rect 16485 18785 16497 18819
rect 16531 18816 16543 18819
rect 16936 18816 16948 18825
rect 16531 18788 16948 18816
rect 16531 18785 16543 18788
rect 16485 18779 16543 18785
rect 16936 18779 16948 18788
rect 16942 18776 16948 18779
rect 17000 18776 17006 18828
rect 17954 18776 17960 18828
rect 18012 18816 18018 18828
rect 19150 18816 19156 18828
rect 18012 18788 19156 18816
rect 18012 18776 18018 18788
rect 19150 18776 19156 18788
rect 19208 18816 19214 18828
rect 19208 18788 19472 18816
rect 19208 18776 19214 18788
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 5224 18720 5365 18748
rect 5224 18708 5230 18720
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 5537 18751 5595 18757
rect 5537 18717 5549 18751
rect 5583 18717 5595 18751
rect 5537 18711 5595 18717
rect 6086 18708 6092 18760
rect 6144 18748 6150 18760
rect 6917 18751 6975 18757
rect 6917 18748 6929 18751
rect 6144 18720 6929 18748
rect 6144 18708 6150 18720
rect 6917 18717 6929 18720
rect 6963 18717 6975 18751
rect 6917 18711 6975 18717
rect 7009 18751 7067 18757
rect 7009 18717 7021 18751
rect 7055 18717 7067 18751
rect 8478 18748 8484 18760
rect 8439 18720 8484 18748
rect 7009 18711 7067 18717
rect 1872 18652 2544 18680
rect 1872 18624 1900 18652
rect 6546 18640 6552 18692
rect 6604 18680 6610 18692
rect 7024 18680 7052 18711
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 8573 18751 8631 18757
rect 8573 18717 8585 18751
rect 8619 18717 8631 18751
rect 8573 18711 8631 18717
rect 6604 18652 7052 18680
rect 6604 18640 6610 18652
rect 7650 18640 7656 18692
rect 7708 18680 7714 18692
rect 8588 18680 8616 18711
rect 10686 18708 10692 18760
rect 10744 18708 10750 18760
rect 15654 18708 15660 18760
rect 15712 18748 15718 18760
rect 16390 18748 16396 18760
rect 15712 18720 16396 18748
rect 15712 18708 15718 18720
rect 16390 18708 16396 18720
rect 16448 18748 16454 18760
rect 19444 18757 19472 18788
rect 19978 18776 19984 18828
rect 20036 18776 20042 18828
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 16448 18720 16681 18748
rect 16448 18708 16454 18720
rect 16669 18717 16681 18720
rect 16715 18717 16727 18751
rect 16669 18711 16727 18717
rect 19429 18751 19487 18757
rect 19429 18717 19441 18751
rect 19475 18717 19487 18751
rect 21358 18748 21364 18760
rect 21319 18720 21364 18748
rect 19429 18711 19487 18717
rect 21358 18708 21364 18720
rect 21416 18708 21422 18760
rect 21468 18757 21496 18856
rect 21542 18844 21548 18896
rect 21600 18884 21606 18896
rect 22278 18884 22284 18896
rect 21600 18856 22284 18884
rect 21600 18844 21606 18856
rect 22278 18844 22284 18856
rect 22336 18844 22342 18896
rect 24946 18884 24952 18896
rect 24907 18856 24952 18884
rect 24946 18844 24952 18856
rect 25004 18844 25010 18896
rect 25590 18884 25596 18896
rect 25551 18856 25596 18884
rect 25590 18844 25596 18856
rect 25648 18844 25654 18896
rect 23014 18776 23020 18828
rect 23072 18816 23078 18828
rect 23293 18819 23351 18825
rect 23293 18816 23305 18819
rect 23072 18788 23305 18816
rect 23072 18776 23078 18788
rect 23293 18785 23305 18788
rect 23339 18785 23351 18819
rect 24305 18819 24363 18825
rect 24305 18816 24317 18819
rect 23293 18779 23351 18785
rect 23400 18788 24317 18816
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18717 21511 18751
rect 21453 18711 21511 18717
rect 21726 18708 21732 18760
rect 21784 18748 21790 18760
rect 23400 18748 23428 18788
rect 24305 18785 24317 18788
rect 24351 18785 24363 18819
rect 24305 18779 24363 18785
rect 24762 18776 24768 18828
rect 24820 18816 24826 18828
rect 25869 18819 25927 18825
rect 25869 18816 25881 18819
rect 24820 18788 25881 18816
rect 24820 18776 24826 18788
rect 25869 18785 25881 18788
rect 25915 18785 25927 18819
rect 25869 18779 25927 18785
rect 21784 18720 23428 18748
rect 21784 18708 21790 18720
rect 23474 18708 23480 18760
rect 23532 18748 23538 18760
rect 23532 18720 23577 18748
rect 23532 18708 23538 18720
rect 25038 18708 25044 18760
rect 25096 18748 25102 18760
rect 25096 18720 25141 18748
rect 25096 18708 25102 18720
rect 9033 18683 9091 18689
rect 9033 18680 9045 18683
rect 7708 18652 9045 18680
rect 7708 18640 7714 18652
rect 9033 18649 9045 18652
rect 9079 18680 9091 18683
rect 9122 18680 9128 18692
rect 9079 18652 9128 18680
rect 9079 18649 9091 18652
rect 9033 18643 9091 18649
rect 9122 18640 9128 18652
rect 9180 18680 9186 18692
rect 9582 18680 9588 18692
rect 9180 18652 9588 18680
rect 9180 18640 9186 18652
rect 9582 18640 9588 18652
rect 9640 18640 9646 18692
rect 20901 18683 20959 18689
rect 20901 18649 20913 18683
rect 20947 18680 20959 18683
rect 22186 18680 22192 18692
rect 20947 18652 22192 18680
rect 20947 18649 20959 18652
rect 20901 18643 20959 18649
rect 22186 18640 22192 18652
rect 22244 18680 22250 18692
rect 22281 18683 22339 18689
rect 22281 18680 22293 18683
rect 22244 18652 22293 18680
rect 22244 18640 22250 18652
rect 22281 18649 22293 18652
rect 22327 18649 22339 18683
rect 22281 18643 22339 18649
rect 22833 18683 22891 18689
rect 22833 18649 22845 18683
rect 22879 18680 22891 18683
rect 23492 18680 23520 18708
rect 22879 18652 23520 18680
rect 22879 18649 22891 18652
rect 22833 18643 22891 18649
rect 23566 18640 23572 18692
rect 23624 18680 23630 18692
rect 24489 18683 24547 18689
rect 24489 18680 24501 18683
rect 23624 18652 24501 18680
rect 23624 18640 23630 18652
rect 24489 18649 24501 18652
rect 24535 18649 24547 18683
rect 24489 18643 24547 18649
rect 25317 18683 25375 18689
rect 25317 18649 25329 18683
rect 25363 18680 25375 18683
rect 25866 18680 25872 18692
rect 25363 18652 25872 18680
rect 25363 18649 25375 18652
rect 25317 18643 25375 18649
rect 25866 18640 25872 18652
rect 25924 18640 25930 18692
rect 1854 18612 1860 18624
rect 1815 18584 1860 18612
rect 1854 18572 1860 18584
rect 1912 18572 1918 18624
rect 1946 18572 1952 18624
rect 2004 18612 2010 18624
rect 2004 18584 2049 18612
rect 2004 18572 2010 18584
rect 2222 18572 2228 18624
rect 2280 18612 2286 18624
rect 3418 18612 3424 18624
rect 2280 18584 3424 18612
rect 2280 18572 2286 18584
rect 3418 18572 3424 18584
rect 3476 18572 3482 18624
rect 6454 18612 6460 18624
rect 6415 18584 6460 18612
rect 6454 18572 6460 18584
rect 6512 18572 6518 18624
rect 8018 18612 8024 18624
rect 7979 18584 8024 18612
rect 8018 18572 8024 18584
rect 8076 18572 8082 18624
rect 11054 18612 11060 18624
rect 11015 18584 11060 18612
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 11422 18612 11428 18624
rect 11335 18584 11428 18612
rect 11422 18572 11428 18584
rect 11480 18612 11486 18624
rect 12342 18612 12348 18624
rect 11480 18584 12348 18612
rect 11480 18572 11486 18584
rect 12342 18572 12348 18584
rect 12400 18572 12406 18624
rect 13998 18572 14004 18624
rect 14056 18612 14062 18624
rect 14093 18615 14151 18621
rect 14093 18612 14105 18615
rect 14056 18584 14105 18612
rect 14056 18572 14062 18584
rect 14093 18581 14105 18584
rect 14139 18581 14151 18615
rect 14093 18575 14151 18581
rect 18049 18615 18107 18621
rect 18049 18581 18061 18615
rect 18095 18612 18107 18615
rect 18138 18612 18144 18624
rect 18095 18584 18144 18612
rect 18095 18581 18107 18584
rect 18049 18575 18107 18581
rect 18138 18572 18144 18584
rect 18196 18572 18202 18624
rect 20346 18612 20352 18624
rect 20307 18584 20352 18612
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 22922 18612 22928 18624
rect 22883 18584 22928 18612
rect 22922 18572 22928 18584
rect 22980 18572 22986 18624
rect 23842 18572 23848 18624
rect 23900 18612 23906 18624
rect 23937 18615 23995 18621
rect 23937 18612 23949 18615
rect 23900 18584 23949 18612
rect 23900 18572 23906 18584
rect 23937 18581 23949 18584
rect 23983 18581 23995 18615
rect 23937 18575 23995 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1394 18368 1400 18420
rect 1452 18408 1458 18420
rect 1581 18411 1639 18417
rect 1581 18408 1593 18411
rect 1452 18380 1593 18408
rect 1452 18368 1458 18380
rect 1581 18377 1593 18380
rect 1627 18377 1639 18411
rect 6546 18408 6552 18420
rect 6507 18380 6552 18408
rect 1581 18371 1639 18377
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 8478 18368 8484 18420
rect 8536 18408 8542 18420
rect 10505 18411 10563 18417
rect 10505 18408 10517 18411
rect 8536 18380 10517 18408
rect 8536 18368 8542 18380
rect 10505 18377 10517 18380
rect 10551 18377 10563 18411
rect 10505 18371 10563 18377
rect 11885 18411 11943 18417
rect 11885 18377 11897 18411
rect 11931 18408 11943 18411
rect 12066 18408 12072 18420
rect 11931 18380 12072 18408
rect 11931 18377 11943 18380
rect 11885 18371 11943 18377
rect 12066 18368 12072 18380
rect 12124 18408 12130 18420
rect 12526 18408 12532 18420
rect 12124 18380 12532 18408
rect 12124 18368 12130 18380
rect 12526 18368 12532 18380
rect 12584 18368 12590 18420
rect 12805 18411 12863 18417
rect 12805 18377 12817 18411
rect 12851 18408 12863 18411
rect 13262 18408 13268 18420
rect 12851 18380 13268 18408
rect 12851 18377 12863 18380
rect 12805 18371 12863 18377
rect 13262 18368 13268 18380
rect 13320 18368 13326 18420
rect 13814 18408 13820 18420
rect 13775 18380 13820 18408
rect 13814 18368 13820 18380
rect 13872 18368 13878 18420
rect 14366 18408 14372 18420
rect 14327 18380 14372 18408
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 15473 18411 15531 18417
rect 15473 18377 15485 18411
rect 15519 18408 15531 18411
rect 15562 18408 15568 18420
rect 15519 18380 15568 18408
rect 15519 18377 15531 18380
rect 15473 18371 15531 18377
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 16301 18411 16359 18417
rect 16301 18377 16313 18411
rect 16347 18408 16359 18411
rect 16942 18408 16948 18420
rect 16347 18380 16948 18408
rect 16347 18377 16359 18380
rect 16301 18371 16359 18377
rect 16942 18368 16948 18380
rect 17000 18368 17006 18420
rect 19518 18408 19524 18420
rect 19479 18380 19524 18408
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 20346 18368 20352 18420
rect 20404 18408 20410 18420
rect 21358 18408 21364 18420
rect 20404 18380 21364 18408
rect 20404 18368 20410 18380
rect 21358 18368 21364 18380
rect 21416 18408 21422 18420
rect 21821 18411 21879 18417
rect 21821 18408 21833 18411
rect 21416 18380 21833 18408
rect 21416 18368 21422 18380
rect 21821 18377 21833 18380
rect 21867 18377 21879 18411
rect 23290 18408 23296 18420
rect 23251 18380 23296 18408
rect 21821 18371 21879 18377
rect 23290 18368 23296 18380
rect 23348 18368 23354 18420
rect 23474 18368 23480 18420
rect 23532 18408 23538 18420
rect 25041 18411 25099 18417
rect 25041 18408 25053 18411
rect 23532 18380 25053 18408
rect 23532 18368 23538 18380
rect 25041 18377 25053 18380
rect 25087 18377 25099 18411
rect 25041 18371 25099 18377
rect 25777 18411 25835 18417
rect 25777 18377 25789 18411
rect 25823 18408 25835 18411
rect 25866 18408 25872 18420
rect 25823 18380 25872 18408
rect 25823 18377 25835 18380
rect 25777 18371 25835 18377
rect 25866 18368 25872 18380
rect 25924 18368 25930 18420
rect 5721 18343 5779 18349
rect 5721 18309 5733 18343
rect 5767 18340 5779 18343
rect 5902 18340 5908 18352
rect 5767 18312 5908 18340
rect 5767 18309 5779 18312
rect 5721 18303 5779 18309
rect 5902 18300 5908 18312
rect 5960 18340 5966 18352
rect 6730 18340 6736 18352
rect 5960 18312 6736 18340
rect 5960 18300 5966 18312
rect 6730 18300 6736 18312
rect 6788 18300 6794 18352
rect 9582 18300 9588 18352
rect 9640 18340 9646 18352
rect 9677 18343 9735 18349
rect 9677 18340 9689 18343
rect 9640 18312 9689 18340
rect 9640 18300 9646 18312
rect 9677 18309 9689 18312
rect 9723 18309 9735 18343
rect 9950 18340 9956 18352
rect 9911 18312 9956 18340
rect 9677 18303 9735 18309
rect 9950 18300 9956 18312
rect 10008 18340 10014 18352
rect 10229 18343 10287 18349
rect 10229 18340 10241 18343
rect 10008 18312 10241 18340
rect 10008 18300 10014 18312
rect 10229 18309 10241 18312
rect 10275 18309 10287 18343
rect 10229 18303 10287 18309
rect 16393 18343 16451 18349
rect 16393 18309 16405 18343
rect 16439 18309 16451 18343
rect 16393 18303 16451 18309
rect 4154 18272 4160 18284
rect 3252 18244 4160 18272
rect 1762 18164 1768 18216
rect 1820 18204 1826 18216
rect 2133 18207 2191 18213
rect 2133 18204 2145 18207
rect 1820 18176 2145 18204
rect 1820 18164 1826 18176
rect 2133 18173 2145 18176
rect 2179 18204 2191 18207
rect 3252 18204 3280 18244
rect 4154 18232 4160 18244
rect 4212 18272 4218 18284
rect 4341 18275 4399 18281
rect 4341 18272 4353 18275
rect 4212 18244 4353 18272
rect 4212 18232 4218 18244
rect 4341 18241 4353 18244
rect 4387 18241 4399 18275
rect 11054 18272 11060 18284
rect 4341 18235 4399 18241
rect 10060 18244 11060 18272
rect 2179 18176 3280 18204
rect 2179 18173 2191 18176
rect 2133 18167 2191 18173
rect 3510 18164 3516 18216
rect 3568 18204 3574 18216
rect 3694 18204 3700 18216
rect 3568 18176 3700 18204
rect 3568 18164 3574 18176
rect 3694 18164 3700 18176
rect 3752 18164 3758 18216
rect 6086 18204 6092 18216
rect 6047 18176 6092 18204
rect 6086 18164 6092 18176
rect 6144 18164 6150 18216
rect 6822 18204 6828 18216
rect 6783 18176 6828 18204
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 8110 18164 8116 18216
rect 8168 18204 8174 18216
rect 8297 18207 8355 18213
rect 8297 18204 8309 18207
rect 8168 18176 8309 18204
rect 8168 18164 8174 18176
rect 8297 18173 8309 18176
rect 8343 18204 8355 18207
rect 8938 18204 8944 18216
rect 8343 18176 8944 18204
rect 8343 18173 8355 18176
rect 8297 18167 8355 18173
rect 8938 18164 8944 18176
rect 8996 18164 9002 18216
rect 10060 18148 10088 18244
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 12250 18272 12256 18284
rect 12163 18244 12256 18272
rect 12250 18232 12256 18244
rect 12308 18272 12314 18284
rect 13449 18275 13507 18281
rect 13449 18272 13461 18275
rect 12308 18244 13461 18272
rect 12308 18232 12314 18244
rect 13449 18241 13461 18244
rect 13495 18272 13507 18275
rect 13998 18272 14004 18284
rect 13495 18244 14004 18272
rect 13495 18241 13507 18244
rect 13449 18235 13507 18241
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 14182 18232 14188 18284
rect 14240 18272 14246 18284
rect 14921 18275 14979 18281
rect 14921 18272 14933 18275
rect 14240 18244 14933 18272
rect 14240 18232 14246 18244
rect 14921 18241 14933 18244
rect 14967 18241 14979 18275
rect 14921 18235 14979 18241
rect 10229 18207 10287 18213
rect 10229 18173 10241 18207
rect 10275 18204 10287 18207
rect 10965 18207 11023 18213
rect 10965 18204 10977 18207
rect 10275 18176 10977 18204
rect 10275 18173 10287 18176
rect 10229 18167 10287 18173
rect 10965 18173 10977 18176
rect 11011 18173 11023 18207
rect 10965 18167 11023 18173
rect 14458 18164 14464 18216
rect 14516 18204 14522 18216
rect 14737 18207 14795 18213
rect 14737 18204 14749 18207
rect 14516 18176 14749 18204
rect 14516 18164 14522 18176
rect 14737 18173 14749 18176
rect 14783 18173 14795 18207
rect 16408 18204 16436 18303
rect 21082 18300 21088 18352
rect 21140 18340 21146 18352
rect 21269 18343 21327 18349
rect 21269 18340 21281 18343
rect 21140 18312 21281 18340
rect 21140 18300 21146 18312
rect 21269 18309 21281 18312
rect 21315 18309 21327 18343
rect 21269 18303 21327 18309
rect 21542 18300 21548 18352
rect 21600 18340 21606 18352
rect 21637 18343 21695 18349
rect 21637 18340 21649 18343
rect 21600 18312 21649 18340
rect 21600 18300 21606 18312
rect 21637 18309 21649 18312
rect 21683 18309 21695 18343
rect 21637 18303 21695 18309
rect 16942 18232 16948 18284
rect 17000 18272 17006 18284
rect 17037 18275 17095 18281
rect 17037 18272 17049 18275
rect 17000 18244 17049 18272
rect 17000 18232 17006 18244
rect 17037 18241 17049 18244
rect 17083 18272 17095 18275
rect 17494 18272 17500 18284
rect 17083 18244 17500 18272
rect 17083 18241 17095 18244
rect 17037 18235 17095 18241
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 17865 18275 17923 18281
rect 17865 18241 17877 18275
rect 17911 18272 17923 18275
rect 18138 18272 18144 18284
rect 17911 18244 18144 18272
rect 17911 18241 17923 18244
rect 17865 18235 17923 18241
rect 18138 18232 18144 18244
rect 18196 18272 18202 18284
rect 18601 18275 18659 18281
rect 18601 18272 18613 18275
rect 18196 18244 18613 18272
rect 18196 18232 18202 18244
rect 18601 18241 18613 18244
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 18966 18232 18972 18284
rect 19024 18272 19030 18284
rect 19518 18272 19524 18284
rect 19024 18244 19524 18272
rect 19024 18232 19030 18244
rect 19518 18232 19524 18244
rect 19576 18272 19582 18284
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 19576 18244 19625 18272
rect 19576 18232 19582 18244
rect 19613 18241 19625 18244
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 21910 18232 21916 18284
rect 21968 18272 21974 18284
rect 22373 18275 22431 18281
rect 22373 18272 22385 18275
rect 21968 18244 22385 18272
rect 21968 18232 21974 18244
rect 22373 18241 22385 18244
rect 22419 18241 22431 18275
rect 22373 18235 22431 18241
rect 25038 18232 25044 18284
rect 25096 18272 25102 18284
rect 25317 18275 25375 18281
rect 25317 18272 25329 18275
rect 25096 18244 25329 18272
rect 25096 18232 25102 18244
rect 25317 18241 25329 18244
rect 25363 18241 25375 18275
rect 25317 18235 25375 18241
rect 17770 18204 17776 18216
rect 16408 18176 17776 18204
rect 14737 18167 14795 18173
rect 17770 18164 17776 18176
rect 17828 18204 17834 18216
rect 18417 18207 18475 18213
rect 18417 18204 18429 18207
rect 17828 18176 18429 18204
rect 17828 18164 17834 18176
rect 18417 18173 18429 18176
rect 18463 18173 18475 18207
rect 18417 18167 18475 18173
rect 18509 18207 18567 18213
rect 18509 18173 18521 18207
rect 18555 18204 18567 18207
rect 18690 18204 18696 18216
rect 18555 18176 18696 18204
rect 18555 18173 18567 18176
rect 18509 18167 18567 18173
rect 18690 18164 18696 18176
rect 18748 18164 18754 18216
rect 19153 18207 19211 18213
rect 19153 18173 19165 18207
rect 19199 18204 19211 18207
rect 19242 18204 19248 18216
rect 19199 18176 19248 18204
rect 19199 18173 19211 18176
rect 19153 18167 19211 18173
rect 19242 18164 19248 18176
rect 19300 18164 19306 18216
rect 22278 18204 22284 18216
rect 22239 18176 22284 18204
rect 22278 18164 22284 18176
rect 22336 18164 22342 18216
rect 23661 18207 23719 18213
rect 23661 18173 23673 18207
rect 23707 18204 23719 18207
rect 24854 18204 24860 18216
rect 23707 18176 24860 18204
rect 23707 18173 23719 18176
rect 23661 18167 23719 18173
rect 24854 18164 24860 18176
rect 24912 18164 24918 18216
rect 2406 18145 2412 18148
rect 2400 18136 2412 18145
rect 2319 18108 2412 18136
rect 2400 18099 2412 18108
rect 2464 18136 2470 18148
rect 3142 18136 3148 18148
rect 2464 18108 3148 18136
rect 2406 18096 2412 18099
rect 2464 18096 2470 18108
rect 3142 18096 3148 18108
rect 3200 18096 3206 18148
rect 4157 18139 4215 18145
rect 4157 18136 4169 18139
rect 3528 18108 4169 18136
rect 2038 18068 2044 18080
rect 1999 18040 2044 18068
rect 2038 18028 2044 18040
rect 2096 18028 2102 18080
rect 2774 18028 2780 18080
rect 2832 18068 2838 18080
rect 3528 18077 3556 18108
rect 4157 18105 4169 18108
rect 4203 18136 4215 18139
rect 4586 18139 4644 18145
rect 4586 18136 4598 18139
rect 4203 18108 4598 18136
rect 4203 18105 4215 18108
rect 4157 18099 4215 18105
rect 4586 18105 4598 18108
rect 4632 18105 4644 18139
rect 7098 18136 7104 18148
rect 7059 18108 7104 18136
rect 4586 18099 4644 18105
rect 7098 18096 7104 18108
rect 7156 18096 7162 18148
rect 8205 18139 8263 18145
rect 8205 18105 8217 18139
rect 8251 18136 8263 18139
rect 8542 18139 8600 18145
rect 8542 18136 8554 18139
rect 8251 18108 8554 18136
rect 8251 18105 8263 18108
rect 8205 18099 8263 18105
rect 8542 18105 8554 18108
rect 8588 18136 8600 18139
rect 10042 18136 10048 18148
rect 8588 18108 10048 18136
rect 8588 18105 8600 18108
rect 8542 18099 8600 18105
rect 10042 18096 10048 18108
rect 10100 18096 10106 18148
rect 10413 18139 10471 18145
rect 10413 18105 10425 18139
rect 10459 18136 10471 18139
rect 10870 18136 10876 18148
rect 10459 18108 10876 18136
rect 10459 18105 10471 18108
rect 10413 18099 10471 18105
rect 3513 18071 3571 18077
rect 3513 18068 3525 18071
rect 2832 18040 3525 18068
rect 2832 18028 2838 18040
rect 3513 18037 3525 18040
rect 3559 18037 3571 18071
rect 3786 18068 3792 18080
rect 3747 18040 3792 18068
rect 3513 18031 3571 18037
rect 3786 18028 3792 18040
rect 3844 18028 3850 18080
rect 7650 18028 7656 18080
rect 7708 18068 7714 18080
rect 7745 18071 7803 18077
rect 7745 18068 7757 18071
rect 7708 18040 7757 18068
rect 7708 18028 7714 18040
rect 7745 18037 7757 18040
rect 7791 18037 7803 18071
rect 7745 18031 7803 18037
rect 9950 18028 9956 18080
rect 10008 18068 10014 18080
rect 10428 18068 10456 18099
rect 10870 18096 10876 18108
rect 10928 18096 10934 18148
rect 13265 18139 13323 18145
rect 13265 18136 13277 18139
rect 12636 18108 13277 18136
rect 12636 18080 12664 18108
rect 13265 18105 13277 18108
rect 13311 18136 13323 18139
rect 13446 18136 13452 18148
rect 13311 18108 13452 18136
rect 13311 18105 13323 18108
rect 13265 18099 13323 18105
rect 13446 18096 13452 18108
rect 13504 18096 13510 18148
rect 15933 18139 15991 18145
rect 15933 18105 15945 18139
rect 15979 18136 15991 18139
rect 16761 18139 16819 18145
rect 15979 18108 16712 18136
rect 15979 18105 15991 18108
rect 15933 18099 15991 18105
rect 12618 18068 12624 18080
rect 10008 18040 10456 18068
rect 12579 18040 12624 18068
rect 10008 18028 10014 18040
rect 12618 18028 12624 18040
rect 12676 18028 12682 18080
rect 12802 18028 12808 18080
rect 12860 18068 12866 18080
rect 13173 18071 13231 18077
rect 13173 18068 13185 18071
rect 12860 18040 13185 18068
rect 12860 18028 12866 18040
rect 13173 18037 13185 18040
rect 13219 18037 13231 18071
rect 14182 18068 14188 18080
rect 14143 18040 14188 18068
rect 13173 18031 13231 18037
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 14366 18028 14372 18080
rect 14424 18068 14430 18080
rect 14829 18071 14887 18077
rect 14829 18068 14841 18071
rect 14424 18040 14841 18068
rect 14424 18028 14430 18040
rect 14829 18037 14841 18040
rect 14875 18037 14887 18071
rect 16684 18068 16712 18108
rect 16761 18105 16773 18139
rect 16807 18136 16819 18139
rect 17862 18136 17868 18148
rect 16807 18108 17868 18136
rect 16807 18105 16819 18108
rect 16761 18099 16819 18105
rect 17862 18096 17868 18108
rect 17920 18096 17926 18148
rect 19880 18139 19938 18145
rect 19880 18105 19892 18139
rect 19926 18136 19938 18139
rect 19978 18136 19984 18148
rect 19926 18108 19984 18136
rect 19926 18105 19938 18108
rect 19880 18099 19938 18105
rect 19978 18096 19984 18108
rect 20036 18096 20042 18148
rect 22186 18136 22192 18148
rect 22147 18108 22192 18136
rect 22186 18096 22192 18108
rect 22244 18096 22250 18148
rect 23842 18096 23848 18148
rect 23900 18145 23906 18148
rect 23900 18139 23964 18145
rect 23900 18105 23918 18139
rect 23952 18105 23964 18139
rect 23900 18099 23964 18105
rect 23900 18096 23906 18099
rect 25590 18096 25596 18148
rect 25648 18136 25654 18148
rect 26053 18139 26111 18145
rect 26053 18136 26065 18139
rect 25648 18108 26065 18136
rect 25648 18096 25654 18108
rect 26053 18105 26065 18108
rect 26099 18105 26111 18139
rect 26053 18099 26111 18105
rect 16850 18068 16856 18080
rect 16684 18040 16856 18068
rect 14829 18031 14887 18037
rect 16850 18028 16856 18040
rect 16908 18028 16914 18080
rect 17494 18068 17500 18080
rect 17455 18040 17500 18068
rect 17494 18028 17500 18040
rect 17552 18028 17558 18080
rect 18049 18071 18107 18077
rect 18049 18037 18061 18071
rect 18095 18068 18107 18071
rect 18230 18068 18236 18080
rect 18095 18040 18236 18068
rect 18095 18037 18107 18040
rect 18049 18031 18107 18037
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 20993 18071 21051 18077
rect 20993 18068 21005 18071
rect 20772 18040 21005 18068
rect 20772 18028 20778 18040
rect 20993 18037 21005 18040
rect 21039 18037 21051 18071
rect 23014 18068 23020 18080
rect 22927 18040 23020 18068
rect 20993 18031 21051 18037
rect 23014 18028 23020 18040
rect 23072 18068 23078 18080
rect 23290 18068 23296 18080
rect 23072 18040 23296 18068
rect 23072 18028 23078 18040
rect 23290 18028 23296 18040
rect 23348 18028 23354 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 3142 17864 3148 17876
rect 3055 17836 3148 17864
rect 3142 17824 3148 17836
rect 3200 17864 3206 17876
rect 3786 17864 3792 17876
rect 3200 17836 3792 17864
rect 3200 17824 3206 17836
rect 3786 17824 3792 17836
rect 3844 17824 3850 17876
rect 4246 17864 4252 17876
rect 4207 17836 4252 17864
rect 4246 17824 4252 17836
rect 4304 17824 4310 17876
rect 4798 17824 4804 17876
rect 4856 17864 4862 17876
rect 4893 17867 4951 17873
rect 4893 17864 4905 17867
rect 4856 17836 4905 17864
rect 4856 17824 4862 17836
rect 4893 17833 4905 17836
rect 4939 17833 4951 17867
rect 5258 17864 5264 17876
rect 5171 17836 5264 17864
rect 4893 17827 4951 17833
rect 5258 17824 5264 17836
rect 5316 17864 5322 17876
rect 6917 17867 6975 17873
rect 6917 17864 6929 17867
rect 5316 17836 6929 17864
rect 5316 17824 5322 17836
rect 6917 17833 6929 17836
rect 6963 17833 6975 17867
rect 6917 17827 6975 17833
rect 8478 17824 8484 17876
rect 8536 17864 8542 17876
rect 9033 17867 9091 17873
rect 9033 17864 9045 17867
rect 8536 17836 9045 17864
rect 8536 17824 8542 17836
rect 9033 17833 9045 17836
rect 9079 17833 9091 17867
rect 9398 17864 9404 17876
rect 9359 17836 9404 17864
rect 9033 17827 9091 17833
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 10042 17824 10048 17876
rect 10100 17864 10106 17876
rect 10597 17867 10655 17873
rect 10597 17864 10609 17867
rect 10100 17836 10609 17864
rect 10100 17824 10106 17836
rect 10597 17833 10609 17836
rect 10643 17864 10655 17867
rect 10870 17864 10876 17876
rect 10643 17836 10876 17864
rect 10643 17833 10655 17836
rect 10597 17827 10655 17833
rect 10870 17824 10876 17836
rect 10928 17824 10934 17876
rect 12342 17824 12348 17876
rect 12400 17864 12406 17876
rect 13173 17867 13231 17873
rect 13173 17864 13185 17867
rect 12400 17836 13185 17864
rect 12400 17824 12406 17836
rect 13173 17833 13185 17836
rect 13219 17833 13231 17867
rect 14366 17864 14372 17876
rect 14327 17836 14372 17864
rect 13173 17827 13231 17833
rect 14366 17824 14372 17836
rect 14424 17824 14430 17876
rect 15565 17867 15623 17873
rect 15565 17833 15577 17867
rect 15611 17864 15623 17867
rect 15746 17864 15752 17876
rect 15611 17836 15752 17864
rect 15611 17833 15623 17836
rect 15565 17827 15623 17833
rect 15746 17824 15752 17836
rect 15804 17824 15810 17876
rect 17494 17824 17500 17876
rect 17552 17864 17558 17876
rect 17865 17867 17923 17873
rect 17865 17864 17877 17867
rect 17552 17836 17877 17864
rect 17552 17824 17558 17836
rect 17865 17833 17877 17836
rect 17911 17833 17923 17867
rect 17865 17827 17923 17833
rect 17954 17824 17960 17876
rect 18012 17864 18018 17876
rect 18141 17867 18199 17873
rect 18141 17864 18153 17867
rect 18012 17836 18153 17864
rect 18012 17824 18018 17836
rect 18141 17833 18153 17836
rect 18187 17864 18199 17867
rect 18693 17867 18751 17873
rect 18693 17864 18705 17867
rect 18187 17836 18705 17864
rect 18187 17833 18199 17836
rect 18141 17827 18199 17833
rect 18693 17833 18705 17836
rect 18739 17833 18751 17867
rect 18693 17827 18751 17833
rect 19978 17824 19984 17876
rect 20036 17864 20042 17876
rect 20073 17867 20131 17873
rect 20073 17864 20085 17867
rect 20036 17836 20085 17864
rect 20036 17824 20042 17836
rect 20073 17833 20085 17836
rect 20119 17864 20131 17867
rect 20625 17867 20683 17873
rect 20625 17864 20637 17867
rect 20119 17836 20637 17864
rect 20119 17833 20131 17836
rect 20073 17827 20131 17833
rect 20625 17833 20637 17836
rect 20671 17833 20683 17867
rect 20898 17864 20904 17876
rect 20859 17836 20904 17864
rect 20625 17827 20683 17833
rect 20898 17824 20904 17836
rect 20956 17824 20962 17876
rect 21358 17864 21364 17876
rect 21319 17836 21364 17864
rect 21358 17824 21364 17836
rect 21416 17824 21422 17876
rect 22278 17864 22284 17876
rect 22239 17836 22284 17864
rect 22278 17824 22284 17836
rect 22336 17824 22342 17876
rect 24946 17824 24952 17876
rect 25004 17864 25010 17876
rect 25041 17867 25099 17873
rect 25041 17864 25053 17867
rect 25004 17836 25053 17864
rect 25004 17824 25010 17836
rect 25041 17833 25053 17836
rect 25087 17833 25099 17867
rect 25041 17827 25099 17833
rect 25590 17824 25596 17876
rect 25648 17864 25654 17876
rect 25777 17867 25835 17873
rect 25777 17864 25789 17867
rect 25648 17836 25789 17864
rect 25648 17824 25654 17836
rect 25777 17833 25789 17836
rect 25823 17833 25835 17867
rect 25777 17827 25835 17833
rect 8110 17796 8116 17808
rect 7392 17768 8116 17796
rect 1762 17728 1768 17740
rect 1723 17700 1768 17728
rect 1762 17688 1768 17700
rect 1820 17688 1826 17740
rect 1854 17688 1860 17740
rect 1912 17728 1918 17740
rect 2032 17731 2090 17737
rect 2032 17728 2044 17731
rect 1912 17700 2044 17728
rect 1912 17688 1918 17700
rect 2032 17697 2044 17700
rect 2078 17728 2090 17731
rect 2590 17728 2596 17740
rect 2078 17700 2596 17728
rect 2078 17697 2090 17700
rect 2032 17691 2090 17697
rect 2590 17688 2596 17700
rect 2648 17688 2654 17740
rect 3881 17731 3939 17737
rect 3881 17697 3893 17731
rect 3927 17728 3939 17731
rect 4062 17728 4068 17740
rect 3927 17700 4068 17728
rect 3927 17697 3939 17700
rect 3881 17691 3939 17697
rect 4062 17688 4068 17700
rect 4120 17688 4126 17740
rect 5629 17731 5687 17737
rect 5629 17697 5641 17731
rect 5675 17728 5687 17731
rect 6270 17728 6276 17740
rect 5675 17700 6276 17728
rect 5675 17697 5687 17700
rect 5629 17691 5687 17697
rect 6270 17688 6276 17700
rect 6328 17688 6334 17740
rect 6914 17688 6920 17740
rect 6972 17728 6978 17740
rect 7392 17737 7420 17768
rect 8110 17756 8116 17768
rect 8168 17756 8174 17808
rect 10137 17799 10195 17805
rect 10137 17765 10149 17799
rect 10183 17796 10195 17799
rect 10778 17796 10784 17808
rect 10183 17768 10784 17796
rect 10183 17765 10195 17768
rect 10137 17759 10195 17765
rect 10778 17756 10784 17768
rect 10836 17756 10842 17808
rect 13814 17796 13820 17808
rect 13727 17768 13820 17796
rect 13814 17756 13820 17768
rect 13872 17796 13878 17808
rect 14734 17796 14740 17808
rect 13872 17768 14740 17796
rect 13872 17756 13878 17768
rect 14734 17756 14740 17768
rect 14792 17756 14798 17808
rect 18046 17756 18052 17808
rect 18104 17796 18110 17808
rect 19061 17799 19119 17805
rect 19061 17796 19073 17799
rect 18104 17768 19073 17796
rect 18104 17756 18110 17768
rect 19061 17765 19073 17768
rect 19107 17765 19119 17799
rect 19061 17759 19119 17765
rect 19150 17756 19156 17808
rect 19208 17756 19214 17808
rect 20714 17756 20720 17808
rect 20772 17796 20778 17808
rect 21910 17796 21916 17808
rect 20772 17768 21916 17796
rect 20772 17756 20778 17768
rect 21910 17756 21916 17768
rect 21968 17756 21974 17808
rect 22833 17799 22891 17805
rect 22833 17765 22845 17799
rect 22879 17796 22891 17799
rect 23750 17796 23756 17808
rect 22879 17768 23756 17796
rect 22879 17765 22891 17768
rect 22833 17759 22891 17765
rect 23750 17756 23756 17768
rect 23808 17796 23814 17808
rect 25409 17799 25467 17805
rect 25409 17796 25421 17799
rect 23808 17768 25421 17796
rect 23808 17756 23814 17768
rect 25409 17765 25421 17768
rect 25455 17765 25467 17799
rect 25409 17759 25467 17765
rect 7650 17737 7656 17740
rect 7193 17731 7251 17737
rect 7193 17728 7205 17731
rect 6972 17700 7205 17728
rect 6972 17688 6978 17700
rect 7193 17697 7205 17700
rect 7239 17697 7251 17731
rect 7193 17691 7251 17697
rect 7377 17731 7435 17737
rect 7377 17697 7389 17731
rect 7423 17697 7435 17731
rect 7644 17728 7656 17737
rect 7611 17700 7656 17728
rect 7377 17691 7435 17697
rect 7644 17691 7656 17700
rect 7650 17688 7656 17691
rect 7708 17688 7714 17740
rect 9858 17728 9864 17740
rect 9819 17700 9864 17728
rect 9858 17688 9864 17700
rect 9916 17688 9922 17740
rect 11422 17737 11428 17740
rect 11416 17728 11428 17737
rect 11335 17700 11428 17728
rect 11416 17691 11428 17700
rect 11480 17728 11486 17740
rect 12250 17728 12256 17740
rect 11480 17700 12256 17728
rect 11422 17688 11428 17691
rect 11480 17688 11486 17700
rect 12250 17688 12256 17700
rect 12308 17688 12314 17740
rect 13446 17688 13452 17740
rect 13504 17728 13510 17740
rect 13725 17731 13783 17737
rect 13725 17728 13737 17731
rect 13504 17700 13737 17728
rect 13504 17688 13510 17700
rect 13725 17697 13737 17700
rect 13771 17697 13783 17731
rect 13725 17691 13783 17697
rect 15381 17731 15439 17737
rect 15381 17697 15393 17731
rect 15427 17728 15439 17731
rect 15562 17728 15568 17740
rect 15427 17700 15568 17728
rect 15427 17697 15439 17700
rect 15381 17691 15439 17697
rect 15562 17688 15568 17700
rect 15620 17688 15626 17740
rect 16298 17728 16304 17740
rect 16259 17700 16304 17728
rect 16298 17688 16304 17700
rect 16356 17688 16362 17740
rect 16752 17731 16810 17737
rect 16752 17697 16764 17731
rect 16798 17728 16810 17731
rect 17678 17728 17684 17740
rect 16798 17700 17684 17728
rect 16798 17697 16810 17700
rect 16752 17691 16810 17697
rect 17678 17688 17684 17700
rect 17736 17688 17742 17740
rect 19168 17728 19196 17756
rect 21269 17731 21327 17737
rect 19168 17700 19288 17728
rect 4430 17620 4436 17672
rect 4488 17660 4494 17672
rect 5721 17663 5779 17669
rect 5721 17660 5733 17663
rect 4488 17632 5733 17660
rect 4488 17620 4494 17632
rect 5721 17629 5733 17632
rect 5767 17629 5779 17663
rect 5902 17660 5908 17672
rect 5863 17632 5908 17660
rect 5721 17623 5779 17629
rect 5902 17620 5908 17632
rect 5960 17620 5966 17672
rect 10686 17620 10692 17672
rect 10744 17660 10750 17672
rect 11054 17660 11060 17672
rect 10744 17632 11060 17660
rect 10744 17620 10750 17632
rect 11054 17620 11060 17632
rect 11112 17660 11118 17672
rect 11149 17663 11207 17669
rect 11149 17660 11161 17663
rect 11112 17632 11161 17660
rect 11112 17620 11118 17632
rect 11149 17629 11161 17632
rect 11195 17629 11207 17663
rect 11149 17623 11207 17629
rect 13262 17620 13268 17672
rect 13320 17660 13326 17672
rect 13909 17663 13967 17669
rect 13909 17660 13921 17663
rect 13320 17632 13921 17660
rect 13320 17620 13326 17632
rect 13909 17629 13921 17632
rect 13955 17629 13967 17663
rect 13909 17623 13967 17629
rect 16390 17620 16396 17672
rect 16448 17660 16454 17672
rect 16485 17663 16543 17669
rect 16485 17660 16497 17663
rect 16448 17632 16497 17660
rect 16448 17620 16454 17632
rect 16485 17629 16497 17632
rect 16531 17629 16543 17663
rect 16485 17623 16543 17629
rect 18782 17620 18788 17672
rect 18840 17660 18846 17672
rect 19260 17669 19288 17700
rect 21269 17697 21281 17731
rect 21315 17728 21327 17731
rect 21542 17728 21548 17740
rect 21315 17700 21548 17728
rect 21315 17697 21327 17700
rect 21269 17691 21327 17697
rect 21542 17688 21548 17700
rect 21600 17688 21606 17740
rect 24394 17728 24400 17740
rect 24355 17700 24400 17728
rect 24394 17688 24400 17700
rect 24452 17688 24458 17740
rect 24489 17731 24547 17737
rect 24489 17697 24501 17731
rect 24535 17728 24547 17731
rect 24762 17728 24768 17740
rect 24535 17700 24768 17728
rect 24535 17697 24547 17700
rect 24489 17691 24547 17697
rect 24762 17688 24768 17700
rect 24820 17688 24826 17740
rect 19153 17663 19211 17669
rect 19153 17660 19165 17663
rect 18840 17632 19165 17660
rect 18840 17620 18846 17632
rect 19153 17629 19165 17632
rect 19199 17629 19211 17663
rect 19153 17623 19211 17629
rect 19245 17663 19303 17669
rect 19245 17629 19257 17663
rect 19291 17660 19303 17663
rect 19705 17663 19763 17669
rect 19705 17660 19717 17663
rect 19291 17632 19717 17660
rect 19291 17629 19303 17632
rect 19245 17623 19303 17629
rect 19705 17629 19717 17632
rect 19751 17629 19763 17663
rect 21450 17660 21456 17672
rect 21411 17632 21456 17660
rect 19705 17623 19763 17629
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 22186 17620 22192 17672
rect 22244 17660 22250 17672
rect 22922 17660 22928 17672
rect 22244 17632 22928 17660
rect 22244 17620 22250 17632
rect 22922 17620 22928 17632
rect 22980 17620 22986 17672
rect 23014 17620 23020 17672
rect 23072 17660 23078 17672
rect 23842 17660 23848 17672
rect 23072 17632 23848 17660
rect 23072 17620 23078 17632
rect 23842 17620 23848 17632
rect 23900 17620 23906 17672
rect 24670 17660 24676 17672
rect 24631 17632 24676 17660
rect 24670 17620 24676 17632
rect 24728 17620 24734 17672
rect 8754 17592 8760 17604
rect 8715 17564 8760 17592
rect 8754 17552 8760 17564
rect 8812 17552 8818 17604
rect 12802 17592 12808 17604
rect 12084 17564 12808 17592
rect 12084 17536 12112 17564
rect 12802 17552 12808 17564
rect 12860 17552 12866 17604
rect 13354 17592 13360 17604
rect 13315 17564 13360 17592
rect 13354 17552 13360 17564
rect 13412 17552 13418 17604
rect 22002 17552 22008 17604
rect 22060 17592 22066 17604
rect 22465 17595 22523 17601
rect 22465 17592 22477 17595
rect 22060 17564 22477 17592
rect 22060 17552 22066 17564
rect 22465 17561 22477 17564
rect 22511 17561 22523 17595
rect 22465 17555 22523 17561
rect 1670 17524 1676 17536
rect 1631 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 3234 17484 3240 17536
rect 3292 17524 3298 17536
rect 3421 17527 3479 17533
rect 3421 17524 3433 17527
rect 3292 17496 3433 17524
rect 3292 17484 3298 17496
rect 3421 17493 3433 17496
rect 3467 17493 3479 17527
rect 3421 17487 3479 17493
rect 6362 17484 6368 17536
rect 6420 17524 6426 17536
rect 6457 17527 6515 17533
rect 6457 17524 6469 17527
rect 6420 17496 6469 17524
rect 6420 17484 6426 17496
rect 6457 17493 6469 17496
rect 6503 17493 6515 17527
rect 6457 17487 6515 17493
rect 7190 17484 7196 17536
rect 7248 17524 7254 17536
rect 9122 17524 9128 17536
rect 7248 17496 9128 17524
rect 7248 17484 7254 17496
rect 9122 17484 9128 17496
rect 9180 17484 9186 17536
rect 11057 17527 11115 17533
rect 11057 17493 11069 17527
rect 11103 17524 11115 17527
rect 11146 17524 11152 17536
rect 11103 17496 11152 17524
rect 11103 17493 11115 17496
rect 11057 17487 11115 17493
rect 11146 17484 11152 17496
rect 11204 17484 11210 17536
rect 12066 17484 12072 17536
rect 12124 17484 12130 17536
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 14826 17524 14832 17536
rect 14787 17496 14832 17524
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 18601 17527 18659 17533
rect 18601 17493 18613 17527
rect 18647 17524 18659 17527
rect 19058 17524 19064 17536
rect 18647 17496 19064 17524
rect 18647 17493 18659 17496
rect 18601 17487 18659 17493
rect 19058 17484 19064 17496
rect 19116 17484 19122 17536
rect 23753 17527 23811 17533
rect 23753 17493 23765 17527
rect 23799 17524 23811 17527
rect 23842 17524 23848 17536
rect 23799 17496 23848 17524
rect 23799 17493 23811 17496
rect 23753 17487 23811 17493
rect 23842 17484 23848 17496
rect 23900 17484 23906 17536
rect 24026 17524 24032 17536
rect 23987 17496 24032 17524
rect 24026 17484 24032 17496
rect 24084 17484 24090 17536
rect 25866 17484 25872 17536
rect 25924 17524 25930 17536
rect 26142 17524 26148 17536
rect 25924 17496 26148 17524
rect 25924 17484 25930 17496
rect 26142 17484 26148 17496
rect 26200 17484 26206 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 3602 17320 3608 17332
rect 3563 17292 3608 17320
rect 3602 17280 3608 17292
rect 3660 17280 3666 17332
rect 5905 17323 5963 17329
rect 5905 17320 5917 17323
rect 4080 17292 5917 17320
rect 2590 17212 2596 17264
rect 2648 17252 2654 17264
rect 2961 17255 3019 17261
rect 2961 17252 2973 17255
rect 2648 17224 2973 17252
rect 2648 17212 2654 17224
rect 2961 17221 2973 17224
rect 3007 17252 3019 17255
rect 4080 17252 4108 17292
rect 5905 17289 5917 17292
rect 5951 17320 5963 17323
rect 6546 17320 6552 17332
rect 5951 17292 6552 17320
rect 5951 17289 5963 17292
rect 5905 17283 5963 17289
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 6641 17323 6699 17329
rect 6641 17289 6653 17323
rect 6687 17320 6699 17323
rect 6730 17320 6736 17332
rect 6687 17292 6736 17320
rect 6687 17289 6699 17292
rect 6641 17283 6699 17289
rect 6730 17280 6736 17292
rect 6788 17280 6794 17332
rect 7561 17323 7619 17329
rect 7561 17289 7573 17323
rect 7607 17320 7619 17323
rect 7650 17320 7656 17332
rect 7607 17292 7656 17320
rect 7607 17289 7619 17292
rect 7561 17283 7619 17289
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 11606 17320 11612 17332
rect 9916 17292 11612 17320
rect 9916 17280 9922 17292
rect 11606 17280 11612 17292
rect 11664 17280 11670 17332
rect 13446 17280 13452 17332
rect 13504 17320 13510 17332
rect 14090 17320 14096 17332
rect 13504 17292 14096 17320
rect 13504 17280 13510 17292
rect 14090 17280 14096 17292
rect 14148 17280 14154 17332
rect 14553 17323 14611 17329
rect 14553 17289 14565 17323
rect 14599 17320 14611 17323
rect 14734 17320 14740 17332
rect 14599 17292 14740 17320
rect 14599 17289 14611 17292
rect 14553 17283 14611 17289
rect 14734 17280 14740 17292
rect 14792 17280 14798 17332
rect 17770 17320 17776 17332
rect 17731 17292 17776 17320
rect 17770 17280 17776 17292
rect 17828 17280 17834 17332
rect 18046 17280 18052 17332
rect 18104 17320 18110 17332
rect 18325 17323 18383 17329
rect 18325 17320 18337 17323
rect 18104 17292 18337 17320
rect 18104 17280 18110 17292
rect 18325 17289 18337 17292
rect 18371 17289 18383 17323
rect 18782 17320 18788 17332
rect 18743 17292 18788 17320
rect 18325 17283 18383 17289
rect 18782 17280 18788 17292
rect 18840 17280 18846 17332
rect 18874 17280 18880 17332
rect 18932 17320 18938 17332
rect 23477 17323 23535 17329
rect 23477 17320 23489 17323
rect 18932 17292 23489 17320
rect 18932 17280 18938 17292
rect 23477 17289 23489 17292
rect 23523 17289 23535 17323
rect 23658 17320 23664 17332
rect 23619 17292 23664 17320
rect 23477 17283 23535 17289
rect 4430 17252 4436 17264
rect 3007 17224 4108 17252
rect 4391 17224 4436 17252
rect 3007 17221 3019 17224
rect 2961 17215 3019 17221
rect 4430 17212 4436 17224
rect 4488 17212 4494 17264
rect 11333 17255 11391 17261
rect 11333 17221 11345 17255
rect 11379 17252 11391 17255
rect 11422 17252 11428 17264
rect 11379 17224 11428 17252
rect 11379 17221 11391 17224
rect 11333 17215 11391 17221
rect 11422 17212 11428 17224
rect 11480 17212 11486 17264
rect 14645 17255 14703 17261
rect 14645 17221 14657 17255
rect 14691 17252 14703 17255
rect 15657 17255 15715 17261
rect 15657 17252 15669 17255
rect 14691 17224 15669 17252
rect 14691 17221 14703 17224
rect 14645 17215 14703 17221
rect 15657 17221 15669 17224
rect 15703 17221 15715 17255
rect 15657 17215 15715 17221
rect 17313 17255 17371 17261
rect 17313 17221 17325 17255
rect 17359 17252 17371 17255
rect 17678 17252 17684 17264
rect 17359 17224 17684 17252
rect 17359 17221 17371 17224
rect 17313 17215 17371 17221
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 2501 17187 2559 17193
rect 2501 17184 2513 17187
rect 1811 17156 2513 17184
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 2501 17153 2513 17156
rect 2547 17184 2559 17187
rect 2682 17184 2688 17196
rect 2547 17156 2688 17184
rect 2547 17153 2559 17156
rect 2501 17147 2559 17153
rect 2682 17144 2688 17156
rect 2740 17144 2746 17196
rect 4154 17144 4160 17196
rect 4212 17184 4218 17196
rect 4338 17184 4344 17196
rect 4212 17156 4344 17184
rect 4212 17144 4218 17156
rect 4338 17144 4344 17156
rect 4396 17184 4402 17196
rect 4525 17187 4583 17193
rect 4525 17184 4537 17187
rect 4396 17156 4537 17184
rect 4396 17144 4402 17156
rect 4525 17153 4537 17156
rect 4571 17153 4583 17187
rect 4525 17147 4583 17153
rect 6086 17144 6092 17196
rect 6144 17184 6150 17196
rect 6546 17184 6552 17196
rect 6144 17156 6552 17184
rect 6144 17144 6150 17156
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 7009 17187 7067 17193
rect 7009 17153 7021 17187
rect 7055 17184 7067 17187
rect 7742 17184 7748 17196
rect 7055 17156 7748 17184
rect 7055 17153 7067 17156
rect 7009 17147 7067 17153
rect 7742 17144 7748 17156
rect 7800 17144 7806 17196
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17184 7987 17187
rect 10137 17187 10195 17193
rect 7975 17156 8156 17184
rect 7975 17153 7987 17156
rect 7929 17147 7987 17153
rect 3234 17116 3240 17128
rect 2240 17088 3240 17116
rect 2240 16992 2268 17088
rect 3234 17076 3240 17088
rect 3292 17076 3298 17128
rect 3421 17119 3479 17125
rect 3421 17085 3433 17119
rect 3467 17116 3479 17119
rect 8018 17116 8024 17128
rect 3467 17088 4108 17116
rect 7979 17088 8024 17116
rect 3467 17085 3479 17088
rect 3421 17079 3479 17085
rect 2317 17051 2375 17057
rect 2317 17017 2329 17051
rect 2363 17048 2375 17051
rect 2958 17048 2964 17060
rect 2363 17020 2964 17048
rect 2363 17017 2375 17020
rect 2317 17011 2375 17017
rect 2958 17008 2964 17020
rect 3016 17048 3022 17060
rect 3329 17051 3387 17057
rect 3329 17048 3341 17051
rect 3016 17020 3341 17048
rect 3016 17008 3022 17020
rect 3329 17017 3341 17020
rect 3375 17017 3387 17051
rect 3329 17011 3387 17017
rect 4080 16992 4108 17088
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 8128 17116 8156 17156
rect 10137 17153 10149 17187
rect 10183 17184 10195 17187
rect 10686 17184 10692 17196
rect 10183 17156 10692 17184
rect 10183 17153 10195 17156
rect 10137 17147 10195 17153
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 10870 17184 10876 17196
rect 10831 17156 10876 17184
rect 10870 17144 10876 17156
rect 10928 17144 10934 17196
rect 14826 17144 14832 17196
rect 14884 17184 14890 17196
rect 15102 17184 15108 17196
rect 14884 17156 15108 17184
rect 14884 17144 14890 17156
rect 15102 17144 15108 17156
rect 15160 17144 15166 17196
rect 15197 17187 15255 17193
rect 15197 17153 15209 17187
rect 15243 17153 15255 17187
rect 15197 17147 15255 17153
rect 8288 17119 8346 17125
rect 8288 17116 8300 17119
rect 8128 17088 8300 17116
rect 8288 17085 8300 17088
rect 8334 17116 8346 17119
rect 8754 17116 8760 17128
rect 8334 17088 8760 17116
rect 8334 17085 8346 17088
rect 8288 17079 8346 17085
rect 8754 17076 8760 17088
rect 8812 17076 8818 17128
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 11112 17088 12449 17116
rect 11112 17076 11118 17088
rect 12437 17085 12449 17088
rect 12483 17116 12495 17119
rect 12986 17116 12992 17128
rect 12483 17088 12992 17116
rect 12483 17085 12495 17088
rect 12437 17079 12495 17085
rect 12986 17076 12992 17088
rect 13044 17076 13050 17128
rect 14642 17076 14648 17128
rect 14700 17116 14706 17128
rect 15212 17116 15240 17147
rect 14700 17088 15240 17116
rect 15672 17116 15700 17215
rect 17678 17212 17684 17224
rect 17736 17212 17742 17264
rect 22922 17212 22928 17264
rect 22980 17252 22986 17264
rect 23017 17255 23075 17261
rect 23017 17252 23029 17255
rect 22980 17224 23029 17252
rect 22980 17212 22986 17224
rect 23017 17221 23029 17224
rect 23063 17221 23075 17255
rect 23017 17215 23075 17221
rect 15838 17144 15844 17196
rect 15896 17184 15902 17196
rect 16117 17187 16175 17193
rect 16117 17184 16129 17187
rect 15896 17156 16129 17184
rect 15896 17144 15902 17156
rect 16117 17153 16129 17156
rect 16163 17184 16175 17187
rect 16761 17187 16819 17193
rect 16761 17184 16773 17187
rect 16163 17156 16773 17184
rect 16163 17153 16175 17156
rect 16117 17147 16175 17153
rect 16761 17153 16773 17156
rect 16807 17153 16819 17187
rect 16761 17147 16819 17153
rect 16577 17119 16635 17125
rect 16577 17116 16589 17119
rect 15672 17088 16589 17116
rect 14700 17076 14706 17088
rect 16577 17085 16589 17088
rect 16623 17085 16635 17119
rect 18966 17116 18972 17128
rect 18927 17088 18972 17116
rect 16577 17079 16635 17085
rect 18966 17076 18972 17088
rect 19024 17076 19030 17128
rect 19058 17076 19064 17128
rect 19116 17116 19122 17128
rect 19242 17125 19248 17128
rect 19225 17119 19248 17125
rect 19225 17116 19237 17119
rect 19116 17088 19237 17116
rect 19116 17076 19122 17088
rect 19225 17085 19237 17088
rect 19225 17079 19248 17085
rect 19242 17076 19248 17079
rect 19300 17076 19306 17128
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 19536 17088 21189 17116
rect 4792 17051 4850 17057
rect 4792 17017 4804 17051
rect 4838 17048 4850 17051
rect 4982 17048 4988 17060
rect 4838 17020 4988 17048
rect 4838 17017 4850 17020
rect 4792 17011 4850 17017
rect 4982 17008 4988 17020
rect 5040 17008 5046 17060
rect 9769 17051 9827 17057
rect 9769 17017 9781 17051
rect 9815 17048 9827 17051
rect 10597 17051 10655 17057
rect 10597 17048 10609 17051
rect 9815 17020 10609 17048
rect 9815 17017 9827 17020
rect 9769 17011 9827 17017
rect 10597 17017 10609 17020
rect 10643 17048 10655 17051
rect 10778 17048 10784 17060
rect 10643 17020 10784 17048
rect 10643 17017 10655 17020
rect 10597 17011 10655 17017
rect 10778 17008 10784 17020
rect 10836 17008 10842 17060
rect 12704 17051 12762 17057
rect 12704 17017 12716 17051
rect 12750 17017 12762 17051
rect 15010 17048 15016 17060
rect 14971 17020 15016 17048
rect 12704 17011 12762 17017
rect 1857 16983 1915 16989
rect 1857 16949 1869 16983
rect 1903 16980 1915 16983
rect 1946 16980 1952 16992
rect 1903 16952 1952 16980
rect 1903 16949 1915 16952
rect 1857 16943 1915 16949
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 2222 16980 2228 16992
rect 2183 16952 2228 16980
rect 2222 16940 2228 16952
rect 2280 16940 2286 16992
rect 4062 16980 4068 16992
rect 4023 16952 4068 16980
rect 4062 16940 4068 16952
rect 4120 16940 4126 16992
rect 6270 16980 6276 16992
rect 6231 16952 6276 16980
rect 6270 16940 6276 16952
rect 6328 16940 6334 16992
rect 9398 16980 9404 16992
rect 9359 16952 9404 16980
rect 9398 16940 9404 16952
rect 9456 16940 9462 16992
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 10192 16952 10241 16980
rect 10192 16940 10198 16952
rect 10229 16949 10241 16952
rect 10275 16949 10287 16983
rect 12158 16980 12164 16992
rect 12119 16952 12164 16980
rect 10229 16943 10287 16949
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 12719 16980 12747 17011
rect 15010 17008 15016 17020
rect 15068 17008 15074 17060
rect 16298 17008 16304 17060
rect 16356 17048 16362 17060
rect 16669 17051 16727 17057
rect 16669 17048 16681 17051
rect 16356 17020 16681 17048
rect 16356 17008 16362 17020
rect 16669 17017 16681 17020
rect 16715 17017 16727 17051
rect 18984 17048 19012 17076
rect 19536 17060 19564 17088
rect 21177 17085 21189 17088
rect 21223 17116 21235 17119
rect 21726 17116 21732 17128
rect 21223 17088 21732 17116
rect 21223 17085 21235 17088
rect 21177 17079 21235 17085
rect 21726 17076 21732 17088
rect 21784 17076 21790 17128
rect 22646 17076 22652 17128
rect 22704 17116 22710 17128
rect 22922 17116 22928 17128
rect 22704 17088 22928 17116
rect 22704 17076 22710 17088
rect 22922 17076 22928 17088
rect 22980 17076 22986 17128
rect 23032 17116 23060 17215
rect 23492 17184 23520 17283
rect 23658 17280 23664 17292
rect 23716 17280 23722 17332
rect 25406 17212 25412 17264
rect 25464 17252 25470 17264
rect 26142 17252 26148 17264
rect 25464 17224 26148 17252
rect 25464 17212 25470 17224
rect 26142 17212 26148 17224
rect 26200 17212 26206 17264
rect 24121 17187 24179 17193
rect 24121 17184 24133 17187
rect 23492 17156 24133 17184
rect 24121 17153 24133 17156
rect 24167 17153 24179 17187
rect 24121 17147 24179 17153
rect 24213 17187 24271 17193
rect 24213 17153 24225 17187
rect 24259 17184 24271 17187
rect 24670 17184 24676 17196
rect 24259 17156 24676 17184
rect 24259 17153 24271 17156
rect 24213 17147 24271 17153
rect 24228 17116 24256 17147
rect 24670 17144 24676 17156
rect 24728 17184 24734 17196
rect 25041 17187 25099 17193
rect 25041 17184 25053 17187
rect 24728 17156 25053 17184
rect 24728 17144 24734 17156
rect 25041 17153 25053 17156
rect 25087 17153 25099 17187
rect 25041 17147 25099 17153
rect 25222 17116 25228 17128
rect 23032 17088 24256 17116
rect 25183 17088 25228 17116
rect 25222 17076 25228 17088
rect 25280 17116 25286 17128
rect 25961 17119 26019 17125
rect 25961 17116 25973 17119
rect 25280 17088 25973 17116
rect 25280 17076 25286 17088
rect 25961 17085 25973 17088
rect 26007 17085 26019 17119
rect 25961 17079 26019 17085
rect 19518 17048 19524 17060
rect 18984 17020 19524 17048
rect 16669 17011 16727 17017
rect 19518 17008 19524 17020
rect 19576 17008 19582 17060
rect 21450 17057 21456 17060
rect 20993 17051 21051 17057
rect 20993 17017 21005 17051
rect 21039 17048 21051 17051
rect 21444 17048 21456 17057
rect 21039 17020 21456 17048
rect 21039 17017 21051 17020
rect 20993 17011 21051 17017
rect 21444 17011 21456 17020
rect 21508 17048 21514 17060
rect 21910 17048 21916 17060
rect 21508 17020 21916 17048
rect 12584 16952 12747 16980
rect 13817 16983 13875 16989
rect 12584 16940 12590 16952
rect 13817 16949 13829 16983
rect 13863 16980 13875 16983
rect 13998 16980 14004 16992
rect 13863 16952 14004 16980
rect 13863 16949 13875 16952
rect 13817 16943 13875 16949
rect 13998 16940 14004 16952
rect 14056 16940 14062 16992
rect 16206 16980 16212 16992
rect 16167 16952 16212 16980
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 20349 16983 20407 16989
rect 20349 16949 20361 16983
rect 20395 16980 20407 16983
rect 21008 16980 21036 17011
rect 21450 17008 21456 17011
rect 21508 17008 21514 17020
rect 21910 17008 21916 17020
rect 21968 17008 21974 17060
rect 25406 17008 25412 17060
rect 25464 17048 25470 17060
rect 25501 17051 25559 17057
rect 25501 17048 25513 17051
rect 25464 17020 25513 17048
rect 25464 17008 25470 17020
rect 25501 17017 25513 17020
rect 25547 17017 25559 17051
rect 25501 17011 25559 17017
rect 20395 16952 21036 16980
rect 22557 16983 22615 16989
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 22557 16949 22569 16983
rect 22603 16980 22615 16983
rect 22646 16980 22652 16992
rect 22603 16952 22652 16980
rect 22603 16949 22615 16952
rect 22557 16943 22615 16949
rect 22646 16940 22652 16952
rect 22704 16940 22710 16992
rect 23842 16940 23848 16992
rect 23900 16980 23906 16992
rect 24026 16980 24032 16992
rect 23900 16952 24032 16980
rect 23900 16940 23906 16952
rect 24026 16940 24032 16952
rect 24084 16940 24090 16992
rect 24670 16980 24676 16992
rect 24631 16952 24676 16980
rect 24670 16940 24676 16952
rect 24728 16940 24734 16992
rect 25590 16940 25596 16992
rect 25648 16980 25654 16992
rect 26329 16983 26387 16989
rect 26329 16980 26341 16983
rect 25648 16952 26341 16980
rect 25648 16940 25654 16952
rect 26329 16949 26341 16952
rect 26375 16949 26387 16983
rect 26329 16943 26387 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1765 16779 1823 16785
rect 1765 16745 1777 16779
rect 1811 16776 1823 16779
rect 2222 16776 2228 16788
rect 1811 16748 2228 16776
rect 1811 16745 1823 16748
rect 1765 16739 1823 16745
rect 2222 16736 2228 16748
rect 2280 16736 2286 16788
rect 3605 16779 3663 16785
rect 3605 16776 3617 16779
rect 2700 16748 3617 16776
rect 2133 16711 2191 16717
rect 2133 16708 2145 16711
rect 1780 16680 2145 16708
rect 1780 16652 1808 16680
rect 2133 16677 2145 16680
rect 2179 16708 2191 16711
rect 2700 16708 2728 16748
rect 3605 16745 3617 16748
rect 3651 16745 3663 16779
rect 3605 16739 3663 16745
rect 3694 16736 3700 16788
rect 3752 16776 3758 16788
rect 4249 16779 4307 16785
rect 4249 16776 4261 16779
rect 3752 16748 4261 16776
rect 3752 16736 3758 16748
rect 4249 16745 4261 16748
rect 4295 16745 4307 16779
rect 5166 16776 5172 16788
rect 5127 16748 5172 16776
rect 4249 16739 4307 16745
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 5350 16736 5356 16788
rect 5408 16776 5414 16788
rect 5629 16779 5687 16785
rect 5629 16776 5641 16779
rect 5408 16748 5641 16776
rect 5408 16736 5414 16748
rect 5629 16745 5641 16748
rect 5675 16745 5687 16779
rect 5629 16739 5687 16745
rect 6178 16736 6184 16788
rect 6236 16736 6242 16788
rect 6914 16776 6920 16788
rect 6875 16748 6920 16776
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 8386 16736 8392 16788
rect 8444 16776 8450 16788
rect 8849 16779 8907 16785
rect 8849 16776 8861 16779
rect 8444 16748 8861 16776
rect 8444 16736 8450 16748
rect 8849 16745 8861 16748
rect 8895 16776 8907 16779
rect 10134 16776 10140 16788
rect 8895 16748 10140 16776
rect 8895 16745 8907 16748
rect 8849 16739 8907 16745
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 10689 16779 10747 16785
rect 10689 16745 10701 16779
rect 10735 16776 10747 16779
rect 10870 16776 10876 16788
rect 10735 16748 10876 16776
rect 10735 16745 10747 16748
rect 10689 16739 10747 16745
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 12897 16779 12955 16785
rect 12897 16745 12909 16779
rect 12943 16776 12955 16779
rect 13722 16776 13728 16788
rect 12943 16748 13728 16776
rect 12943 16745 12955 16748
rect 12897 16739 12955 16745
rect 13722 16736 13728 16748
rect 13780 16736 13786 16788
rect 14642 16776 14648 16788
rect 14603 16748 14648 16776
rect 14642 16736 14648 16748
rect 14700 16736 14706 16788
rect 15010 16776 15016 16788
rect 14971 16748 15016 16776
rect 15010 16736 15016 16748
rect 15068 16736 15074 16788
rect 16850 16736 16856 16788
rect 16908 16776 16914 16788
rect 17681 16779 17739 16785
rect 17681 16776 17693 16779
rect 16908 16748 17693 16776
rect 16908 16736 16914 16748
rect 17681 16745 17693 16748
rect 17727 16745 17739 16779
rect 17681 16739 17739 16745
rect 18601 16779 18659 16785
rect 18601 16745 18613 16779
rect 18647 16776 18659 16779
rect 18785 16779 18843 16785
rect 18785 16776 18797 16779
rect 18647 16748 18797 16776
rect 18647 16745 18659 16748
rect 18601 16739 18659 16745
rect 18785 16745 18797 16748
rect 18831 16776 18843 16779
rect 19058 16776 19064 16788
rect 18831 16748 19064 16776
rect 18831 16745 18843 16748
rect 18785 16739 18843 16745
rect 19058 16736 19064 16748
rect 19116 16736 19122 16788
rect 19153 16779 19211 16785
rect 19153 16745 19165 16779
rect 19199 16776 19211 16779
rect 19242 16776 19248 16788
rect 19199 16748 19248 16776
rect 19199 16745 19211 16748
rect 19153 16739 19211 16745
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 19978 16736 19984 16788
rect 20036 16776 20042 16788
rect 20257 16779 20315 16785
rect 20257 16776 20269 16779
rect 20036 16748 20269 16776
rect 20036 16736 20042 16748
rect 20257 16745 20269 16748
rect 20303 16776 20315 16779
rect 20533 16779 20591 16785
rect 20533 16776 20545 16779
rect 20303 16748 20545 16776
rect 20303 16745 20315 16748
rect 20257 16739 20315 16745
rect 20533 16745 20545 16748
rect 20579 16745 20591 16779
rect 20533 16739 20591 16745
rect 20901 16779 20959 16785
rect 20901 16745 20913 16779
rect 20947 16745 20959 16779
rect 20901 16739 20959 16745
rect 2866 16708 2872 16720
rect 2179 16680 2728 16708
rect 2827 16680 2872 16708
rect 2179 16677 2191 16680
rect 2133 16671 2191 16677
rect 2866 16668 2872 16680
rect 2924 16668 2930 16720
rect 3326 16708 3332 16720
rect 3287 16680 3332 16708
rect 3326 16668 3332 16680
rect 3384 16668 3390 16720
rect 6196 16708 6224 16736
rect 6454 16708 6460 16720
rect 6196 16680 6460 16708
rect 6454 16668 6460 16680
rect 6512 16668 6518 16720
rect 7650 16708 7656 16720
rect 7611 16680 7656 16708
rect 7650 16668 7656 16680
rect 7708 16708 7714 16720
rect 8754 16708 8760 16720
rect 7708 16680 8760 16708
rect 7708 16668 7714 16680
rect 8754 16668 8760 16680
rect 8812 16708 8818 16720
rect 9217 16711 9275 16717
rect 9217 16708 9229 16711
rect 8812 16680 9229 16708
rect 8812 16668 8818 16680
rect 9217 16677 9229 16680
rect 9263 16677 9275 16711
rect 16298 16708 16304 16720
rect 9217 16671 9275 16677
rect 15488 16680 16304 16708
rect 1762 16600 1768 16652
rect 1820 16600 1826 16652
rect 3050 16600 3056 16652
rect 3108 16640 3114 16652
rect 3602 16640 3608 16652
rect 3108 16612 3608 16640
rect 3108 16600 3114 16612
rect 3602 16600 3608 16612
rect 3660 16600 3666 16652
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 5537 16643 5595 16649
rect 5537 16609 5549 16643
rect 5583 16640 5595 16643
rect 6178 16640 6184 16652
rect 5583 16612 6184 16640
rect 5583 16609 5595 16612
rect 5537 16603 5595 16609
rect 2222 16572 2228 16584
rect 2183 16544 2228 16572
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 2406 16572 2412 16584
rect 2367 16544 2412 16572
rect 2406 16532 2412 16544
rect 2464 16532 2470 16584
rect 4080 16572 4108 16603
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 6546 16640 6552 16652
rect 6288 16612 6552 16640
rect 4154 16572 4160 16584
rect 4080 16544 4160 16572
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 5813 16575 5871 16581
rect 5813 16541 5825 16575
rect 5859 16572 5871 16575
rect 5994 16572 6000 16584
rect 5859 16544 6000 16572
rect 5859 16541 5871 16544
rect 5813 16535 5871 16541
rect 5994 16532 6000 16544
rect 6052 16532 6058 16584
rect 6288 16572 6316 16612
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 6730 16640 6736 16652
rect 6691 16612 6736 16640
rect 6730 16600 6736 16612
rect 6788 16640 6794 16652
rect 7285 16643 7343 16649
rect 7285 16640 7297 16643
rect 6788 16612 7297 16640
rect 6788 16600 6794 16612
rect 7285 16609 7297 16612
rect 7331 16609 7343 16643
rect 8202 16640 8208 16652
rect 8163 16612 8208 16640
rect 7285 16603 7343 16609
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 9858 16640 9864 16652
rect 9819 16612 9864 16640
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 10137 16643 10195 16649
rect 10137 16609 10149 16643
rect 10183 16640 10195 16643
rect 10962 16640 10968 16652
rect 10183 16612 10968 16640
rect 10183 16609 10195 16612
rect 10137 16603 10195 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 11422 16649 11428 16652
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 11112 16612 11161 16640
rect 11112 16600 11118 16612
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 11416 16640 11428 16649
rect 11383 16612 11428 16640
rect 11149 16603 11207 16609
rect 11416 16603 11428 16612
rect 11422 16600 11428 16603
rect 11480 16600 11486 16652
rect 11790 16600 11796 16652
rect 11848 16640 11854 16652
rect 13173 16643 13231 16649
rect 13173 16640 13185 16643
rect 11848 16612 13185 16640
rect 11848 16600 11854 16612
rect 13173 16609 13185 16612
rect 13219 16640 13231 16643
rect 13262 16640 13268 16652
rect 13219 16612 13268 16640
rect 13219 16609 13231 16612
rect 13173 16603 13231 16609
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 13538 16600 13544 16652
rect 13596 16640 13602 16652
rect 15488 16649 15516 16680
rect 16298 16668 16304 16680
rect 16356 16708 16362 16720
rect 16758 16708 16764 16720
rect 16356 16680 16764 16708
rect 16356 16668 16362 16680
rect 16758 16668 16764 16680
rect 16816 16668 16822 16720
rect 17589 16711 17647 16717
rect 17589 16677 17601 16711
rect 17635 16708 17647 16711
rect 19613 16711 19671 16717
rect 19613 16708 19625 16711
rect 17635 16680 19625 16708
rect 17635 16677 17647 16680
rect 17589 16671 17647 16677
rect 19613 16677 19625 16680
rect 19659 16708 19671 16711
rect 20916 16708 20944 16739
rect 21266 16736 21272 16788
rect 21324 16776 21330 16788
rect 21361 16779 21419 16785
rect 21361 16776 21373 16779
rect 21324 16748 21373 16776
rect 21324 16736 21330 16748
rect 21361 16745 21373 16748
rect 21407 16745 21419 16779
rect 21910 16776 21916 16788
rect 21871 16748 21916 16776
rect 21361 16739 21419 16745
rect 21910 16736 21916 16748
rect 21968 16736 21974 16788
rect 22557 16779 22615 16785
rect 22557 16745 22569 16779
rect 22603 16776 22615 16779
rect 23014 16776 23020 16788
rect 22603 16748 23020 16776
rect 22603 16745 22615 16748
rect 22557 16739 22615 16745
rect 23014 16736 23020 16748
rect 23072 16776 23078 16788
rect 24121 16779 24179 16785
rect 24121 16776 24133 16779
rect 23072 16748 24133 16776
rect 23072 16736 23078 16748
rect 24121 16745 24133 16748
rect 24167 16745 24179 16779
rect 24854 16776 24860 16788
rect 24815 16748 24860 16776
rect 24121 16739 24179 16745
rect 24854 16736 24860 16748
rect 24912 16736 24918 16788
rect 25130 16776 25136 16788
rect 25091 16748 25136 16776
rect 25130 16736 25136 16748
rect 25188 16736 25194 16788
rect 25501 16711 25559 16717
rect 25501 16708 25513 16711
rect 19659 16680 20944 16708
rect 22756 16680 25513 16708
rect 19659 16677 19671 16680
rect 19613 16671 19671 16677
rect 15746 16649 15752 16652
rect 13725 16643 13783 16649
rect 13725 16640 13737 16643
rect 13596 16612 13737 16640
rect 13596 16600 13602 16612
rect 13725 16609 13737 16612
rect 13771 16609 13783 16643
rect 13725 16603 13783 16609
rect 15473 16643 15531 16649
rect 15473 16609 15485 16643
rect 15519 16609 15531 16643
rect 15740 16640 15752 16649
rect 15707 16612 15752 16640
rect 15473 16603 15531 16609
rect 15740 16603 15752 16612
rect 15746 16600 15752 16603
rect 15804 16600 15810 16652
rect 18049 16643 18107 16649
rect 18049 16640 18061 16643
rect 17696 16612 18061 16640
rect 8297 16575 8355 16581
rect 8297 16572 8309 16575
rect 6104 16544 6316 16572
rect 8220 16544 8309 16572
rect 4798 16464 4804 16516
rect 4856 16504 4862 16516
rect 6104 16504 6132 16544
rect 8220 16516 8248 16544
rect 8297 16541 8309 16544
rect 8343 16541 8355 16575
rect 8297 16535 8355 16541
rect 8481 16575 8539 16581
rect 8481 16541 8493 16575
rect 8527 16572 8539 16575
rect 8938 16572 8944 16584
rect 8527 16544 8944 16572
rect 8527 16541 8539 16544
rect 8481 16535 8539 16541
rect 8938 16532 8944 16544
rect 8996 16532 9002 16584
rect 12894 16532 12900 16584
rect 12952 16572 12958 16584
rect 13817 16575 13875 16581
rect 13817 16572 13829 16575
rect 12952 16544 13829 16572
rect 12952 16532 12958 16544
rect 13817 16541 13829 16544
rect 13863 16541 13875 16575
rect 13817 16535 13875 16541
rect 13906 16532 13912 16584
rect 13964 16572 13970 16584
rect 13964 16544 14009 16572
rect 13964 16532 13970 16544
rect 17218 16532 17224 16584
rect 17276 16572 17282 16584
rect 17696 16572 17724 16612
rect 18049 16609 18061 16612
rect 18095 16609 18107 16643
rect 18049 16603 18107 16609
rect 18141 16643 18199 16649
rect 18141 16609 18153 16643
rect 18187 16609 18199 16643
rect 18601 16643 18659 16649
rect 18601 16640 18613 16643
rect 18141 16603 18199 16609
rect 18340 16612 18613 16640
rect 17276 16544 17724 16572
rect 17276 16532 17282 16544
rect 17770 16532 17776 16584
rect 17828 16572 17834 16584
rect 18156 16572 18184 16603
rect 18340 16581 18368 16612
rect 18601 16609 18613 16612
rect 18647 16609 18659 16643
rect 18601 16603 18659 16609
rect 20622 16600 20628 16652
rect 20680 16640 20686 16652
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 20680 16612 21281 16640
rect 20680 16600 20686 16612
rect 21269 16609 21281 16612
rect 21315 16609 21327 16643
rect 21269 16603 21327 16609
rect 21726 16600 21732 16652
rect 21784 16640 21790 16652
rect 22370 16640 22376 16652
rect 21784 16612 22376 16640
rect 21784 16600 21790 16612
rect 22370 16600 22376 16612
rect 22428 16640 22434 16652
rect 22756 16649 22784 16680
rect 25501 16677 25513 16680
rect 25547 16708 25559 16711
rect 25590 16708 25596 16720
rect 25547 16680 25596 16708
rect 25547 16677 25559 16680
rect 25501 16671 25559 16677
rect 25590 16668 25596 16680
rect 25648 16668 25654 16720
rect 23014 16649 23020 16652
rect 22741 16643 22799 16649
rect 22741 16640 22753 16643
rect 22428 16612 22753 16640
rect 22428 16600 22434 16612
rect 22741 16609 22753 16612
rect 22787 16609 22799 16643
rect 23008 16640 23020 16649
rect 22975 16612 23020 16640
rect 22741 16603 22799 16609
rect 23008 16603 23020 16612
rect 23014 16600 23020 16603
rect 23072 16600 23078 16652
rect 24946 16640 24952 16652
rect 24907 16612 24952 16640
rect 24946 16600 24952 16612
rect 25004 16600 25010 16652
rect 17828 16544 18184 16572
rect 18325 16575 18383 16581
rect 17828 16532 17834 16544
rect 18325 16541 18337 16575
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 4856 16476 6132 16504
rect 4856 16464 4862 16476
rect 8202 16464 8208 16516
rect 8260 16464 8266 16516
rect 16853 16507 16911 16513
rect 16853 16473 16865 16507
rect 16899 16504 16911 16507
rect 17034 16504 17040 16516
rect 16899 16476 17040 16504
rect 16899 16473 16911 16476
rect 16853 16467 16911 16473
rect 17034 16464 17040 16476
rect 17092 16504 17098 16516
rect 18340 16504 18368 16535
rect 18506 16532 18512 16584
rect 18564 16572 18570 16584
rect 19702 16572 19708 16584
rect 18564 16544 19708 16572
rect 18564 16532 18570 16544
rect 19702 16532 19708 16544
rect 19760 16532 19766 16584
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16541 19855 16575
rect 19797 16535 19855 16541
rect 20533 16575 20591 16581
rect 20533 16541 20545 16575
rect 20579 16572 20591 16575
rect 21082 16572 21088 16584
rect 20579 16544 21088 16572
rect 20579 16541 20591 16544
rect 20533 16535 20591 16541
rect 17092 16476 18368 16504
rect 17092 16464 17098 16476
rect 19150 16464 19156 16516
rect 19208 16504 19214 16516
rect 19245 16507 19303 16513
rect 19245 16504 19257 16507
rect 19208 16476 19257 16504
rect 19208 16464 19214 16476
rect 19245 16473 19257 16476
rect 19291 16473 19303 16507
rect 19245 16467 19303 16473
rect 19334 16464 19340 16516
rect 19392 16504 19398 16516
rect 19812 16504 19840 16535
rect 21082 16532 21088 16544
rect 21140 16572 21146 16584
rect 21453 16575 21511 16581
rect 21453 16572 21465 16575
rect 21140 16544 21465 16572
rect 21140 16532 21146 16544
rect 21453 16541 21465 16544
rect 21499 16541 21511 16575
rect 21453 16535 21511 16541
rect 22002 16532 22008 16584
rect 22060 16572 22066 16584
rect 22462 16572 22468 16584
rect 22060 16544 22468 16572
rect 22060 16532 22066 16544
rect 22462 16532 22468 16544
rect 22520 16532 22526 16584
rect 19392 16476 19840 16504
rect 19392 16464 19398 16476
rect 23842 16464 23848 16516
rect 23900 16504 23906 16516
rect 24118 16504 24124 16516
rect 23900 16476 24124 16504
rect 23900 16464 23906 16476
rect 24118 16464 24124 16476
rect 24176 16464 24182 16516
rect 1673 16439 1731 16445
rect 1673 16405 1685 16439
rect 1719 16436 1731 16439
rect 1762 16436 1768 16448
rect 1719 16408 1768 16436
rect 1719 16405 1731 16408
rect 1673 16399 1731 16405
rect 1762 16396 1768 16408
rect 1820 16396 1826 16448
rect 4709 16439 4767 16445
rect 4709 16405 4721 16439
rect 4755 16436 4767 16439
rect 4982 16436 4988 16448
rect 4755 16408 4988 16436
rect 4755 16405 4767 16408
rect 4709 16399 4767 16405
rect 4982 16396 4988 16408
rect 5040 16396 5046 16448
rect 5077 16439 5135 16445
rect 5077 16405 5089 16439
rect 5123 16436 5135 16439
rect 5166 16436 5172 16448
rect 5123 16408 5172 16436
rect 5123 16405 5135 16408
rect 5077 16399 5135 16405
rect 5166 16396 5172 16408
rect 5224 16396 5230 16448
rect 6270 16436 6276 16448
rect 6183 16408 6276 16436
rect 6270 16396 6276 16408
rect 6328 16436 6334 16448
rect 7006 16436 7012 16448
rect 6328 16408 7012 16436
rect 6328 16396 6334 16408
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 7098 16396 7104 16448
rect 7156 16436 7162 16448
rect 7837 16439 7895 16445
rect 7837 16436 7849 16439
rect 7156 16408 7849 16436
rect 7156 16396 7162 16408
rect 7837 16405 7849 16408
rect 7883 16405 7895 16439
rect 11054 16436 11060 16448
rect 11015 16408 11060 16436
rect 7837 16399 7895 16405
rect 11054 16396 11060 16408
rect 11112 16396 11118 16448
rect 12526 16436 12532 16448
rect 12487 16408 12532 16436
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 13357 16439 13415 16445
rect 13357 16405 13369 16439
rect 13403 16436 13415 16439
rect 13446 16436 13452 16448
rect 13403 16408 13452 16436
rect 13403 16405 13415 16408
rect 13357 16399 13415 16405
rect 13446 16396 13452 16408
rect 13504 16396 13510 16448
rect 17221 16439 17279 16445
rect 17221 16405 17233 16439
rect 17267 16436 17279 16439
rect 17402 16436 17408 16448
rect 17267 16408 17408 16436
rect 17267 16405 17279 16408
rect 17221 16399 17279 16405
rect 17402 16396 17408 16408
rect 17460 16396 17466 16448
rect 20622 16436 20628 16448
rect 20583 16408 20628 16436
rect 20622 16396 20628 16408
rect 20680 16396 20686 16448
rect 22462 16396 22468 16448
rect 22520 16436 22526 16448
rect 24489 16439 24547 16445
rect 24489 16436 24501 16439
rect 22520 16408 24501 16436
rect 22520 16396 22526 16408
rect 24489 16405 24501 16408
rect 24535 16436 24547 16439
rect 24854 16436 24860 16448
rect 24535 16408 24860 16436
rect 24535 16405 24547 16408
rect 24489 16399 24547 16405
rect 24854 16396 24860 16408
rect 24912 16396 24918 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2225 16235 2283 16241
rect 2225 16201 2237 16235
rect 2271 16232 2283 16235
rect 2406 16232 2412 16244
rect 2271 16204 2412 16232
rect 2271 16201 2283 16204
rect 2225 16195 2283 16201
rect 2406 16192 2412 16204
rect 2464 16232 2470 16244
rect 2682 16232 2688 16244
rect 2464 16204 2688 16232
rect 2464 16192 2470 16204
rect 2682 16192 2688 16204
rect 2740 16192 2746 16244
rect 4338 16192 4344 16244
rect 4396 16232 4402 16244
rect 4433 16235 4491 16241
rect 4433 16232 4445 16235
rect 4396 16204 4445 16232
rect 4396 16192 4402 16204
rect 4433 16201 4445 16204
rect 4479 16201 4491 16235
rect 4433 16195 4491 16201
rect 5077 16235 5135 16241
rect 5077 16201 5089 16235
rect 5123 16232 5135 16235
rect 5350 16232 5356 16244
rect 5123 16204 5356 16232
rect 5123 16201 5135 16204
rect 5077 16195 5135 16201
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 6549 16235 6607 16241
rect 6549 16232 6561 16235
rect 6052 16204 6561 16232
rect 6052 16192 6058 16204
rect 6549 16201 6561 16204
rect 6595 16201 6607 16235
rect 6549 16195 6607 16201
rect 7837 16235 7895 16241
rect 7837 16201 7849 16235
rect 7883 16232 7895 16235
rect 8110 16232 8116 16244
rect 7883 16204 8116 16232
rect 7883 16201 7895 16204
rect 7837 16195 7895 16201
rect 8110 16192 8116 16204
rect 8168 16192 8174 16244
rect 8938 16192 8944 16244
rect 8996 16232 9002 16244
rect 9309 16235 9367 16241
rect 9309 16232 9321 16235
rect 8996 16204 9321 16232
rect 8996 16192 9002 16204
rect 9309 16201 9321 16204
rect 9355 16201 9367 16235
rect 9674 16232 9680 16244
rect 9635 16204 9680 16232
rect 9309 16195 9367 16201
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 10321 16235 10379 16241
rect 10321 16201 10333 16235
rect 10367 16232 10379 16235
rect 11422 16232 11428 16244
rect 10367 16204 11428 16232
rect 10367 16201 10379 16204
rect 10321 16195 10379 16201
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 13538 16232 13544 16244
rect 13499 16204 13544 16232
rect 13538 16192 13544 16204
rect 13596 16192 13602 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 14001 16235 14059 16241
rect 14001 16232 14013 16235
rect 13872 16204 14013 16232
rect 13872 16192 13878 16204
rect 14001 16201 14013 16204
rect 14047 16201 14059 16235
rect 17034 16232 17040 16244
rect 16995 16204 17040 16232
rect 14001 16195 14059 16201
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 19702 16192 19708 16244
rect 19760 16232 19766 16244
rect 20441 16235 20499 16241
rect 20441 16232 20453 16235
rect 19760 16204 20453 16232
rect 19760 16192 19766 16204
rect 20441 16201 20453 16204
rect 20487 16201 20499 16235
rect 20441 16195 20499 16201
rect 21266 16192 21272 16244
rect 21324 16232 21330 16244
rect 21453 16235 21511 16241
rect 21453 16232 21465 16235
rect 21324 16204 21465 16232
rect 21324 16192 21330 16204
rect 21453 16201 21465 16204
rect 21499 16201 21511 16235
rect 21453 16195 21511 16201
rect 22005 16235 22063 16241
rect 22005 16201 22017 16235
rect 22051 16232 22063 16235
rect 22186 16232 22192 16244
rect 22051 16204 22192 16232
rect 22051 16201 22063 16204
rect 22005 16195 22063 16201
rect 22186 16192 22192 16204
rect 22244 16192 22250 16244
rect 23661 16235 23719 16241
rect 22296 16204 23152 16232
rect 2869 16167 2927 16173
rect 2869 16133 2881 16167
rect 2915 16164 2927 16167
rect 2958 16164 2964 16176
rect 2915 16136 2964 16164
rect 2915 16133 2927 16136
rect 2869 16127 2927 16133
rect 2958 16124 2964 16136
rect 3016 16124 3022 16176
rect 5442 16124 5448 16176
rect 5500 16164 5506 16176
rect 6178 16164 6184 16176
rect 5500 16136 6184 16164
rect 5500 16124 5506 16136
rect 6178 16124 6184 16136
rect 6236 16124 6242 16176
rect 10689 16167 10747 16173
rect 10689 16133 10701 16167
rect 10735 16164 10747 16167
rect 12158 16164 12164 16176
rect 10735 16136 12164 16164
rect 10735 16133 10747 16136
rect 10689 16127 10747 16133
rect 2774 16056 2780 16108
rect 2832 16096 2838 16108
rect 3421 16099 3479 16105
rect 3421 16096 3433 16099
rect 2832 16068 3433 16096
rect 2832 16056 2838 16068
rect 3421 16065 3433 16068
rect 3467 16065 3479 16099
rect 3421 16059 3479 16065
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 5994 16096 6000 16108
rect 5859 16068 6000 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11348 16105 11376 16136
rect 12158 16124 12164 16136
rect 12216 16164 12222 16176
rect 12526 16164 12532 16176
rect 12216 16136 12532 16164
rect 12216 16124 12222 16136
rect 12526 16124 12532 16136
rect 12584 16124 12590 16176
rect 19978 16164 19984 16176
rect 19939 16136 19984 16164
rect 19978 16124 19984 16136
rect 20036 16124 20042 16176
rect 21913 16167 21971 16173
rect 21913 16164 21925 16167
rect 21836 16136 21925 16164
rect 11241 16099 11299 16105
rect 11241 16096 11253 16099
rect 11112 16068 11253 16096
rect 11112 16056 11118 16068
rect 11241 16065 11253 16068
rect 11287 16065 11299 16099
rect 11241 16059 11299 16065
rect 11333 16099 11391 16105
rect 11333 16065 11345 16099
rect 11379 16065 11391 16099
rect 11882 16096 11888 16108
rect 11795 16068 11888 16096
rect 11333 16059 11391 16065
rect 11882 16056 11888 16068
rect 11940 16096 11946 16108
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 11940 16068 13001 16096
rect 11940 16056 11946 16068
rect 12989 16065 13001 16068
rect 13035 16096 13047 16099
rect 13538 16096 13544 16108
rect 13035 16068 13544 16096
rect 13035 16065 13047 16068
rect 12989 16059 13047 16065
rect 13538 16056 13544 16068
rect 13596 16096 13602 16108
rect 13906 16096 13912 16108
rect 13596 16068 13912 16096
rect 13596 16056 13602 16068
rect 13906 16056 13912 16068
rect 13964 16096 13970 16108
rect 14366 16096 14372 16108
rect 13964 16068 14372 16096
rect 13964 16056 13970 16068
rect 14366 16056 14372 16068
rect 14424 16096 14430 16108
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 14424 16068 14565 16096
rect 14424 16056 14430 16068
rect 14553 16065 14565 16068
rect 14599 16096 14611 16099
rect 15013 16099 15071 16105
rect 15013 16096 15025 16099
rect 14599 16068 15025 16096
rect 14599 16065 14611 16068
rect 14553 16059 14611 16065
rect 15013 16065 15025 16068
rect 15059 16065 15071 16099
rect 15013 16059 15071 16065
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16096 15531 16099
rect 15746 16096 15752 16108
rect 15519 16068 15752 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 15746 16056 15752 16068
rect 15804 16096 15810 16108
rect 16209 16099 16267 16105
rect 16209 16096 16221 16099
rect 15804 16068 16221 16096
rect 15804 16056 15810 16068
rect 16209 16065 16221 16068
rect 16255 16096 16267 16099
rect 16666 16096 16672 16108
rect 16255 16068 16672 16096
rect 16255 16065 16267 16068
rect 16209 16059 16267 16065
rect 16666 16056 16672 16068
rect 16724 16056 16730 16108
rect 21082 16096 21088 16108
rect 21043 16068 21088 16096
rect 21082 16056 21088 16068
rect 21140 16056 21146 16108
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1762 16028 1768 16040
rect 1443 16000 1768 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 2866 15988 2872 16040
rect 2924 16028 2930 16040
rect 3329 16031 3387 16037
rect 3329 16028 3341 16031
rect 2924 16000 3341 16028
rect 2924 15988 2930 16000
rect 3329 15997 3341 16000
rect 3375 15997 3387 16031
rect 3329 15991 3387 15997
rect 4617 16031 4675 16037
rect 4617 15997 4629 16031
rect 4663 16028 4675 16031
rect 4798 16028 4804 16040
rect 4663 16000 4804 16028
rect 4663 15997 4675 16000
rect 4617 15991 4675 15997
rect 4798 15988 4804 16000
rect 4856 15988 4862 16040
rect 5166 15988 5172 16040
rect 5224 16028 5230 16040
rect 5629 16031 5687 16037
rect 5629 16028 5641 16031
rect 5224 16000 5641 16028
rect 5224 15988 5230 16000
rect 5629 15997 5641 16000
rect 5675 16028 5687 16031
rect 7098 16028 7104 16040
rect 5675 16000 7104 16028
rect 5675 15997 5687 16000
rect 5629 15991 5687 15997
rect 7098 15988 7104 16000
rect 7156 15988 7162 16040
rect 7926 16028 7932 16040
rect 7887 16000 7932 16028
rect 7926 15988 7932 16000
rect 7984 15988 7990 16040
rect 14458 16028 14464 16040
rect 14419 16000 14464 16028
rect 14458 15988 14464 16000
rect 14516 15988 14522 16040
rect 18046 16028 18052 16040
rect 18007 16000 18052 16028
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 1486 15920 1492 15972
rect 1544 15960 1550 15972
rect 1673 15963 1731 15969
rect 1673 15960 1685 15963
rect 1544 15932 1685 15960
rect 1544 15920 1550 15932
rect 1673 15929 1685 15932
rect 1719 15929 1731 15963
rect 1673 15923 1731 15929
rect 2406 15920 2412 15972
rect 2464 15960 2470 15972
rect 7469 15963 7527 15969
rect 2464 15932 6960 15960
rect 2464 15920 2470 15932
rect 3237 15895 3295 15901
rect 3237 15861 3249 15895
rect 3283 15892 3295 15895
rect 3326 15892 3332 15904
rect 3283 15864 3332 15892
rect 3283 15861 3295 15864
rect 3237 15855 3295 15861
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 4154 15892 4160 15904
rect 4115 15864 4160 15892
rect 4154 15852 4160 15864
rect 4212 15852 4218 15904
rect 5169 15895 5227 15901
rect 5169 15861 5181 15895
rect 5215 15892 5227 15895
rect 5258 15892 5264 15904
rect 5215 15864 5264 15892
rect 5215 15861 5227 15864
rect 5169 15855 5227 15861
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 5537 15895 5595 15901
rect 5537 15861 5549 15895
rect 5583 15892 5595 15895
rect 6270 15892 6276 15904
rect 5583 15864 6276 15892
rect 5583 15861 5595 15864
rect 5537 15855 5595 15861
rect 6270 15852 6276 15864
rect 6328 15852 6334 15904
rect 6638 15852 6644 15904
rect 6696 15892 6702 15904
rect 6825 15895 6883 15901
rect 6825 15892 6837 15895
rect 6696 15864 6837 15892
rect 6696 15852 6702 15864
rect 6825 15861 6837 15864
rect 6871 15861 6883 15895
rect 6932 15892 6960 15932
rect 7469 15929 7481 15963
rect 7515 15960 7527 15963
rect 8196 15963 8254 15969
rect 8196 15960 8208 15963
rect 7515 15932 8208 15960
rect 7515 15929 7527 15932
rect 7469 15923 7527 15929
rect 8196 15929 8208 15932
rect 8242 15960 8254 15963
rect 9398 15960 9404 15972
rect 8242 15932 9404 15960
rect 8242 15929 8254 15932
rect 8196 15923 8254 15929
rect 9398 15920 9404 15932
rect 9456 15920 9462 15972
rect 10134 15920 10140 15972
rect 10192 15960 10198 15972
rect 11330 15960 11336 15972
rect 10192 15932 11336 15960
rect 10192 15920 10198 15932
rect 11330 15920 11336 15932
rect 11388 15920 11394 15972
rect 12253 15963 12311 15969
rect 12253 15929 12265 15963
rect 12299 15960 12311 15963
rect 12618 15960 12624 15972
rect 12299 15932 12624 15960
rect 12299 15929 12311 15932
rect 12253 15923 12311 15929
rect 12618 15920 12624 15932
rect 12676 15960 12682 15972
rect 12805 15963 12863 15969
rect 12676 15932 12756 15960
rect 12676 15920 12682 15932
rect 9030 15892 9036 15904
rect 6932 15864 9036 15892
rect 6825 15855 6883 15861
rect 9030 15852 9036 15864
rect 9088 15852 9094 15904
rect 10778 15892 10784 15904
rect 10739 15864 10784 15892
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 11146 15892 11152 15904
rect 11107 15864 11152 15892
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 12728 15892 12756 15932
rect 12805 15929 12817 15963
rect 12851 15960 12863 15963
rect 13078 15960 13084 15972
rect 12851 15932 13084 15960
rect 12851 15929 12863 15932
rect 12805 15923 12863 15929
rect 13078 15920 13084 15932
rect 13136 15920 13142 15972
rect 13909 15963 13967 15969
rect 13909 15929 13921 15963
rect 13955 15960 13967 15963
rect 14369 15963 14427 15969
rect 14369 15960 14381 15963
rect 13955 15932 14381 15960
rect 13955 15929 13967 15932
rect 13909 15923 13967 15929
rect 14369 15929 14381 15932
rect 14415 15960 14427 15963
rect 14550 15960 14556 15972
rect 14415 15932 14556 15960
rect 14415 15929 14427 15932
rect 14369 15923 14427 15929
rect 14550 15920 14556 15932
rect 14608 15920 14614 15972
rect 17218 15920 17224 15972
rect 17276 15960 17282 15972
rect 17313 15963 17371 15969
rect 17313 15960 17325 15963
rect 17276 15932 17325 15960
rect 17276 15920 17282 15932
rect 17313 15929 17325 15932
rect 17359 15929 17371 15963
rect 17313 15923 17371 15929
rect 18138 15920 18144 15972
rect 18196 15960 18202 15972
rect 18294 15963 18352 15969
rect 18294 15960 18306 15963
rect 18196 15932 18306 15960
rect 18196 15920 18202 15932
rect 18294 15929 18306 15932
rect 18340 15929 18352 15963
rect 18294 15923 18352 15929
rect 20349 15963 20407 15969
rect 20349 15929 20361 15963
rect 20395 15960 20407 15963
rect 20809 15963 20867 15969
rect 20809 15960 20821 15963
rect 20395 15932 20821 15960
rect 20395 15929 20407 15932
rect 20349 15923 20407 15929
rect 20809 15929 20821 15932
rect 20855 15960 20867 15963
rect 21082 15960 21088 15972
rect 20855 15932 21088 15960
rect 20855 15929 20867 15932
rect 20809 15923 20867 15929
rect 21082 15920 21088 15932
rect 21140 15920 21146 15972
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 12492 15864 12537 15892
rect 12728 15864 12909 15892
rect 12492 15852 12498 15864
rect 12897 15861 12909 15864
rect 12943 15892 12955 15895
rect 12986 15892 12992 15904
rect 12943 15864 12992 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 12986 15852 12992 15864
rect 13044 15852 13050 15904
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 13630 15892 13636 15904
rect 13412 15864 13636 15892
rect 13412 15852 13418 15864
rect 13630 15852 13636 15864
rect 13688 15852 13694 15904
rect 15562 15892 15568 15904
rect 15523 15864 15568 15892
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 15930 15892 15936 15904
rect 15891 15864 15936 15892
rect 15930 15852 15936 15864
rect 15988 15852 15994 15904
rect 16025 15895 16083 15901
rect 16025 15861 16037 15895
rect 16071 15892 16083 15895
rect 16114 15892 16120 15904
rect 16071 15864 16120 15892
rect 16071 15861 16083 15864
rect 16025 15855 16083 15861
rect 16114 15852 16120 15864
rect 16172 15852 16178 15904
rect 16666 15892 16672 15904
rect 16627 15864 16672 15892
rect 16666 15852 16672 15864
rect 16724 15852 16730 15904
rect 17770 15892 17776 15904
rect 17731 15864 17776 15892
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 19429 15895 19487 15901
rect 19429 15861 19441 15895
rect 19475 15892 19487 15895
rect 20254 15892 20260 15904
rect 19475 15864 20260 15892
rect 19475 15861 19487 15864
rect 19429 15855 19487 15861
rect 20254 15852 20260 15864
rect 20312 15852 20318 15904
rect 20898 15892 20904 15904
rect 20859 15864 20904 15892
rect 20898 15852 20904 15864
rect 20956 15852 20962 15904
rect 21836 15892 21864 16136
rect 21913 16133 21925 16136
rect 21959 16164 21971 16167
rect 22296 16164 22324 16204
rect 23014 16164 23020 16176
rect 21959 16136 22324 16164
rect 22572 16136 23020 16164
rect 21959 16133 21971 16136
rect 21913 16127 21971 16133
rect 22572 16108 22600 16136
rect 23014 16124 23020 16136
rect 23072 16124 23078 16176
rect 23124 16164 23152 16204
rect 23661 16201 23673 16235
rect 23707 16232 23719 16235
rect 23750 16232 23756 16244
rect 23707 16204 23756 16232
rect 23707 16201 23719 16204
rect 23661 16195 23719 16201
rect 23750 16192 23756 16204
rect 23808 16192 23814 16244
rect 24946 16232 24952 16244
rect 24907 16204 24952 16232
rect 24946 16192 24952 16204
rect 25004 16192 25010 16244
rect 25409 16235 25467 16241
rect 25409 16201 25421 16235
rect 25455 16232 25467 16235
rect 25498 16232 25504 16244
rect 25455 16204 25504 16232
rect 25455 16201 25467 16204
rect 25409 16195 25467 16201
rect 25498 16192 25504 16204
rect 25556 16192 25562 16244
rect 25590 16192 25596 16244
rect 25648 16232 25654 16244
rect 26145 16235 26203 16241
rect 26145 16232 26157 16235
rect 25648 16204 26157 16232
rect 25648 16192 25654 16204
rect 26145 16201 26157 16204
rect 26191 16201 26203 16235
rect 26145 16195 26203 16201
rect 26234 16164 26240 16176
rect 23124 16136 26240 16164
rect 26234 16124 26240 16136
rect 26292 16124 26298 16176
rect 22554 16096 22560 16108
rect 22515 16068 22560 16096
rect 22554 16056 22560 16068
rect 22612 16056 22618 16108
rect 22738 16056 22744 16108
rect 22796 16056 22802 16108
rect 24210 16096 24216 16108
rect 24171 16068 24216 16096
rect 24210 16056 24216 16068
rect 24268 16056 24274 16108
rect 22186 15988 22192 16040
rect 22244 16028 22250 16040
rect 22756 16028 22784 16056
rect 22244 16000 22784 16028
rect 23109 16031 23167 16037
rect 22244 15988 22250 16000
rect 23109 15997 23121 16031
rect 23155 16028 23167 16031
rect 25222 16028 25228 16040
rect 23155 16000 24256 16028
rect 25183 16000 25228 16028
rect 23155 15997 23167 16000
rect 23109 15991 23167 15997
rect 24121 15963 24179 15969
rect 24121 15960 24133 15963
rect 23492 15932 24133 15960
rect 22373 15895 22431 15901
rect 22373 15892 22385 15895
rect 21836 15864 22385 15892
rect 22373 15861 22385 15864
rect 22419 15861 22431 15895
rect 22373 15855 22431 15861
rect 22462 15852 22468 15904
rect 22520 15892 22526 15904
rect 22520 15864 22565 15892
rect 22520 15852 22526 15864
rect 23106 15852 23112 15904
rect 23164 15892 23170 15904
rect 23492 15901 23520 15932
rect 24121 15929 24133 15932
rect 24167 15929 24179 15963
rect 24121 15923 24179 15929
rect 23477 15895 23535 15901
rect 23477 15892 23489 15895
rect 23164 15864 23489 15892
rect 23164 15852 23170 15864
rect 23477 15861 23489 15864
rect 23523 15861 23535 15895
rect 23477 15855 23535 15861
rect 24029 15895 24087 15901
rect 24029 15861 24041 15895
rect 24075 15892 24087 15895
rect 24228 15892 24256 16000
rect 25222 15988 25228 16000
rect 25280 16028 25286 16040
rect 25777 16031 25835 16037
rect 25777 16028 25789 16031
rect 25280 16000 25789 16028
rect 25280 15988 25286 16000
rect 25777 15997 25789 16000
rect 25823 15997 25835 16031
rect 25777 15991 25835 15997
rect 24762 15892 24768 15904
rect 24075 15864 24768 15892
rect 24075 15861 24087 15864
rect 24029 15855 24087 15861
rect 24762 15852 24768 15864
rect 24820 15852 24826 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1949 15691 2007 15697
rect 1949 15657 1961 15691
rect 1995 15688 2007 15691
rect 2222 15688 2228 15700
rect 1995 15660 2228 15688
rect 1995 15657 2007 15660
rect 1949 15651 2007 15657
rect 2222 15648 2228 15660
rect 2280 15688 2286 15700
rect 3329 15691 3387 15697
rect 3329 15688 3341 15691
rect 2280 15660 3341 15688
rect 2280 15648 2286 15660
rect 3329 15657 3341 15660
rect 3375 15657 3387 15691
rect 3329 15651 3387 15657
rect 4338 15648 4344 15700
rect 4396 15648 4402 15700
rect 8021 15691 8079 15697
rect 8021 15657 8033 15691
rect 8067 15688 8079 15691
rect 8202 15688 8208 15700
rect 8067 15660 8208 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 8389 15691 8447 15697
rect 8389 15657 8401 15691
rect 8435 15688 8447 15691
rect 8478 15688 8484 15700
rect 8435 15660 8484 15688
rect 8435 15657 8447 15660
rect 8389 15651 8447 15657
rect 8478 15648 8484 15660
rect 8536 15688 8542 15700
rect 9306 15688 9312 15700
rect 8536 15660 9312 15688
rect 8536 15648 8542 15660
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 12989 15691 13047 15697
rect 12989 15688 13001 15691
rect 11112 15660 13001 15688
rect 11112 15648 11118 15660
rect 12989 15657 13001 15660
rect 13035 15657 13047 15691
rect 13446 15688 13452 15700
rect 13407 15660 13452 15688
rect 12989 15651 13047 15657
rect 13446 15648 13452 15660
rect 13504 15648 13510 15700
rect 14366 15688 14372 15700
rect 14327 15660 14372 15688
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 16666 15688 16672 15700
rect 16627 15660 16672 15688
rect 16666 15648 16672 15660
rect 16724 15648 16730 15700
rect 17402 15688 17408 15700
rect 17363 15660 17408 15688
rect 17402 15648 17408 15660
rect 17460 15648 17466 15700
rect 17678 15688 17684 15700
rect 17639 15660 17684 15688
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 18138 15688 18144 15700
rect 18099 15660 18144 15688
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 18506 15688 18512 15700
rect 18467 15660 18512 15688
rect 18506 15648 18512 15660
rect 18564 15648 18570 15700
rect 19334 15648 19340 15700
rect 19392 15648 19398 15700
rect 19978 15688 19984 15700
rect 19939 15660 19984 15688
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 20806 15648 20812 15700
rect 20864 15688 20870 15700
rect 22097 15691 22155 15697
rect 20864 15660 21312 15688
rect 20864 15648 20870 15660
rect 2406 15620 2412 15632
rect 2367 15592 2412 15620
rect 2406 15580 2412 15592
rect 2464 15580 2470 15632
rect 4356 15620 4384 15648
rect 4080 15592 4384 15620
rect 2314 15552 2320 15564
rect 2275 15524 2320 15552
rect 2314 15512 2320 15524
rect 2372 15512 2378 15564
rect 2774 15512 2780 15564
rect 2832 15552 2838 15564
rect 4080 15561 4108 15592
rect 7650 15580 7656 15632
rect 7708 15620 7714 15632
rect 7929 15623 7987 15629
rect 7929 15620 7941 15623
rect 7708 15592 7941 15620
rect 7708 15580 7714 15592
rect 7929 15589 7941 15592
rect 7975 15620 7987 15623
rect 8938 15620 8944 15632
rect 7975 15592 8944 15620
rect 7975 15589 7987 15592
rect 7929 15583 7987 15589
rect 8938 15580 8944 15592
rect 8996 15580 9002 15632
rect 10689 15623 10747 15629
rect 10689 15589 10701 15623
rect 10735 15620 10747 15623
rect 11146 15620 11152 15632
rect 10735 15592 11152 15620
rect 10735 15589 10747 15592
rect 10689 15583 10747 15589
rect 11146 15580 11152 15592
rect 11204 15620 11210 15632
rect 12342 15620 12348 15632
rect 11204 15592 12348 15620
rect 11204 15580 11210 15592
rect 12342 15580 12348 15592
rect 12400 15580 12406 15632
rect 12434 15580 12440 15632
rect 12492 15620 12498 15632
rect 13357 15623 13415 15629
rect 13357 15620 13369 15623
rect 12492 15592 13369 15620
rect 12492 15580 12498 15592
rect 13357 15589 13369 15592
rect 13403 15620 13415 15623
rect 14737 15623 14795 15629
rect 14737 15620 14749 15623
rect 13403 15592 14749 15620
rect 13403 15589 13415 15592
rect 13357 15583 13415 15589
rect 14737 15589 14749 15592
rect 14783 15589 14795 15623
rect 14737 15583 14795 15589
rect 16390 15580 16396 15632
rect 16448 15620 16454 15632
rect 17420 15620 17448 15648
rect 16448 15592 17448 15620
rect 19352 15620 19380 15648
rect 20714 15620 20720 15632
rect 19352 15592 20720 15620
rect 16448 15580 16454 15592
rect 20714 15580 20720 15592
rect 20772 15580 20778 15632
rect 21284 15629 21312 15660
rect 22097 15657 22109 15691
rect 22143 15688 22155 15691
rect 22554 15688 22560 15700
rect 22143 15660 22560 15688
rect 22143 15657 22155 15660
rect 22097 15651 22155 15657
rect 22554 15648 22560 15660
rect 22612 15688 22618 15700
rect 23845 15691 23903 15697
rect 23845 15688 23857 15691
rect 22612 15660 23857 15688
rect 22612 15648 22618 15660
rect 23845 15657 23857 15660
rect 23891 15688 23903 15691
rect 24121 15691 24179 15697
rect 24121 15688 24133 15691
rect 23891 15660 24133 15688
rect 23891 15657 23903 15660
rect 23845 15651 23903 15657
rect 24121 15657 24133 15660
rect 24167 15688 24179 15691
rect 24210 15688 24216 15700
rect 24167 15660 24216 15688
rect 24167 15657 24179 15660
rect 24121 15651 24179 15657
rect 24210 15648 24216 15660
rect 24268 15688 24274 15700
rect 24489 15691 24547 15697
rect 24489 15688 24501 15691
rect 24268 15660 24501 15688
rect 24268 15648 24274 15660
rect 24489 15657 24501 15660
rect 24535 15657 24547 15691
rect 24489 15651 24547 15657
rect 25038 15648 25044 15700
rect 25096 15688 25102 15700
rect 25133 15691 25191 15697
rect 25133 15688 25145 15691
rect 25096 15660 25145 15688
rect 25096 15648 25102 15660
rect 25133 15657 25145 15660
rect 25179 15657 25191 15691
rect 25133 15651 25191 15657
rect 21269 15623 21327 15629
rect 21269 15589 21281 15623
rect 21315 15620 21327 15623
rect 21450 15620 21456 15632
rect 21315 15592 21456 15620
rect 21315 15589 21327 15592
rect 21269 15583 21327 15589
rect 21450 15580 21456 15592
rect 21508 15580 21514 15632
rect 22646 15580 22652 15632
rect 22704 15629 22710 15632
rect 22704 15623 22768 15629
rect 22704 15589 22722 15623
rect 22756 15589 22768 15623
rect 22704 15583 22768 15589
rect 22704 15580 22710 15583
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 2832 15524 4077 15552
rect 2832 15512 2838 15524
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 4154 15512 4160 15564
rect 4212 15552 4218 15564
rect 4321 15555 4379 15561
rect 4321 15552 4333 15555
rect 4212 15524 4333 15552
rect 4212 15512 4218 15524
rect 4321 15521 4333 15524
rect 4367 15521 4379 15555
rect 4321 15515 4379 15521
rect 6454 15512 6460 15564
rect 6512 15552 6518 15564
rect 6641 15555 6699 15561
rect 6641 15552 6653 15555
rect 6512 15524 6653 15552
rect 6512 15512 6518 15524
rect 6641 15521 6653 15524
rect 6687 15521 6699 15555
rect 6641 15515 6699 15521
rect 8386 15512 8392 15564
rect 8444 15552 8450 15564
rect 11054 15561 11060 15564
rect 8481 15555 8539 15561
rect 8481 15552 8493 15555
rect 8444 15524 8493 15552
rect 8444 15512 8450 15524
rect 8481 15521 8493 15524
rect 8527 15521 8539 15555
rect 11048 15552 11060 15561
rect 10967 15524 11060 15552
rect 8481 15515 8539 15521
rect 11048 15515 11060 15524
rect 11112 15552 11118 15564
rect 11882 15552 11888 15564
rect 11112 15524 11888 15552
rect 11054 15512 11060 15515
rect 11112 15512 11118 15524
rect 11882 15512 11888 15524
rect 11940 15512 11946 15564
rect 12894 15552 12900 15564
rect 12855 15524 12900 15552
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 14093 15555 14151 15561
rect 14093 15521 14105 15555
rect 14139 15552 14151 15555
rect 14458 15552 14464 15564
rect 14139 15524 14464 15552
rect 14139 15521 14151 15524
rect 14093 15515 14151 15521
rect 14458 15512 14464 15524
rect 14516 15512 14522 15564
rect 15556 15555 15614 15561
rect 15556 15521 15568 15555
rect 15602 15552 15614 15555
rect 15838 15552 15844 15564
rect 15602 15524 15844 15552
rect 15602 15521 15614 15524
rect 15556 15515 15614 15521
rect 15838 15512 15844 15524
rect 15896 15512 15902 15564
rect 17310 15512 17316 15564
rect 17368 15552 17374 15564
rect 18874 15561 18880 15564
rect 17497 15555 17555 15561
rect 17497 15552 17509 15555
rect 17368 15524 17509 15552
rect 17368 15512 17374 15524
rect 17497 15521 17509 15524
rect 17543 15521 17555 15555
rect 18868 15552 18880 15561
rect 18835 15524 18880 15552
rect 17497 15515 17555 15521
rect 18868 15515 18880 15524
rect 18874 15512 18880 15515
rect 18932 15512 18938 15564
rect 20530 15512 20536 15564
rect 20588 15552 20594 15564
rect 21361 15555 21419 15561
rect 21361 15552 21373 15555
rect 20588 15524 21373 15552
rect 20588 15512 20594 15524
rect 21361 15521 21373 15524
rect 21407 15521 21419 15555
rect 21361 15515 21419 15521
rect 22370 15512 22376 15564
rect 22428 15552 22434 15564
rect 22465 15555 22523 15561
rect 22465 15552 22477 15555
rect 22428 15524 22477 15552
rect 22428 15512 22434 15524
rect 22465 15521 22477 15524
rect 22511 15552 22523 15555
rect 23290 15552 23296 15564
rect 22511 15524 23296 15552
rect 22511 15521 22523 15524
rect 22465 15515 22523 15521
rect 23290 15512 23296 15524
rect 23348 15512 23354 15564
rect 25038 15552 25044 15564
rect 24999 15524 25044 15552
rect 25038 15512 25044 15524
rect 25096 15512 25102 15564
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15484 2559 15487
rect 2590 15484 2596 15496
rect 2547 15456 2596 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 2222 15376 2228 15428
rect 2280 15416 2286 15428
rect 2516 15416 2544 15447
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 3878 15484 3884 15496
rect 3839 15456 3884 15484
rect 3878 15444 3884 15456
rect 3936 15444 3942 15496
rect 6730 15484 6736 15496
rect 6691 15456 6736 15484
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 6917 15487 6975 15493
rect 6917 15453 6929 15487
rect 6963 15453 6975 15487
rect 6917 15447 6975 15453
rect 8665 15487 8723 15493
rect 8665 15453 8677 15487
rect 8711 15484 8723 15487
rect 9398 15484 9404 15496
rect 8711 15456 9404 15484
rect 8711 15453 8723 15456
rect 8665 15447 8723 15453
rect 2280 15388 2544 15416
rect 2280 15376 2286 15388
rect 5534 15376 5540 15428
rect 5592 15416 5598 15428
rect 6273 15419 6331 15425
rect 6273 15416 6285 15419
rect 5592 15388 6285 15416
rect 5592 15376 5598 15388
rect 6273 15385 6285 15388
rect 6319 15385 6331 15419
rect 6273 15379 6331 15385
rect 1670 15348 1676 15360
rect 1631 15320 1676 15348
rect 1670 15308 1676 15320
rect 1728 15308 1734 15360
rect 3050 15348 3056 15360
rect 3011 15320 3056 15348
rect 3050 15308 3056 15320
rect 3108 15308 3114 15360
rect 4798 15308 4804 15360
rect 4856 15348 4862 15360
rect 4982 15348 4988 15360
rect 4856 15320 4988 15348
rect 4856 15308 4862 15320
rect 4982 15308 4988 15320
rect 5040 15348 5046 15360
rect 5445 15351 5503 15357
rect 5445 15348 5457 15351
rect 5040 15320 5457 15348
rect 5040 15308 5046 15320
rect 5445 15317 5457 15320
rect 5491 15317 5503 15351
rect 5445 15311 5503 15317
rect 5813 15351 5871 15357
rect 5813 15317 5825 15351
rect 5859 15348 5871 15351
rect 5994 15348 6000 15360
rect 5859 15320 6000 15348
rect 5859 15317 5871 15320
rect 5813 15311 5871 15317
rect 5994 15308 6000 15320
rect 6052 15348 6058 15360
rect 6089 15351 6147 15357
rect 6089 15348 6101 15351
rect 6052 15320 6101 15348
rect 6052 15308 6058 15320
rect 6089 15317 6101 15320
rect 6135 15348 6147 15351
rect 6932 15348 6960 15447
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 9766 15484 9772 15496
rect 9727 15456 9772 15484
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 9858 15444 9864 15496
rect 9916 15484 9922 15496
rect 10318 15484 10324 15496
rect 9916 15456 10324 15484
rect 9916 15444 9922 15456
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 10686 15444 10692 15496
rect 10744 15484 10750 15496
rect 10781 15487 10839 15493
rect 10781 15484 10793 15487
rect 10744 15456 10793 15484
rect 10744 15444 10750 15456
rect 10781 15453 10793 15456
rect 10827 15453 10839 15487
rect 10781 15447 10839 15453
rect 12434 15444 12440 15496
rect 12492 15484 12498 15496
rect 13446 15484 13452 15496
rect 12492 15456 13452 15484
rect 12492 15444 12498 15456
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 13630 15484 13636 15496
rect 13591 15456 13636 15484
rect 13630 15444 13636 15456
rect 13688 15444 13694 15496
rect 15286 15484 15292 15496
rect 15247 15456 15292 15484
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15453 18659 15487
rect 18601 15447 18659 15453
rect 6135 15320 6960 15348
rect 7377 15351 7435 15357
rect 6135 15317 6147 15320
rect 6089 15311 6147 15317
rect 7377 15317 7389 15351
rect 7423 15348 7435 15351
rect 7558 15348 7564 15360
rect 7423 15320 7564 15348
rect 7423 15317 7435 15320
rect 7377 15311 7435 15317
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 7926 15308 7932 15360
rect 7984 15348 7990 15360
rect 9125 15351 9183 15357
rect 9125 15348 9137 15351
rect 7984 15320 9137 15348
rect 7984 15308 7990 15320
rect 9125 15317 9137 15320
rect 9171 15348 9183 15351
rect 9493 15351 9551 15357
rect 9493 15348 9505 15351
rect 9171 15320 9505 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 9493 15317 9505 15320
rect 9539 15348 9551 15351
rect 9674 15348 9680 15360
rect 9539 15320 9680 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 11422 15308 11428 15360
rect 11480 15348 11486 15360
rect 12158 15348 12164 15360
rect 11480 15320 12164 15348
rect 11480 15308 11486 15320
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 12529 15351 12587 15357
rect 12529 15317 12541 15351
rect 12575 15348 12587 15351
rect 13078 15348 13084 15360
rect 12575 15320 13084 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 13078 15308 13084 15320
rect 13136 15308 13142 15360
rect 15930 15308 15936 15360
rect 15988 15348 15994 15360
rect 16945 15351 17003 15357
rect 16945 15348 16957 15351
rect 15988 15320 16957 15348
rect 15988 15308 15994 15320
rect 16945 15317 16957 15320
rect 16991 15317 17003 15351
rect 18616 15348 18644 15447
rect 20254 15444 20260 15496
rect 20312 15484 20318 15496
rect 21453 15487 21511 15493
rect 21453 15484 21465 15487
rect 20312 15456 21465 15484
rect 20312 15444 20318 15456
rect 21453 15453 21465 15456
rect 21499 15453 21511 15487
rect 21453 15447 21511 15453
rect 23750 15444 23756 15496
rect 23808 15484 23814 15496
rect 24854 15484 24860 15496
rect 23808 15456 24860 15484
rect 23808 15444 23814 15456
rect 24854 15444 24860 15456
rect 24912 15444 24918 15496
rect 25314 15484 25320 15496
rect 25275 15456 25320 15484
rect 25314 15444 25320 15456
rect 25372 15444 25378 15496
rect 24118 15376 24124 15428
rect 24176 15416 24182 15428
rect 24673 15419 24731 15425
rect 24673 15416 24685 15419
rect 24176 15388 24685 15416
rect 24176 15376 24182 15388
rect 24673 15385 24685 15388
rect 24719 15385 24731 15419
rect 24673 15379 24731 15385
rect 18966 15348 18972 15360
rect 18616 15320 18972 15348
rect 16945 15311 17003 15317
rect 18966 15308 18972 15320
rect 19024 15348 19030 15360
rect 19242 15348 19248 15360
rect 19024 15320 19248 15348
rect 19024 15308 19030 15320
rect 19242 15308 19248 15320
rect 19300 15308 19306 15360
rect 20533 15351 20591 15357
rect 20533 15317 20545 15351
rect 20579 15348 20591 15351
rect 20714 15348 20720 15360
rect 20579 15320 20720 15348
rect 20579 15317 20591 15320
rect 20533 15311 20591 15317
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 20806 15308 20812 15360
rect 20864 15348 20870 15360
rect 20901 15351 20959 15357
rect 20901 15348 20913 15351
rect 20864 15320 20913 15348
rect 20864 15308 20870 15320
rect 20901 15317 20913 15320
rect 20947 15317 20959 15351
rect 20901 15311 20959 15317
rect 22738 15308 22744 15360
rect 22796 15348 22802 15360
rect 23658 15348 23664 15360
rect 22796 15320 23664 15348
rect 22796 15308 22802 15320
rect 23658 15308 23664 15320
rect 23716 15308 23722 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2314 15104 2320 15156
rect 2372 15144 2378 15156
rect 2501 15147 2559 15153
rect 2501 15144 2513 15147
rect 2372 15116 2513 15144
rect 2372 15104 2378 15116
rect 2501 15113 2513 15116
rect 2547 15144 2559 15147
rect 2685 15147 2743 15153
rect 2685 15144 2697 15147
rect 2547 15116 2697 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 2685 15113 2697 15116
rect 2731 15113 2743 15147
rect 5166 15144 5172 15156
rect 5127 15116 5172 15144
rect 2685 15107 2743 15113
rect 5166 15104 5172 15116
rect 5224 15104 5230 15156
rect 6270 15104 6276 15156
rect 6328 15144 6334 15156
rect 6549 15147 6607 15153
rect 6549 15144 6561 15147
rect 6328 15116 6561 15144
rect 6328 15104 6334 15116
rect 6549 15113 6561 15116
rect 6595 15144 6607 15147
rect 6825 15147 6883 15153
rect 6825 15144 6837 15147
rect 6595 15116 6837 15144
rect 6595 15113 6607 15116
rect 6549 15107 6607 15113
rect 6825 15113 6837 15116
rect 6871 15113 6883 15147
rect 7006 15144 7012 15156
rect 6967 15116 7012 15144
rect 6825 15107 6883 15113
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 8478 15144 8484 15156
rect 8439 15116 8484 15144
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 9125 15147 9183 15153
rect 9125 15113 9137 15147
rect 9171 15144 9183 15147
rect 9398 15144 9404 15156
rect 9171 15116 9404 15144
rect 9171 15113 9183 15116
rect 9125 15107 9183 15113
rect 9398 15104 9404 15116
rect 9456 15104 9462 15156
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11149 15147 11207 15153
rect 11149 15144 11161 15147
rect 11112 15116 11161 15144
rect 11112 15104 11118 15116
rect 11149 15113 11161 15116
rect 11195 15144 11207 15147
rect 11425 15147 11483 15153
rect 11425 15144 11437 15147
rect 11195 15116 11437 15144
rect 11195 15113 11207 15116
rect 11149 15107 11207 15113
rect 11425 15113 11437 15116
rect 11471 15113 11483 15147
rect 12158 15144 12164 15156
rect 12119 15116 12164 15144
rect 11425 15107 11483 15113
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 12342 15104 12348 15156
rect 12400 15144 12406 15156
rect 12437 15147 12495 15153
rect 12437 15144 12449 15147
rect 12400 15116 12449 15144
rect 12400 15104 12406 15116
rect 12437 15113 12449 15116
rect 12483 15113 12495 15147
rect 13538 15144 13544 15156
rect 13499 15116 13544 15144
rect 12437 15107 12495 15113
rect 13538 15104 13544 15116
rect 13596 15104 13602 15156
rect 13630 15104 13636 15156
rect 13688 15144 13694 15156
rect 13817 15147 13875 15153
rect 13817 15144 13829 15147
rect 13688 15116 13829 15144
rect 13688 15104 13694 15116
rect 13817 15113 13829 15116
rect 13863 15113 13875 15147
rect 17034 15144 17040 15156
rect 16995 15116 17040 15144
rect 13817 15107 13875 15113
rect 17034 15104 17040 15116
rect 17092 15104 17098 15156
rect 17862 15144 17868 15156
rect 17775 15116 17868 15144
rect 17862 15104 17868 15116
rect 17920 15144 17926 15156
rect 18874 15144 18880 15156
rect 17920 15116 18880 15144
rect 17920 15104 17926 15116
rect 18874 15104 18880 15116
rect 18932 15144 18938 15156
rect 19521 15147 19579 15153
rect 19521 15144 19533 15147
rect 18932 15116 19533 15144
rect 18932 15104 18938 15116
rect 19521 15113 19533 15116
rect 19567 15113 19579 15147
rect 20254 15144 20260 15156
rect 20215 15116 20260 15144
rect 19521 15107 19579 15113
rect 20254 15104 20260 15116
rect 20312 15104 20318 15156
rect 22002 15104 22008 15156
rect 22060 15144 22066 15156
rect 22370 15144 22376 15156
rect 22060 15116 22376 15144
rect 22060 15104 22066 15116
rect 22370 15104 22376 15116
rect 22428 15104 22434 15156
rect 22646 15144 22652 15156
rect 22607 15116 22652 15144
rect 22646 15104 22652 15116
rect 22704 15104 22710 15156
rect 23661 15147 23719 15153
rect 23661 15113 23673 15147
rect 23707 15144 23719 15147
rect 23934 15144 23940 15156
rect 23707 15116 23940 15144
rect 23707 15113 23719 15116
rect 23661 15107 23719 15113
rect 23934 15104 23940 15116
rect 23992 15104 23998 15156
rect 24762 15144 24768 15156
rect 24723 15116 24768 15144
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 24949 15147 25007 15153
rect 24949 15113 24961 15147
rect 24995 15144 25007 15147
rect 25041 15147 25099 15153
rect 25041 15144 25053 15147
rect 24995 15116 25053 15144
rect 24995 15113 25007 15116
rect 24949 15107 25007 15113
rect 25041 15113 25053 15116
rect 25087 15144 25099 15147
rect 25314 15144 25320 15156
rect 25087 15116 25320 15144
rect 25087 15113 25099 15116
rect 25041 15107 25099 15113
rect 25314 15104 25320 15116
rect 25372 15104 25378 15156
rect 2225 15079 2283 15085
rect 2225 15045 2237 15079
rect 2271 15076 2283 15079
rect 2406 15076 2412 15088
rect 2271 15048 2412 15076
rect 2271 15045 2283 15048
rect 2225 15039 2283 15045
rect 2406 15036 2412 15048
rect 2464 15036 2470 15088
rect 8113 15079 8171 15085
rect 8113 15045 8125 15079
rect 8159 15076 8171 15079
rect 8386 15076 8392 15088
rect 8159 15048 8392 15076
rect 8159 15045 8171 15048
rect 8113 15039 8171 15045
rect 8386 15036 8392 15048
rect 8444 15036 8450 15088
rect 12176 15076 12204 15104
rect 12176 15048 13124 15076
rect 1670 15008 1676 15020
rect 1412 14980 1676 15008
rect 1412 14949 1440 14980
rect 1670 14968 1676 14980
rect 1728 14968 1734 15020
rect 2774 14968 2780 15020
rect 2832 15008 2838 15020
rect 5077 15011 5135 15017
rect 2832 14980 2877 15008
rect 2832 14968 2838 14980
rect 5077 14977 5089 15011
rect 5123 15008 5135 15011
rect 5721 15011 5779 15017
rect 5721 15008 5733 15011
rect 5123 14980 5733 15008
rect 5123 14977 5135 14980
rect 5077 14971 5135 14977
rect 5721 14977 5733 14980
rect 5767 15008 5779 15011
rect 6546 15008 6552 15020
rect 5767 14980 6552 15008
rect 5767 14977 5779 14980
rect 5721 14971 5779 14977
rect 6546 14968 6552 14980
rect 6604 14968 6610 15020
rect 7650 15008 7656 15020
rect 7611 14980 7656 15008
rect 7650 14968 7656 14980
rect 7708 14968 7714 15020
rect 8570 15008 8576 15020
rect 8531 14980 8576 15008
rect 8570 14968 8576 14980
rect 8628 14968 8634 15020
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 15008 11943 15011
rect 12434 15008 12440 15020
rect 11931 14980 12440 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 12434 14968 12440 14980
rect 12492 14968 12498 15020
rect 13096 15017 13124 15048
rect 13081 15011 13139 15017
rect 13081 14977 13093 15011
rect 13127 15008 13139 15011
rect 13648 15008 13676 15104
rect 22186 15036 22192 15088
rect 22244 15076 22250 15088
rect 22554 15076 22560 15088
rect 22244 15048 22560 15076
rect 22244 15036 22250 15048
rect 22554 15036 22560 15048
rect 22612 15036 22618 15088
rect 24670 15036 24676 15088
rect 24728 15076 24734 15088
rect 25409 15079 25467 15085
rect 25409 15076 25421 15079
rect 24728 15048 25421 15076
rect 24728 15036 24734 15048
rect 25409 15045 25421 15048
rect 25455 15045 25467 15079
rect 25409 15039 25467 15045
rect 13127 14980 13676 15008
rect 13127 14977 13139 14980
rect 13081 14971 13139 14977
rect 17218 14968 17224 15020
rect 17276 15008 17282 15020
rect 19889 15011 19947 15017
rect 17276 14980 18276 15008
rect 17276 14968 17282 14980
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14909 1455 14943
rect 1397 14903 1455 14909
rect 1670 14872 1676 14884
rect 1631 14844 1676 14872
rect 1670 14832 1676 14844
rect 1728 14832 1734 14884
rect 2792 14872 2820 14968
rect 3050 14949 3056 14952
rect 3044 14940 3056 14949
rect 3011 14912 3056 14940
rect 3044 14903 3056 14912
rect 3050 14900 3056 14903
rect 3108 14900 3114 14952
rect 5534 14940 5540 14952
rect 5495 14912 5540 14940
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 6270 14940 6276 14952
rect 6183 14912 6276 14940
rect 6270 14900 6276 14912
rect 6328 14940 6334 14952
rect 7668 14940 7696 14968
rect 9766 14940 9772 14952
rect 6328 14912 7696 14940
rect 9679 14912 9772 14940
rect 6328 14900 6334 14912
rect 9766 14900 9772 14912
rect 9824 14940 9830 14952
rect 12897 14943 12955 14949
rect 9824 14912 10732 14940
rect 9824 14900 9830 14912
rect 10704 14884 10732 14912
rect 12897 14909 12909 14943
rect 12943 14940 12955 14943
rect 13722 14940 13728 14952
rect 12943 14912 13728 14940
rect 12943 14909 12955 14912
rect 12897 14903 12955 14909
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 14366 14900 14372 14952
rect 14424 14940 14430 14952
rect 14645 14943 14703 14949
rect 14645 14940 14657 14943
rect 14424 14912 14657 14940
rect 14424 14900 14430 14912
rect 14645 14909 14657 14912
rect 14691 14940 14703 14943
rect 15286 14940 15292 14952
rect 14691 14912 15292 14940
rect 14691 14909 14703 14912
rect 14645 14903 14703 14909
rect 15286 14900 15292 14912
rect 15344 14900 15350 14952
rect 16853 14943 16911 14949
rect 16853 14940 16865 14943
rect 16684 14912 16865 14940
rect 2958 14872 2964 14884
rect 2792 14844 2964 14872
rect 2958 14832 2964 14844
rect 3016 14832 3022 14884
rect 6825 14875 6883 14881
rect 6825 14841 6837 14875
rect 6871 14872 6883 14875
rect 7374 14872 7380 14884
rect 6871 14844 7380 14872
rect 6871 14841 6883 14844
rect 6825 14835 6883 14841
rect 7374 14832 7380 14844
rect 7432 14832 7438 14884
rect 9677 14875 9735 14881
rect 9677 14841 9689 14875
rect 9723 14872 9735 14875
rect 10036 14875 10094 14881
rect 10036 14872 10048 14875
rect 9723 14844 10048 14872
rect 9723 14841 9735 14844
rect 9677 14835 9735 14841
rect 10036 14841 10048 14844
rect 10082 14872 10094 14875
rect 10134 14872 10140 14884
rect 10082 14844 10140 14872
rect 10082 14841 10094 14844
rect 10036 14835 10094 14841
rect 10134 14832 10140 14844
rect 10192 14832 10198 14884
rect 10686 14832 10692 14884
rect 10744 14832 10750 14884
rect 14553 14875 14611 14881
rect 14553 14841 14565 14875
rect 14599 14872 14611 14875
rect 14734 14872 14740 14884
rect 14599 14844 14740 14872
rect 14599 14841 14611 14844
rect 14553 14835 14611 14841
rect 14734 14832 14740 14844
rect 14792 14872 14798 14884
rect 14890 14875 14948 14881
rect 14890 14872 14902 14875
rect 14792 14844 14902 14872
rect 14792 14832 14798 14844
rect 14890 14841 14902 14844
rect 14936 14841 14948 14875
rect 14890 14835 14948 14841
rect 16684 14816 16712 14912
rect 16853 14909 16865 14912
rect 16899 14909 16911 14943
rect 16853 14903 16911 14909
rect 17770 14900 17776 14952
rect 17828 14940 17834 14952
rect 18046 14940 18052 14952
rect 17828 14912 18052 14940
rect 17828 14900 17834 14912
rect 18046 14900 18052 14912
rect 18104 14940 18110 14952
rect 18141 14943 18199 14949
rect 18141 14940 18153 14943
rect 18104 14912 18153 14940
rect 18104 14900 18110 14912
rect 18141 14909 18153 14912
rect 18187 14909 18199 14943
rect 18248 14940 18276 14980
rect 19889 14977 19901 15011
rect 19935 15008 19947 15011
rect 20806 15008 20812 15020
rect 19935 14980 20812 15008
rect 19935 14977 19947 14980
rect 19889 14971 19947 14977
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 20898 14968 20904 15020
rect 20956 15008 20962 15020
rect 23109 15011 23167 15017
rect 20956 14980 21001 15008
rect 20956 14968 20962 14980
rect 23109 14977 23121 15011
rect 23155 15008 23167 15011
rect 24213 15011 24271 15017
rect 24213 15008 24225 15011
rect 23155 14980 24225 15008
rect 23155 14977 23167 14980
rect 23109 14971 23167 14977
rect 24213 14977 24225 14980
rect 24259 15008 24271 15011
rect 24949 15011 25007 15017
rect 24949 15008 24961 15011
rect 24259 14980 24961 15008
rect 24259 14977 24271 14980
rect 24213 14971 24271 14977
rect 24949 14977 24961 14980
rect 24995 14977 25007 15011
rect 24949 14971 25007 14977
rect 20162 14940 20168 14952
rect 18248 14912 20168 14940
rect 18141 14903 18199 14909
rect 20162 14900 20168 14912
rect 20220 14940 20226 14952
rect 20530 14940 20536 14952
rect 20220 14912 20536 14940
rect 20220 14900 20226 14912
rect 20530 14900 20536 14912
rect 20588 14940 20594 14952
rect 21361 14943 21419 14949
rect 21361 14940 21373 14943
rect 20588 14912 21373 14940
rect 20588 14900 20594 14912
rect 21361 14909 21373 14912
rect 21407 14909 21419 14943
rect 21910 14940 21916 14952
rect 21871 14912 21916 14940
rect 21361 14903 21419 14909
rect 21910 14900 21916 14912
rect 21968 14900 21974 14952
rect 23658 14900 23664 14952
rect 23716 14940 23722 14952
rect 24029 14943 24087 14949
rect 24029 14940 24041 14943
rect 23716 14912 24041 14940
rect 23716 14900 23722 14912
rect 24029 14909 24041 14912
rect 24075 14909 24087 14943
rect 25225 14943 25283 14949
rect 25225 14940 25237 14943
rect 24029 14903 24087 14909
rect 24136 14912 25237 14940
rect 17497 14875 17555 14881
rect 17497 14841 17509 14875
rect 17543 14872 17555 14875
rect 18408 14875 18466 14881
rect 18408 14872 18420 14875
rect 17543 14844 18420 14872
rect 17543 14841 17555 14844
rect 17497 14835 17555 14841
rect 18408 14841 18420 14844
rect 18454 14872 18466 14875
rect 19242 14872 19248 14884
rect 18454 14844 19248 14872
rect 18454 14841 18466 14844
rect 18408 14835 18466 14841
rect 19242 14832 19248 14844
rect 19300 14832 19306 14884
rect 19978 14832 19984 14884
rect 20036 14872 20042 14884
rect 20717 14875 20775 14881
rect 20717 14872 20729 14875
rect 20036 14844 20729 14872
rect 20036 14832 20042 14844
rect 20717 14841 20729 14844
rect 20763 14841 20775 14875
rect 20717 14835 20775 14841
rect 20806 14832 20812 14884
rect 20864 14872 20870 14884
rect 21450 14872 21456 14884
rect 20864 14844 21456 14872
rect 20864 14832 20870 14844
rect 21450 14832 21456 14844
rect 21508 14872 21514 14884
rect 21729 14875 21787 14881
rect 21729 14872 21741 14875
rect 21508 14844 21741 14872
rect 21508 14832 21514 14844
rect 21729 14841 21741 14844
rect 21775 14841 21787 14875
rect 22186 14872 22192 14884
rect 22147 14844 22192 14872
rect 21729 14835 21787 14841
rect 22186 14832 22192 14844
rect 22244 14832 22250 14884
rect 23474 14872 23480 14884
rect 23435 14844 23480 14872
rect 23474 14832 23480 14844
rect 23532 14872 23538 14884
rect 24136 14881 24164 14912
rect 25225 14909 25237 14912
rect 25271 14940 25283 14943
rect 25777 14943 25835 14949
rect 25777 14940 25789 14943
rect 25271 14912 25789 14940
rect 25271 14909 25283 14912
rect 25225 14903 25283 14909
rect 25777 14909 25789 14912
rect 25823 14909 25835 14943
rect 25777 14903 25835 14909
rect 24121 14875 24179 14881
rect 24121 14872 24133 14875
rect 23532 14844 24133 14872
rect 23532 14832 23538 14844
rect 24121 14841 24133 14844
rect 24167 14841 24179 14875
rect 24121 14835 24179 14841
rect 2685 14807 2743 14813
rect 2685 14773 2697 14807
rect 2731 14804 2743 14807
rect 2774 14804 2780 14816
rect 2731 14776 2780 14804
rect 2731 14773 2743 14776
rect 2685 14767 2743 14773
rect 2774 14764 2780 14776
rect 2832 14764 2838 14816
rect 4154 14804 4160 14816
rect 4115 14776 4160 14804
rect 4154 14764 4160 14776
rect 4212 14804 4218 14816
rect 4433 14807 4491 14813
rect 4433 14804 4445 14807
rect 4212 14776 4445 14804
rect 4212 14764 4218 14776
rect 4433 14773 4445 14776
rect 4479 14773 4491 14807
rect 5626 14804 5632 14816
rect 5587 14776 5632 14804
rect 4433 14767 4491 14773
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 7469 14807 7527 14813
rect 7469 14773 7481 14807
rect 7515 14804 7527 14807
rect 7558 14804 7564 14816
rect 7515 14776 7564 14804
rect 7515 14773 7527 14776
rect 7469 14767 7527 14773
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 12802 14804 12808 14816
rect 12763 14776 12808 14804
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 15838 14764 15844 14816
rect 15896 14804 15902 14816
rect 16025 14807 16083 14813
rect 16025 14804 16037 14807
rect 15896 14776 16037 14804
rect 15896 14764 15902 14776
rect 16025 14773 16037 14776
rect 16071 14773 16083 14807
rect 16025 14767 16083 14773
rect 16114 14764 16120 14816
rect 16172 14804 16178 14816
rect 16301 14807 16359 14813
rect 16301 14804 16313 14807
rect 16172 14776 16313 14804
rect 16172 14764 16178 14776
rect 16301 14773 16313 14776
rect 16347 14773 16359 14807
rect 16666 14804 16672 14816
rect 16627 14776 16672 14804
rect 16301 14767 16359 14773
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 20346 14804 20352 14816
rect 20307 14776 20352 14804
rect 20346 14764 20352 14776
rect 20404 14764 20410 14816
rect 21818 14764 21824 14816
rect 21876 14804 21882 14816
rect 22646 14804 22652 14816
rect 21876 14776 22652 14804
rect 21876 14764 21882 14776
rect 22646 14764 22652 14776
rect 22704 14764 22710 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1949 14603 2007 14609
rect 1949 14569 1961 14603
rect 1995 14600 2007 14603
rect 2222 14600 2228 14612
rect 1995 14572 2228 14600
rect 1995 14569 2007 14572
rect 1949 14563 2007 14569
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 2409 14603 2467 14609
rect 2409 14569 2421 14603
rect 2455 14600 2467 14603
rect 2498 14600 2504 14612
rect 2455 14572 2504 14600
rect 2455 14569 2467 14572
rect 2409 14563 2467 14569
rect 2498 14560 2504 14572
rect 2556 14560 2562 14612
rect 2869 14603 2927 14609
rect 2869 14569 2881 14603
rect 2915 14600 2927 14603
rect 3237 14603 3295 14609
rect 3237 14600 3249 14603
rect 2915 14572 3249 14600
rect 2915 14569 2927 14572
rect 2869 14563 2927 14569
rect 3237 14569 3249 14572
rect 3283 14600 3295 14603
rect 3602 14600 3608 14612
rect 3283 14572 3608 14600
rect 3283 14569 3295 14572
rect 3237 14563 3295 14569
rect 3602 14560 3608 14572
rect 3660 14560 3666 14612
rect 3878 14600 3884 14612
rect 3839 14572 3884 14600
rect 3878 14560 3884 14572
rect 3936 14560 3942 14612
rect 4249 14603 4307 14609
rect 4249 14569 4261 14603
rect 4295 14600 4307 14603
rect 5721 14603 5779 14609
rect 5721 14600 5733 14603
rect 4295 14572 5733 14600
rect 4295 14569 4307 14572
rect 4249 14563 4307 14569
rect 5721 14569 5733 14572
rect 5767 14600 5779 14603
rect 6730 14600 6736 14612
rect 5767 14572 6736 14600
rect 5767 14569 5779 14572
rect 5721 14563 5779 14569
rect 6730 14560 6736 14572
rect 6788 14560 6794 14612
rect 8018 14600 8024 14612
rect 7979 14572 8024 14600
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 8389 14603 8447 14609
rect 8389 14569 8401 14603
rect 8435 14600 8447 14603
rect 8478 14600 8484 14612
rect 8435 14572 8484 14600
rect 8435 14569 8447 14572
rect 8389 14563 8447 14569
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 8754 14560 8760 14612
rect 8812 14600 8818 14612
rect 9033 14603 9091 14609
rect 9033 14600 9045 14603
rect 8812 14572 9045 14600
rect 8812 14560 8818 14572
rect 9033 14569 9045 14572
rect 9079 14569 9091 14603
rect 9033 14563 9091 14569
rect 9493 14603 9551 14609
rect 9493 14569 9505 14603
rect 9539 14600 9551 14603
rect 9766 14600 9772 14612
rect 9539 14572 9772 14600
rect 9539 14569 9551 14572
rect 9493 14563 9551 14569
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 10778 14600 10784 14612
rect 10643 14572 10784 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 4617 14535 4675 14541
rect 4617 14501 4629 14535
rect 4663 14532 4675 14535
rect 4890 14532 4896 14544
rect 4663 14504 4896 14532
rect 4663 14501 4675 14504
rect 4617 14495 4675 14501
rect 4890 14492 4896 14504
rect 4948 14492 4954 14544
rect 5350 14532 5356 14544
rect 5311 14504 5356 14532
rect 5350 14492 5356 14504
rect 5408 14492 5414 14544
rect 6080 14535 6138 14541
rect 6080 14532 6092 14535
rect 5736 14504 6092 14532
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 4706 14464 4712 14476
rect 2832 14436 4712 14464
rect 2832 14424 2838 14436
rect 4706 14424 4712 14436
rect 4764 14464 4770 14476
rect 5442 14464 5448 14476
rect 4764 14436 5448 14464
rect 4764 14424 4770 14436
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14396 1455 14399
rect 2038 14396 2044 14408
rect 1443 14368 2044 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 2038 14356 2044 14368
rect 2096 14356 2102 14408
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14396 2375 14399
rect 3053 14399 3111 14405
rect 3053 14396 3065 14399
rect 2363 14368 3065 14396
rect 2363 14365 2375 14368
rect 2317 14359 2375 14365
rect 3053 14365 3065 14368
rect 3099 14396 3111 14399
rect 4798 14396 4804 14408
rect 3099 14368 4804 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 4798 14356 4804 14368
rect 4856 14356 4862 14408
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14396 4951 14399
rect 5736 14396 5764 14504
rect 6080 14501 6092 14504
rect 6126 14532 6138 14535
rect 6270 14532 6276 14544
rect 6126 14504 6276 14532
rect 6126 14501 6138 14504
rect 6080 14495 6138 14501
rect 6270 14492 6276 14504
rect 6328 14492 6334 14544
rect 10612 14532 10640 14563
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 10962 14600 10968 14612
rect 10923 14572 10968 14600
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 12713 14603 12771 14609
rect 12713 14600 12725 14603
rect 12676 14572 12725 14600
rect 12676 14560 12682 14572
rect 12713 14569 12725 14572
rect 12759 14569 12771 14603
rect 12713 14563 12771 14569
rect 9784 14504 10640 14532
rect 11324 14535 11382 14541
rect 5813 14467 5871 14473
rect 5813 14433 5825 14467
rect 5859 14464 5871 14467
rect 6822 14464 6828 14476
rect 5859 14436 6828 14464
rect 5859 14433 5871 14436
rect 5813 14427 5871 14433
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 8386 14424 8392 14476
rect 8444 14464 8450 14476
rect 9784 14473 9812 14504
rect 11324 14501 11336 14535
rect 11370 14532 11382 14535
rect 11974 14532 11980 14544
rect 11370 14504 11980 14532
rect 11370 14501 11382 14504
rect 11324 14495 11382 14501
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 12728 14532 12756 14563
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 13265 14603 13323 14609
rect 13265 14600 13277 14603
rect 12860 14572 13277 14600
rect 12860 14560 12866 14572
rect 13265 14569 13277 14572
rect 13311 14569 13323 14603
rect 13265 14563 13323 14569
rect 15105 14603 15163 14609
rect 15105 14569 15117 14603
rect 15151 14600 15163 14603
rect 16209 14603 16267 14609
rect 16209 14600 16221 14603
rect 15151 14572 16221 14600
rect 15151 14569 15163 14572
rect 15105 14563 15163 14569
rect 16209 14569 16221 14572
rect 16255 14600 16267 14603
rect 16390 14600 16396 14612
rect 16255 14572 16396 14600
rect 16255 14569 16267 14572
rect 16209 14563 16267 14569
rect 16390 14560 16396 14572
rect 16448 14560 16454 14612
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 16669 14603 16727 14609
rect 16669 14600 16681 14603
rect 16632 14572 16681 14600
rect 16632 14560 16638 14572
rect 16669 14569 16681 14572
rect 16715 14569 16727 14603
rect 16669 14563 16727 14569
rect 17310 14560 17316 14612
rect 17368 14600 17374 14612
rect 17497 14603 17555 14609
rect 17497 14600 17509 14603
rect 17368 14572 17509 14600
rect 17368 14560 17374 14572
rect 17497 14569 17509 14572
rect 17543 14569 17555 14603
rect 19242 14600 19248 14612
rect 19155 14572 19248 14600
rect 17497 14563 17555 14569
rect 19242 14560 19248 14572
rect 19300 14600 19306 14612
rect 20441 14603 20499 14609
rect 20441 14600 20453 14603
rect 19300 14572 20453 14600
rect 19300 14560 19306 14572
rect 20441 14569 20453 14572
rect 20487 14600 20499 14603
rect 20898 14600 20904 14612
rect 20487 14572 20904 14600
rect 20487 14569 20499 14572
rect 20441 14563 20499 14569
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 20990 14560 20996 14612
rect 21048 14600 21054 14612
rect 21085 14603 21143 14609
rect 21085 14600 21097 14603
rect 21048 14572 21097 14600
rect 21048 14560 21054 14572
rect 21085 14569 21097 14572
rect 21131 14569 21143 14603
rect 21542 14600 21548 14612
rect 21503 14572 21548 14600
rect 21085 14563 21143 14569
rect 21542 14560 21548 14572
rect 21600 14560 21606 14612
rect 22002 14600 22008 14612
rect 21963 14572 22008 14600
rect 22002 14560 22008 14572
rect 22060 14560 22066 14612
rect 22373 14603 22431 14609
rect 22373 14569 22385 14603
rect 22419 14600 22431 14603
rect 22462 14600 22468 14612
rect 22419 14572 22468 14600
rect 22419 14569 22431 14572
rect 22373 14563 22431 14569
rect 22462 14560 22468 14572
rect 22520 14600 22526 14612
rect 22649 14603 22707 14609
rect 22649 14600 22661 14603
rect 22520 14572 22661 14600
rect 22520 14560 22526 14572
rect 22649 14569 22661 14572
rect 22695 14569 22707 14603
rect 22649 14563 22707 14569
rect 22922 14560 22928 14612
rect 22980 14600 22986 14612
rect 23106 14600 23112 14612
rect 22980 14572 23112 14600
rect 22980 14560 22986 14572
rect 23106 14560 23112 14572
rect 23164 14560 23170 14612
rect 23290 14560 23296 14612
rect 23348 14600 23354 14612
rect 24029 14603 24087 14609
rect 24029 14600 24041 14603
rect 23348 14572 24041 14600
rect 23348 14560 23354 14572
rect 24029 14569 24041 14572
rect 24075 14569 24087 14603
rect 24029 14563 24087 14569
rect 25041 14603 25099 14609
rect 25041 14569 25053 14603
rect 25087 14600 25099 14603
rect 25130 14600 25136 14612
rect 25087 14572 25136 14600
rect 25087 14569 25099 14572
rect 25041 14563 25099 14569
rect 25130 14560 25136 14572
rect 25188 14560 25194 14612
rect 13633 14535 13691 14541
rect 13633 14532 13645 14535
rect 12728 14504 13645 14532
rect 13633 14501 13645 14504
rect 13679 14501 13691 14535
rect 13633 14495 13691 14501
rect 13722 14492 13728 14544
rect 13780 14532 13786 14544
rect 15378 14532 15384 14544
rect 13780 14504 15384 14532
rect 13780 14492 13786 14504
rect 15378 14492 15384 14504
rect 15436 14492 15442 14544
rect 16482 14492 16488 14544
rect 16540 14532 16546 14544
rect 16761 14535 16819 14541
rect 16761 14532 16773 14535
rect 16540 14504 16773 14532
rect 16540 14492 16546 14504
rect 16761 14501 16773 14504
rect 16807 14501 16819 14535
rect 16761 14495 16819 14501
rect 17586 14492 17592 14544
rect 17644 14532 17650 14544
rect 18132 14535 18190 14541
rect 18132 14532 18144 14535
rect 17644 14504 18144 14532
rect 17644 14492 17650 14504
rect 18132 14501 18144 14504
rect 18178 14532 18190 14535
rect 19610 14532 19616 14544
rect 18178 14504 19616 14532
rect 18178 14501 18190 14504
rect 18132 14495 18190 14501
rect 19610 14492 19616 14504
rect 19668 14532 19674 14544
rect 19705 14535 19763 14541
rect 19705 14532 19717 14535
rect 19668 14504 19717 14532
rect 19668 14492 19674 14504
rect 19705 14501 19717 14504
rect 19751 14532 19763 14535
rect 20254 14532 20260 14544
rect 19751 14504 20260 14532
rect 19751 14501 19763 14504
rect 19705 14495 19763 14501
rect 20254 14492 20260 14504
rect 20312 14492 20318 14544
rect 8481 14467 8539 14473
rect 8481 14464 8493 14467
rect 8444 14436 8493 14464
rect 8444 14424 8450 14436
rect 8481 14433 8493 14436
rect 8527 14433 8539 14467
rect 8481 14427 8539 14433
rect 9769 14467 9827 14473
rect 9769 14433 9781 14467
rect 9815 14433 9827 14467
rect 10042 14464 10048 14476
rect 10003 14436 10048 14464
rect 9769 14427 9827 14433
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 10686 14424 10692 14476
rect 10744 14464 10750 14476
rect 11057 14467 11115 14473
rect 11057 14464 11069 14467
rect 10744 14436 11069 14464
rect 10744 14424 10750 14436
rect 11057 14433 11069 14436
rect 11103 14433 11115 14467
rect 11057 14427 11115 14433
rect 13538 14424 13544 14476
rect 13596 14464 13602 14476
rect 13596 14436 13860 14464
rect 13596 14424 13602 14436
rect 7466 14396 7472 14408
rect 4939 14368 5764 14396
rect 7427 14368 7472 14396
rect 4939 14365 4951 14368
rect 4893 14359 4951 14365
rect 1946 14288 1952 14340
rect 2004 14328 2010 14340
rect 3421 14331 3479 14337
rect 3421 14328 3433 14331
rect 2004 14300 3433 14328
rect 2004 14288 2010 14300
rect 3421 14297 3433 14300
rect 3467 14297 3479 14331
rect 3421 14291 3479 14297
rect 3878 14288 3884 14340
rect 3936 14328 3942 14340
rect 4908 14328 4936 14359
rect 7466 14356 7472 14368
rect 7524 14356 7530 14408
rect 8665 14399 8723 14405
rect 8665 14365 8677 14399
rect 8711 14396 8723 14399
rect 10134 14396 10140 14408
rect 8711 14368 10140 14396
rect 8711 14365 8723 14368
rect 8665 14359 8723 14365
rect 3936 14300 4936 14328
rect 7929 14331 7987 14337
rect 3936 14288 3942 14300
rect 7929 14297 7941 14331
rect 7975 14328 7987 14331
rect 8680 14328 8708 14359
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 12802 14356 12808 14408
rect 12860 14396 12866 14408
rect 13173 14399 13231 14405
rect 13173 14396 13185 14399
rect 12860 14368 13185 14396
rect 12860 14356 12866 14368
rect 13173 14365 13185 14368
rect 13219 14396 13231 14399
rect 13722 14396 13728 14408
rect 13219 14368 13728 14396
rect 13219 14365 13231 14368
rect 13173 14359 13231 14365
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 13832 14405 13860 14436
rect 20530 14424 20536 14476
rect 20588 14464 20594 14476
rect 20717 14467 20775 14473
rect 20717 14464 20729 14467
rect 20588 14436 20729 14464
rect 20588 14424 20594 14436
rect 20717 14433 20729 14436
rect 20763 14433 20775 14467
rect 20717 14427 20775 14433
rect 20901 14467 20959 14473
rect 20901 14433 20913 14467
rect 20947 14464 20959 14467
rect 20990 14464 20996 14476
rect 20947 14436 20996 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 20990 14424 20996 14436
rect 21048 14464 21054 14476
rect 21358 14464 21364 14476
rect 21048 14436 21364 14464
rect 21048 14424 21054 14436
rect 21358 14424 21364 14436
rect 21416 14424 21422 14476
rect 22370 14424 22376 14476
rect 22428 14464 22434 14476
rect 23017 14467 23075 14473
rect 23017 14464 23029 14467
rect 22428 14436 23029 14464
rect 22428 14424 22434 14436
rect 23017 14433 23029 14436
rect 23063 14464 23075 14467
rect 23382 14464 23388 14476
rect 23063 14436 23388 14464
rect 23063 14433 23075 14436
rect 23017 14427 23075 14433
rect 23382 14424 23388 14436
rect 23440 14424 23446 14476
rect 24210 14464 24216 14476
rect 24171 14436 24216 14464
rect 24210 14424 24216 14436
rect 24268 14424 24274 14476
rect 13817 14399 13875 14405
rect 13817 14365 13829 14399
rect 13863 14365 13875 14399
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 13817 14359 13875 14365
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 16758 14356 16764 14408
rect 16816 14396 16822 14408
rect 16945 14399 17003 14405
rect 16945 14396 16957 14399
rect 16816 14368 16957 14396
rect 16816 14356 16822 14368
rect 16945 14365 16957 14368
rect 16991 14396 17003 14399
rect 17586 14396 17592 14408
rect 16991 14368 17592 14396
rect 16991 14365 17003 14368
rect 16945 14359 17003 14365
rect 17586 14356 17592 14368
rect 17644 14356 17650 14408
rect 17770 14356 17776 14408
rect 17828 14396 17834 14408
rect 17865 14399 17923 14405
rect 17865 14396 17877 14399
rect 17828 14368 17877 14396
rect 17828 14356 17834 14368
rect 17865 14365 17877 14368
rect 17911 14365 17923 14399
rect 19978 14396 19984 14408
rect 19939 14368 19984 14396
rect 17865 14359 17923 14365
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 23106 14396 23112 14408
rect 20220 14368 23112 14396
rect 20220 14356 20226 14368
rect 23106 14356 23112 14368
rect 23164 14356 23170 14408
rect 23201 14399 23259 14405
rect 23201 14365 23213 14399
rect 23247 14365 23259 14399
rect 23201 14359 23259 14365
rect 24489 14399 24547 14405
rect 24489 14365 24501 14399
rect 24535 14396 24547 14399
rect 24670 14396 24676 14408
rect 24535 14368 24676 14396
rect 24535 14365 24547 14368
rect 24489 14359 24547 14365
rect 16298 14328 16304 14340
rect 7975 14300 8708 14328
rect 16259 14300 16304 14328
rect 7975 14297 7987 14300
rect 7929 14291 7987 14297
rect 16298 14288 16304 14300
rect 16356 14288 16362 14340
rect 20898 14288 20904 14340
rect 20956 14328 20962 14340
rect 21634 14328 21640 14340
rect 20956 14300 21640 14328
rect 20956 14288 20962 14300
rect 21634 14288 21640 14300
rect 21692 14288 21698 14340
rect 21818 14288 21824 14340
rect 21876 14328 21882 14340
rect 23216 14328 23244 14359
rect 24670 14356 24676 14368
rect 24728 14356 24734 14408
rect 21876 14300 23244 14328
rect 21876 14288 21882 14300
rect 3234 14260 3240 14272
rect 3195 14232 3240 14260
rect 3234 14220 3240 14232
rect 3292 14220 3298 14272
rect 5994 14220 6000 14272
rect 6052 14260 6058 14272
rect 7193 14263 7251 14269
rect 7193 14260 7205 14263
rect 6052 14232 7205 14260
rect 6052 14220 6058 14232
rect 7193 14229 7205 14232
rect 7239 14229 7251 14263
rect 7193 14223 7251 14229
rect 9674 14220 9680 14272
rect 9732 14260 9738 14272
rect 11790 14260 11796 14272
rect 9732 14232 11796 14260
rect 9732 14220 9738 14232
rect 11790 14220 11796 14232
rect 11848 14220 11854 14272
rect 12158 14220 12164 14272
rect 12216 14260 12222 14272
rect 12437 14263 12495 14269
rect 12437 14260 12449 14263
rect 12216 14232 12449 14260
rect 12216 14220 12222 14232
rect 12437 14229 12449 14232
rect 12483 14229 12495 14263
rect 12437 14223 12495 14229
rect 13998 14220 14004 14272
rect 14056 14260 14062 14272
rect 14277 14263 14335 14269
rect 14277 14260 14289 14263
rect 14056 14232 14289 14260
rect 14056 14220 14062 14232
rect 14277 14229 14289 14232
rect 14323 14229 14335 14263
rect 14642 14260 14648 14272
rect 14603 14232 14648 14260
rect 14277 14223 14335 14229
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 15838 14260 15844 14272
rect 15799 14232 15844 14260
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 19518 14260 19524 14272
rect 19392 14232 19524 14260
rect 19392 14220 19398 14232
rect 19518 14220 19524 14232
rect 19576 14260 19582 14272
rect 20533 14263 20591 14269
rect 20533 14260 20545 14263
rect 19576 14232 20545 14260
rect 19576 14220 19582 14232
rect 20533 14229 20545 14232
rect 20579 14229 20591 14263
rect 20533 14223 20591 14229
rect 22278 14220 22284 14272
rect 22336 14260 22342 14272
rect 22554 14260 22560 14272
rect 22336 14232 22560 14260
rect 22336 14220 22342 14232
rect 22554 14220 22560 14232
rect 22612 14220 22618 14272
rect 23658 14260 23664 14272
rect 23619 14232 23664 14260
rect 23658 14220 23664 14232
rect 23716 14220 23722 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2501 14059 2559 14065
rect 2501 14025 2513 14059
rect 2547 14056 2559 14059
rect 2547 14028 2820 14056
rect 2547 14025 2559 14028
rect 2501 14019 2559 14025
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 1854 13920 1860 13932
rect 1719 13892 1860 13920
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 1946 13852 1952 13864
rect 1443 13824 1952 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 2792 13716 2820 14028
rect 3050 14016 3056 14068
rect 3108 14056 3114 14068
rect 4249 14059 4307 14065
rect 4249 14056 4261 14059
rect 3108 14028 4261 14056
rect 3108 14016 3114 14028
rect 4249 14025 4261 14028
rect 4295 14025 4307 14059
rect 4249 14019 4307 14025
rect 4617 14059 4675 14065
rect 4617 14025 4629 14059
rect 4663 14056 4675 14059
rect 4706 14056 4712 14068
rect 4663 14028 4712 14056
rect 4663 14025 4675 14028
rect 4617 14019 4675 14025
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 4890 14056 4896 14068
rect 4851 14028 4896 14056
rect 4890 14016 4896 14028
rect 4948 14016 4954 14068
rect 5166 14056 5172 14068
rect 5127 14028 5172 14056
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 6270 14056 6276 14068
rect 6231 14028 6276 14056
rect 6270 14016 6276 14028
rect 6328 14016 6334 14068
rect 6546 14056 6552 14068
rect 6507 14028 6552 14056
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 8849 14059 8907 14065
rect 8849 14056 8861 14059
rect 8536 14028 8861 14056
rect 8536 14016 8542 14028
rect 8849 14025 8861 14028
rect 8895 14025 8907 14059
rect 8849 14019 8907 14025
rect 10134 14016 10140 14068
rect 10192 14056 10198 14068
rect 10413 14059 10471 14065
rect 10413 14056 10425 14059
rect 10192 14028 10425 14056
rect 10192 14016 10198 14028
rect 10413 14025 10425 14028
rect 10459 14025 10471 14059
rect 10413 14019 10471 14025
rect 14734 14016 14740 14068
rect 14792 14056 14798 14068
rect 15749 14059 15807 14065
rect 15749 14056 15761 14059
rect 14792 14028 15761 14056
rect 14792 14016 14798 14028
rect 15749 14025 15761 14028
rect 15795 14025 15807 14059
rect 15749 14019 15807 14025
rect 16022 14016 16028 14068
rect 16080 14056 16086 14068
rect 16393 14059 16451 14065
rect 16393 14056 16405 14059
rect 16080 14028 16405 14056
rect 16080 14016 16086 14028
rect 16393 14025 16405 14028
rect 16439 14056 16451 14059
rect 16482 14056 16488 14068
rect 16439 14028 16488 14056
rect 16439 14025 16451 14028
rect 16393 14019 16451 14025
rect 16482 14016 16488 14028
rect 16540 14016 16546 14068
rect 17497 14059 17555 14065
rect 17497 14025 17509 14059
rect 17543 14056 17555 14059
rect 17586 14056 17592 14068
rect 17543 14028 17592 14056
rect 17543 14025 17555 14028
rect 17497 14019 17555 14025
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 17862 14056 17868 14068
rect 17823 14028 17868 14056
rect 17862 14016 17868 14028
rect 17920 14016 17926 14068
rect 19153 14059 19211 14065
rect 19153 14056 19165 14059
rect 18524 14028 19165 14056
rect 5534 13920 5540 13932
rect 4080 13892 5540 13920
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13852 2927 13855
rect 2958 13852 2964 13864
rect 2915 13824 2964 13852
rect 2915 13821 2927 13824
rect 2869 13815 2927 13821
rect 2958 13812 2964 13824
rect 3016 13852 3022 13864
rect 4080 13852 4108 13892
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 5626 13880 5632 13932
rect 5684 13920 5690 13932
rect 5813 13923 5871 13929
rect 5813 13920 5825 13923
rect 5684 13892 5825 13920
rect 5684 13880 5690 13892
rect 5813 13889 5825 13892
rect 5859 13920 5871 13923
rect 6288 13920 6316 14016
rect 5859 13892 6316 13920
rect 6564 13920 6592 14016
rect 12434 13948 12440 14000
rect 12492 13988 12498 14000
rect 12492 13960 12537 13988
rect 12492 13948 12498 13960
rect 17402 13948 17408 14000
rect 17460 13988 17466 14000
rect 18049 13991 18107 13997
rect 18049 13988 18061 13991
rect 17460 13960 18061 13988
rect 17460 13948 17466 13960
rect 18049 13957 18061 13960
rect 18095 13957 18107 13991
rect 18049 13951 18107 13957
rect 6564 13892 6960 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 3016 13824 4108 13852
rect 3016 13812 3022 13824
rect 5350 13812 5356 13864
rect 5408 13852 5414 13864
rect 6822 13852 6828 13864
rect 5408 13824 5488 13852
rect 6783 13824 6828 13852
rect 5408 13812 5414 13824
rect 3136 13787 3194 13793
rect 3136 13753 3148 13787
rect 3182 13784 3194 13787
rect 3602 13784 3608 13796
rect 3182 13756 3608 13784
rect 3182 13753 3194 13756
rect 3136 13747 3194 13753
rect 3602 13744 3608 13756
rect 3660 13744 3666 13796
rect 5460 13784 5488 13824
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 6932 13852 6960 13892
rect 8386 13880 8392 13932
rect 8444 13920 8450 13932
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 8444 13892 8493 13920
rect 8444 13880 8450 13892
rect 8481 13889 8493 13892
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13920 10839 13923
rect 12158 13920 12164 13932
rect 10827 13892 12020 13920
rect 12119 13892 12164 13920
rect 10827 13889 10839 13892
rect 10781 13883 10839 13889
rect 7098 13861 7104 13864
rect 7081 13855 7104 13861
rect 7081 13852 7093 13855
rect 6932 13824 7093 13852
rect 7081 13821 7093 13824
rect 7156 13852 7162 13864
rect 9033 13855 9091 13861
rect 7156 13824 7229 13852
rect 7081 13815 7104 13821
rect 7098 13812 7104 13815
rect 7156 13812 7162 13824
rect 9033 13821 9045 13855
rect 9079 13852 9091 13855
rect 9766 13852 9772 13864
rect 9079 13824 9772 13852
rect 9079 13821 9091 13824
rect 9033 13815 9091 13821
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 11882 13852 11888 13864
rect 11843 13824 11888 13852
rect 11882 13812 11888 13824
rect 11940 13812 11946 13864
rect 11992 13852 12020 13892
rect 12158 13880 12164 13892
rect 12216 13920 12222 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12216 13892 13001 13920
rect 12216 13880 12222 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 13998 13920 14004 13932
rect 13959 13892 14004 13920
rect 12989 13883 13047 13889
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 16942 13920 16948 13932
rect 16903 13892 16948 13920
rect 16942 13880 16948 13892
rect 17000 13880 17006 13932
rect 18524 13929 18552 14028
rect 19153 14025 19165 14028
rect 19199 14056 19211 14059
rect 20346 14056 20352 14068
rect 19199 14028 20352 14056
rect 19199 14025 19211 14028
rect 19153 14019 19211 14025
rect 20346 14016 20352 14028
rect 20404 14016 20410 14068
rect 20990 14056 20996 14068
rect 20951 14028 20996 14056
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 21818 14056 21824 14068
rect 21779 14028 21824 14056
rect 21818 14016 21824 14028
rect 21876 14016 21882 14068
rect 22094 14016 22100 14068
rect 22152 14056 22158 14068
rect 23106 14056 23112 14068
rect 22152 14028 22197 14056
rect 23067 14028 23112 14056
rect 22152 14016 22158 14028
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 23474 14056 23480 14068
rect 23435 14028 23480 14056
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 21453 13991 21511 13997
rect 21453 13957 21465 13991
rect 21499 13988 21511 13991
rect 21910 13988 21916 14000
rect 21499 13960 21916 13988
rect 21499 13957 21511 13960
rect 21453 13951 21511 13957
rect 21910 13948 21916 13960
rect 21968 13948 21974 14000
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13889 18567 13923
rect 18509 13883 18567 13889
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 12434 13852 12440 13864
rect 11992 13824 12440 13852
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12544 13824 12909 13852
rect 5537 13787 5595 13793
rect 5537 13784 5549 13787
rect 5460 13756 5549 13784
rect 5537 13753 5549 13756
rect 5583 13753 5595 13787
rect 5537 13747 5595 13753
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 9278 13787 9336 13793
rect 9278 13784 9290 13787
rect 9180 13756 9290 13784
rect 9180 13744 9186 13756
rect 9278 13753 9290 13756
rect 9324 13753 9336 13787
rect 11238 13784 11244 13796
rect 11199 13756 11244 13784
rect 9278 13747 9336 13753
rect 11238 13744 11244 13756
rect 11296 13744 11302 13796
rect 12250 13744 12256 13796
rect 12308 13784 12314 13796
rect 12544 13784 12572 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 14366 13852 14372 13864
rect 14327 13824 14372 13852
rect 12897 13815 12955 13821
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 14642 13861 14648 13864
rect 14636 13852 14648 13861
rect 14603 13824 14648 13852
rect 14636 13815 14648 13824
rect 14642 13812 14648 13815
rect 14700 13812 14706 13864
rect 16669 13855 16727 13861
rect 16669 13821 16681 13855
rect 16715 13852 16727 13855
rect 17402 13852 17408 13864
rect 16715 13824 17408 13852
rect 16715 13821 16727 13824
rect 16669 13815 16727 13821
rect 17402 13812 17408 13824
rect 17460 13812 17466 13864
rect 17862 13812 17868 13864
rect 17920 13852 17926 13864
rect 18616 13852 18644 13883
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 19610 13920 19616 13932
rect 19300 13892 19616 13920
rect 19300 13880 19306 13892
rect 19610 13880 19616 13892
rect 19668 13920 19674 13932
rect 20165 13923 20223 13929
rect 20165 13920 20177 13923
rect 19668 13892 20177 13920
rect 19668 13880 19674 13892
rect 20165 13889 20177 13892
rect 20211 13889 20223 13923
rect 23492 13920 23520 14016
rect 23492 13892 23796 13920
rect 20165 13883 20223 13889
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 17920 13824 18644 13852
rect 18708 13824 19533 13852
rect 17920 13812 17926 13824
rect 12308 13756 12572 13784
rect 12308 13744 12314 13756
rect 12618 13744 12624 13796
rect 12676 13784 12682 13796
rect 13909 13787 13967 13793
rect 13909 13784 13921 13787
rect 12676 13756 13921 13784
rect 12676 13744 12682 13756
rect 13909 13753 13921 13756
rect 13955 13753 13967 13787
rect 13909 13747 13967 13753
rect 18598 13744 18604 13796
rect 18656 13784 18662 13796
rect 18708 13784 18736 13824
rect 19521 13821 19533 13824
rect 19567 13852 19579 13855
rect 20073 13855 20131 13861
rect 20073 13852 20085 13855
rect 19567 13824 20085 13852
rect 19567 13821 19579 13824
rect 19521 13815 19579 13821
rect 20073 13821 20085 13824
rect 20119 13852 20131 13855
rect 20254 13852 20260 13864
rect 20119 13824 20260 13852
rect 20119 13821 20131 13824
rect 20073 13815 20131 13821
rect 20254 13812 20260 13824
rect 20312 13812 20318 13864
rect 21913 13855 21971 13861
rect 21913 13821 21925 13855
rect 21959 13852 21971 13855
rect 22002 13852 22008 13864
rect 21959 13824 22008 13852
rect 21959 13821 21971 13824
rect 21913 13815 21971 13821
rect 22002 13812 22008 13824
rect 22060 13812 22066 13864
rect 22741 13855 22799 13861
rect 22741 13821 22753 13855
rect 22787 13852 22799 13855
rect 23382 13852 23388 13864
rect 22787 13824 23388 13852
rect 22787 13821 22799 13824
rect 22741 13815 22799 13821
rect 23382 13812 23388 13824
rect 23440 13812 23446 13864
rect 23658 13852 23664 13864
rect 23619 13824 23664 13852
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 23768 13852 23796 13892
rect 23917 13855 23975 13861
rect 23917 13852 23929 13855
rect 23768 13824 23929 13852
rect 23917 13821 23929 13824
rect 23963 13821 23975 13855
rect 23917 13815 23975 13821
rect 18656 13756 18736 13784
rect 18656 13744 18662 13756
rect 19334 13744 19340 13796
rect 19392 13784 19398 13796
rect 19981 13787 20039 13793
rect 19981 13784 19993 13787
rect 19392 13756 19993 13784
rect 19392 13744 19398 13756
rect 19981 13753 19993 13756
rect 20027 13753 20039 13787
rect 19981 13747 20039 13753
rect 3234 13716 3240 13728
rect 2792 13688 3240 13716
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 4430 13676 4436 13728
rect 4488 13716 4494 13728
rect 5166 13716 5172 13728
rect 4488 13688 5172 13716
rect 4488 13676 4494 13688
rect 5166 13676 5172 13688
rect 5224 13716 5230 13728
rect 5629 13719 5687 13725
rect 5629 13716 5641 13719
rect 5224 13688 5641 13716
rect 5224 13676 5230 13688
rect 5629 13685 5641 13688
rect 5675 13685 5687 13719
rect 5629 13679 5687 13685
rect 8205 13719 8263 13725
rect 8205 13685 8217 13719
rect 8251 13716 8263 13719
rect 8478 13716 8484 13728
rect 8251 13688 8484 13716
rect 8251 13685 8263 13688
rect 8205 13679 8263 13685
rect 8478 13676 8484 13688
rect 8536 13676 8542 13728
rect 11149 13719 11207 13725
rect 11149 13685 11161 13719
rect 11195 13716 11207 13719
rect 11974 13716 11980 13728
rect 11195 13688 11980 13716
rect 11195 13685 11207 13688
rect 11149 13679 11207 13685
rect 11974 13676 11980 13688
rect 12032 13676 12038 13728
rect 12526 13676 12532 13728
rect 12584 13716 12590 13728
rect 12805 13719 12863 13725
rect 12805 13716 12817 13719
rect 12584 13688 12817 13716
rect 12584 13676 12590 13688
rect 12805 13685 12817 13688
rect 12851 13716 12863 13719
rect 13449 13719 13507 13725
rect 13449 13716 13461 13719
rect 12851 13688 13461 13716
rect 12851 13685 12863 13688
rect 12805 13679 12863 13685
rect 13449 13685 13461 13688
rect 13495 13685 13507 13719
rect 13814 13716 13820 13728
rect 13775 13688 13820 13716
rect 13449 13679 13507 13685
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 18230 13676 18236 13728
rect 18288 13716 18294 13728
rect 18417 13719 18475 13725
rect 18417 13716 18429 13719
rect 18288 13688 18429 13716
rect 18288 13676 18294 13688
rect 18417 13685 18429 13688
rect 18463 13685 18475 13719
rect 18417 13679 18475 13685
rect 18690 13676 18696 13728
rect 18748 13716 18754 13728
rect 19613 13719 19671 13725
rect 19613 13716 19625 13719
rect 18748 13688 19625 13716
rect 18748 13676 18754 13688
rect 19613 13685 19625 13688
rect 19659 13685 19671 13719
rect 25038 13716 25044 13728
rect 24999 13688 25044 13716
rect 19613 13679 19671 13685
rect 25038 13676 25044 13688
rect 25096 13676 25102 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1762 13472 1768 13524
rect 1820 13512 1826 13524
rect 2409 13515 2467 13521
rect 2409 13512 2421 13515
rect 1820 13484 2421 13512
rect 1820 13472 1826 13484
rect 2409 13481 2421 13484
rect 2455 13481 2467 13515
rect 2409 13475 2467 13481
rect 2590 13472 2596 13524
rect 2648 13512 2654 13524
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2648 13484 2881 13512
rect 2648 13472 2654 13484
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 2869 13475 2927 13481
rect 3786 13472 3792 13524
rect 3844 13512 3850 13524
rect 4433 13515 4491 13521
rect 4433 13512 4445 13515
rect 3844 13484 4445 13512
rect 3844 13472 3850 13484
rect 4433 13481 4445 13484
rect 4479 13512 4491 13515
rect 4890 13512 4896 13524
rect 4479 13484 4896 13512
rect 4479 13481 4491 13484
rect 4433 13475 4491 13481
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 5166 13512 5172 13524
rect 5127 13484 5172 13512
rect 5166 13472 5172 13484
rect 5224 13472 5230 13524
rect 5626 13512 5632 13524
rect 5587 13484 5632 13512
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 7098 13512 7104 13524
rect 7059 13484 7104 13512
rect 7098 13472 7104 13484
rect 7156 13472 7162 13524
rect 9122 13512 9128 13524
rect 9083 13484 9128 13512
rect 9122 13472 9128 13484
rect 9180 13472 9186 13524
rect 9493 13515 9551 13521
rect 9493 13481 9505 13515
rect 9539 13512 9551 13515
rect 9766 13512 9772 13524
rect 9539 13484 9772 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 10045 13515 10103 13521
rect 10045 13481 10057 13515
rect 10091 13512 10103 13515
rect 10686 13512 10692 13524
rect 10091 13484 10692 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 2317 13447 2375 13453
rect 2317 13413 2329 13447
rect 2363 13444 2375 13447
rect 2682 13444 2688 13456
rect 2363 13416 2688 13444
rect 2363 13413 2375 13416
rect 2317 13407 2375 13413
rect 2682 13404 2688 13416
rect 2740 13404 2746 13456
rect 3878 13444 3884 13456
rect 3839 13416 3884 13444
rect 3878 13404 3884 13416
rect 3936 13404 3942 13456
rect 3970 13404 3976 13456
rect 4028 13444 4034 13456
rect 4246 13444 4252 13456
rect 4028 13416 4252 13444
rect 4028 13404 4034 13416
rect 4246 13404 4252 13416
rect 4304 13444 4310 13456
rect 4525 13447 4583 13453
rect 4525 13444 4537 13447
rect 4304 13416 4537 13444
rect 4304 13404 4310 13416
rect 4525 13413 4537 13416
rect 4571 13413 4583 13447
rect 6822 13444 6828 13456
rect 4525 13407 4583 13413
rect 5736 13416 6828 13444
rect 2498 13336 2504 13388
rect 2556 13376 2562 13388
rect 5736 13385 5764 13416
rect 6822 13404 6828 13416
rect 6880 13404 6886 13456
rect 8018 13404 8024 13456
rect 8076 13444 8082 13456
rect 8297 13447 8355 13453
rect 8297 13444 8309 13447
rect 8076 13416 8309 13444
rect 8076 13404 8082 13416
rect 8297 13413 8309 13416
rect 8343 13444 8355 13447
rect 10060 13444 10088 13475
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 11885 13515 11943 13521
rect 11885 13481 11897 13515
rect 11931 13512 11943 13515
rect 11974 13512 11980 13524
rect 11931 13484 11980 13512
rect 11931 13481 11943 13484
rect 11885 13475 11943 13481
rect 11974 13472 11980 13484
rect 12032 13472 12038 13524
rect 12618 13512 12624 13524
rect 12579 13484 12624 13512
rect 12618 13472 12624 13484
rect 12676 13512 12682 13524
rect 15289 13515 15347 13521
rect 12676 13484 12848 13512
rect 12676 13472 12682 13484
rect 8343 13416 10088 13444
rect 8343 13413 8355 13416
rect 8297 13407 8355 13413
rect 5994 13385 6000 13388
rect 2777 13379 2835 13385
rect 2777 13376 2789 13379
rect 2556 13348 2789 13376
rect 2556 13336 2562 13348
rect 2777 13345 2789 13348
rect 2823 13345 2835 13379
rect 2777 13339 2835 13345
rect 5721 13379 5779 13385
rect 5721 13345 5733 13379
rect 5767 13345 5779 13379
rect 5988 13376 6000 13385
rect 5955 13348 6000 13376
rect 5721 13339 5779 13345
rect 5988 13339 6000 13348
rect 5994 13336 6000 13339
rect 6052 13336 6058 13388
rect 10761 13379 10819 13385
rect 10761 13376 10773 13379
rect 10244 13348 10773 13376
rect 10244 13320 10272 13348
rect 10761 13345 10773 13348
rect 10807 13345 10819 13379
rect 10761 13339 10819 13345
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 12492 13348 12725 13376
rect 12492 13336 12498 13348
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 2958 13308 2964 13320
rect 2919 13280 2964 13308
rect 2958 13268 2964 13280
rect 3016 13308 3022 13320
rect 4154 13308 4160 13320
rect 3016 13280 4160 13308
rect 3016 13268 3022 13280
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 4890 13308 4896 13320
rect 4755 13280 4896 13308
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 8294 13268 8300 13320
rect 8352 13308 8358 13320
rect 8389 13311 8447 13317
rect 8389 13308 8401 13311
rect 8352 13280 8401 13308
rect 8352 13268 8358 13280
rect 8389 13277 8401 13280
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 10134 13308 10140 13320
rect 8536 13280 8581 13308
rect 10095 13280 10140 13308
rect 8536 13268 8542 13280
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 10505 13311 10563 13317
rect 10284 13280 10329 13308
rect 10284 13268 10290 13280
rect 10505 13277 10517 13311
rect 10551 13277 10563 13311
rect 10505 13271 10563 13277
rect 4062 13240 4068 13252
rect 4023 13212 4068 13240
rect 4062 13200 4068 13212
rect 4120 13200 4126 13252
rect 6822 13200 6828 13252
rect 6880 13240 6886 13252
rect 7469 13243 7527 13249
rect 7469 13240 7481 13243
rect 6880 13212 7481 13240
rect 6880 13200 6886 13212
rect 7469 13209 7481 13212
rect 7515 13240 7527 13243
rect 7834 13240 7840 13252
rect 7515 13212 7840 13240
rect 7515 13209 7527 13212
rect 7469 13203 7527 13209
rect 7834 13200 7840 13212
rect 7892 13200 7898 13252
rect 9766 13200 9772 13252
rect 9824 13240 9830 13252
rect 10042 13240 10048 13252
rect 9824 13212 10048 13240
rect 9824 13200 9830 13212
rect 10042 13200 10048 13212
rect 10100 13240 10106 13252
rect 10520 13240 10548 13271
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 12820 13308 12848 13484
rect 15289 13481 15301 13515
rect 15335 13512 15347 13515
rect 15930 13512 15936 13524
rect 15335 13484 15936 13512
rect 15335 13481 15347 13484
rect 15289 13475 15347 13481
rect 15930 13472 15936 13484
rect 15988 13472 15994 13524
rect 16393 13515 16451 13521
rect 16393 13481 16405 13515
rect 16439 13512 16451 13515
rect 16482 13512 16488 13524
rect 16439 13484 16488 13512
rect 16439 13481 16451 13484
rect 16393 13475 16451 13481
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 16758 13512 16764 13524
rect 16719 13484 16764 13512
rect 16758 13472 16764 13484
rect 16816 13472 16822 13524
rect 16850 13472 16856 13524
rect 16908 13512 16914 13524
rect 17402 13512 17408 13524
rect 16908 13484 16953 13512
rect 17363 13484 17408 13512
rect 16908 13472 16914 13484
rect 17402 13472 17408 13484
rect 17460 13472 17466 13524
rect 17773 13515 17831 13521
rect 17773 13481 17785 13515
rect 17819 13512 17831 13515
rect 18230 13512 18236 13524
rect 17819 13484 18236 13512
rect 17819 13481 17831 13484
rect 17773 13475 17831 13481
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 18322 13472 18328 13524
rect 18380 13512 18386 13524
rect 18601 13515 18659 13521
rect 18601 13512 18613 13515
rect 18380 13484 18613 13512
rect 18380 13472 18386 13484
rect 18601 13481 18613 13484
rect 18647 13512 18659 13515
rect 18690 13512 18696 13524
rect 18647 13484 18696 13512
rect 18647 13481 18659 13484
rect 18601 13475 18659 13481
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 19797 13515 19855 13521
rect 19797 13481 19809 13515
rect 19843 13512 19855 13515
rect 20622 13512 20628 13524
rect 19843 13484 20628 13512
rect 19843 13481 19855 13484
rect 19797 13475 19855 13481
rect 20622 13472 20628 13484
rect 20680 13472 20686 13524
rect 21634 13512 21640 13524
rect 21595 13484 21640 13512
rect 21634 13472 21640 13484
rect 21692 13472 21698 13524
rect 22741 13515 22799 13521
rect 22741 13481 22753 13515
rect 22787 13512 22799 13515
rect 23198 13512 23204 13524
rect 22787 13484 23204 13512
rect 22787 13481 22799 13484
rect 22741 13475 22799 13481
rect 23198 13472 23204 13484
rect 23256 13472 23262 13524
rect 23290 13472 23296 13524
rect 23348 13512 23354 13524
rect 23658 13512 23664 13524
rect 23348 13484 23664 13512
rect 23348 13472 23354 13484
rect 23658 13472 23664 13484
rect 23716 13472 23722 13524
rect 24854 13512 24860 13524
rect 24815 13484 24860 13512
rect 24854 13472 24860 13484
rect 24912 13472 24918 13524
rect 25501 13515 25559 13521
rect 25501 13481 25513 13515
rect 25547 13512 25559 13515
rect 26050 13512 26056 13524
rect 25547 13484 26056 13512
rect 25547 13481 25559 13484
rect 25501 13475 25559 13481
rect 26050 13472 26056 13484
rect 26108 13472 26114 13524
rect 14274 13404 14280 13456
rect 14332 13444 14338 13456
rect 14550 13444 14556 13456
rect 14332 13416 14556 13444
rect 14332 13404 14338 13416
rect 14550 13404 14556 13416
rect 14608 13404 14614 13456
rect 15657 13447 15715 13453
rect 15657 13413 15669 13447
rect 15703 13444 15715 13447
rect 15746 13444 15752 13456
rect 15703 13416 15752 13444
rect 15703 13413 15715 13416
rect 15657 13407 15715 13413
rect 15746 13404 15752 13416
rect 15804 13404 15810 13456
rect 18046 13376 18052 13388
rect 18007 13348 18052 13376
rect 18046 13336 18052 13348
rect 18104 13376 18110 13388
rect 18414 13376 18420 13388
rect 18104 13348 18420 13376
rect 18104 13336 18110 13348
rect 18414 13336 18420 13348
rect 18472 13376 18478 13388
rect 20530 13376 20536 13388
rect 18472 13348 20536 13376
rect 18472 13336 18478 13348
rect 20530 13336 20536 13348
rect 20588 13336 20594 13388
rect 21453 13379 21511 13385
rect 21453 13345 21465 13379
rect 21499 13376 21511 13379
rect 21910 13376 21916 13388
rect 21499 13348 21916 13376
rect 21499 13345 21511 13348
rect 21453 13339 21511 13345
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 22554 13376 22560 13388
rect 22515 13348 22560 13376
rect 22554 13336 22560 13348
rect 22612 13336 22618 13388
rect 22646 13336 22652 13388
rect 22704 13376 22710 13388
rect 23198 13376 23204 13388
rect 22704 13348 23204 13376
rect 22704 13336 22710 13348
rect 23198 13336 23204 13348
rect 23256 13336 23262 13388
rect 24026 13376 24032 13388
rect 23987 13348 24032 13376
rect 24026 13336 24032 13348
rect 24084 13336 24090 13388
rect 25314 13376 25320 13388
rect 25275 13348 25320 13376
rect 25314 13336 25320 13348
rect 25372 13336 25378 13388
rect 15749 13311 15807 13317
rect 15749 13308 15761 13311
rect 12676 13280 12848 13308
rect 15028 13280 15761 13308
rect 12676 13268 12682 13280
rect 10100 13212 10548 13240
rect 10100 13200 10106 13212
rect 13814 13200 13820 13252
rect 13872 13240 13878 13252
rect 14001 13243 14059 13249
rect 14001 13240 14013 13243
rect 13872 13212 14013 13240
rect 13872 13200 13878 13212
rect 14001 13209 14013 13212
rect 14047 13209 14059 13243
rect 14001 13203 14059 13209
rect 1946 13172 1952 13184
rect 1907 13144 1952 13172
rect 1946 13132 1952 13144
rect 2004 13132 2010 13184
rect 3513 13175 3571 13181
rect 3513 13141 3525 13175
rect 3559 13172 3571 13175
rect 3602 13172 3608 13184
rect 3559 13144 3608 13172
rect 3559 13141 3571 13144
rect 3513 13135 3571 13141
rect 3602 13132 3608 13144
rect 3660 13132 3666 13184
rect 7926 13172 7932 13184
rect 7887 13144 7932 13172
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 9677 13175 9735 13181
rect 9677 13141 9689 13175
rect 9723 13172 9735 13175
rect 11146 13172 11152 13184
rect 9723 13144 11152 13172
rect 9723 13141 9735 13144
rect 9677 13135 9735 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 12250 13172 12256 13184
rect 12211 13144 12256 13172
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 14550 13132 14556 13184
rect 14608 13172 14614 13184
rect 15028 13181 15056 13280
rect 15749 13277 15761 13280
rect 15795 13277 15807 13311
rect 15749 13271 15807 13277
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 18690 13308 18696 13320
rect 15896 13280 15941 13308
rect 18651 13280 18696 13308
rect 15896 13268 15902 13280
rect 18690 13268 18696 13280
rect 18748 13268 18754 13320
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 19150 13308 19156 13320
rect 18923 13280 19156 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 19150 13268 19156 13280
rect 19208 13268 19214 13320
rect 24210 13308 24216 13320
rect 24171 13280 24216 13308
rect 24210 13268 24216 13280
rect 24268 13268 24274 13320
rect 17770 13200 17776 13252
rect 17828 13240 17834 13252
rect 17865 13243 17923 13249
rect 17865 13240 17877 13243
rect 17828 13212 17877 13240
rect 17828 13200 17834 13212
rect 17865 13209 17877 13212
rect 17911 13240 17923 13243
rect 18230 13240 18236 13252
rect 17911 13212 18236 13240
rect 17911 13209 17923 13212
rect 17865 13203 17923 13209
rect 18230 13200 18236 13212
rect 18288 13240 18294 13252
rect 19245 13243 19303 13249
rect 19245 13240 19257 13243
rect 18288 13212 19257 13240
rect 18288 13200 18294 13212
rect 19245 13209 19257 13212
rect 19291 13240 19303 13243
rect 19886 13240 19892 13252
rect 19291 13212 19892 13240
rect 19291 13209 19303 13212
rect 19245 13203 19303 13209
rect 19886 13200 19892 13212
rect 19944 13200 19950 13252
rect 15013 13175 15071 13181
rect 15013 13172 15025 13175
rect 14608 13144 15025 13172
rect 14608 13132 14614 13144
rect 15013 13141 15025 13144
rect 15059 13141 15071 13175
rect 15013 13135 15071 13141
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 19613 13175 19671 13181
rect 19613 13172 19625 13175
rect 19392 13144 19625 13172
rect 19392 13132 19398 13144
rect 19613 13141 19625 13144
rect 19659 13141 19671 13175
rect 19613 13135 19671 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 4249 12971 4307 12977
rect 4249 12968 4261 12971
rect 2832 12940 4261 12968
rect 2832 12928 2838 12940
rect 4249 12937 4261 12940
rect 4295 12937 4307 12971
rect 4249 12931 4307 12937
rect 5813 12971 5871 12977
rect 5813 12937 5825 12971
rect 5859 12968 5871 12971
rect 5994 12968 6000 12980
rect 5859 12940 6000 12968
rect 5859 12937 5871 12940
rect 5813 12931 5871 12937
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 6086 12928 6092 12980
rect 6144 12968 6150 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 6144 12940 6837 12968
rect 6144 12928 6150 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 8018 12968 8024 12980
rect 7979 12940 8024 12968
rect 6825 12931 6883 12937
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 9309 12971 9367 12977
rect 9309 12937 9321 12971
rect 9355 12968 9367 12971
rect 10226 12968 10232 12980
rect 9355 12940 10232 12968
rect 9355 12937 9367 12940
rect 9309 12931 9367 12937
rect 10226 12928 10232 12940
rect 10284 12928 10290 12980
rect 10321 12971 10379 12977
rect 10321 12937 10333 12971
rect 10367 12968 10379 12971
rect 10686 12968 10692 12980
rect 10367 12940 10692 12968
rect 10367 12937 10379 12940
rect 10321 12931 10379 12937
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 14366 12968 14372 12980
rect 13004 12940 14372 12968
rect 2501 12903 2559 12909
rect 2501 12869 2513 12903
rect 2547 12900 2559 12903
rect 2958 12900 2964 12912
rect 2547 12872 2964 12900
rect 2547 12869 2559 12872
rect 2501 12863 2559 12869
rect 2958 12860 2964 12872
rect 3016 12860 3022 12912
rect 5261 12903 5319 12909
rect 5261 12900 5273 12903
rect 3252 12872 5273 12900
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12832 2191 12835
rect 3050 12832 3056 12844
rect 2179 12804 3056 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 3050 12792 3056 12804
rect 3108 12832 3114 12844
rect 3252 12841 3280 12872
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 3108 12804 3249 12832
rect 3108 12792 3114 12804
rect 3237 12801 3249 12804
rect 3283 12801 3295 12835
rect 3786 12832 3792 12844
rect 3747 12804 3792 12832
rect 3237 12795 3295 12801
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12832 4215 12835
rect 4246 12832 4252 12844
rect 4203 12804 4252 12832
rect 4203 12801 4215 12804
rect 4157 12795 4215 12801
rect 4246 12792 4252 12804
rect 4304 12792 4310 12844
rect 4706 12832 4712 12844
rect 4667 12804 4712 12832
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 4816 12841 4844 12872
rect 5261 12869 5273 12872
rect 5307 12869 5319 12903
rect 5261 12863 5319 12869
rect 8294 12860 8300 12912
rect 8352 12900 8358 12912
rect 9585 12903 9643 12909
rect 9585 12900 9597 12903
rect 8352 12872 9597 12900
rect 8352 12860 8358 12872
rect 9585 12869 9597 12872
rect 9631 12900 9643 12903
rect 10134 12900 10140 12912
rect 9631 12872 10140 12900
rect 9631 12869 9643 12872
rect 9585 12863 9643 12869
rect 10134 12860 10140 12872
rect 10192 12860 10198 12912
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12801 4859 12835
rect 4801 12795 4859 12801
rect 4890 12792 4896 12844
rect 4948 12832 4954 12844
rect 6273 12835 6331 12841
rect 6273 12832 6285 12835
rect 4948 12804 6285 12832
rect 4948 12792 4954 12804
rect 6273 12801 6285 12804
rect 6319 12832 6331 12835
rect 7469 12835 7527 12841
rect 7469 12832 7481 12835
rect 6319 12804 7481 12832
rect 6319 12801 6331 12804
rect 6273 12795 6331 12801
rect 7469 12801 7481 12804
rect 7515 12832 7527 12835
rect 8662 12832 8668 12844
rect 7515 12804 7880 12832
rect 8623 12804 8668 12832
rect 7515 12801 7527 12804
rect 7469 12795 7527 12801
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 1486 12764 1492 12776
rect 1443 12736 1492 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1486 12724 1492 12736
rect 1544 12724 1550 12776
rect 4062 12724 4068 12776
rect 4120 12764 4126 12776
rect 4617 12767 4675 12773
rect 4617 12764 4629 12767
rect 4120 12736 4629 12764
rect 4120 12724 4126 12736
rect 4617 12733 4629 12736
rect 4663 12733 4675 12767
rect 7282 12764 7288 12776
rect 7195 12736 7288 12764
rect 4617 12727 4675 12733
rect 7282 12724 7288 12736
rect 7340 12764 7346 12776
rect 7742 12764 7748 12776
rect 7340 12736 7748 12764
rect 7340 12724 7346 12736
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 1946 12656 1952 12708
rect 2004 12696 2010 12708
rect 3053 12699 3111 12705
rect 3053 12696 3065 12699
rect 2004 12668 3065 12696
rect 2004 12656 2010 12668
rect 3053 12665 3065 12668
rect 3099 12665 3111 12699
rect 3053 12659 3111 12665
rect 6641 12699 6699 12705
rect 6641 12665 6653 12699
rect 6687 12696 6699 12699
rect 7190 12696 7196 12708
rect 6687 12668 7196 12696
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 7190 12656 7196 12668
rect 7248 12656 7254 12708
rect 7852 12696 7880 12804
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 10244 12832 10272 12928
rect 11238 12832 11244 12844
rect 10244 12804 11244 12832
rect 11238 12792 11244 12804
rect 11296 12832 11302 12844
rect 13004 12841 13032 12940
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 14737 12971 14795 12977
rect 14737 12937 14749 12971
rect 14783 12968 14795 12971
rect 15013 12971 15071 12977
rect 15013 12968 15025 12971
rect 14783 12940 15025 12968
rect 14783 12937 14795 12940
rect 14737 12931 14795 12937
rect 15013 12937 15025 12940
rect 15059 12937 15071 12971
rect 15013 12931 15071 12937
rect 15197 12971 15255 12977
rect 15197 12937 15209 12971
rect 15243 12968 15255 12971
rect 16114 12968 16120 12980
rect 15243 12940 16120 12968
rect 15243 12937 15255 12940
rect 15197 12931 15255 12937
rect 11333 12835 11391 12841
rect 11333 12832 11345 12835
rect 11296 12804 11345 12832
rect 11296 12792 11302 12804
rect 11333 12801 11345 12804
rect 11379 12832 11391 12835
rect 11793 12835 11851 12841
rect 11793 12832 11805 12835
rect 11379 12804 11805 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 11793 12801 11805 12804
rect 11839 12801 11851 12835
rect 11793 12795 11851 12801
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 15028 12832 15056 12931
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 17497 12971 17555 12977
rect 17497 12937 17509 12971
rect 17543 12968 17555 12971
rect 18322 12968 18328 12980
rect 17543 12940 18328 12968
rect 17543 12937 17555 12940
rect 17497 12931 17555 12937
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 18874 12968 18880 12980
rect 18748 12940 18880 12968
rect 18748 12928 18754 12940
rect 18874 12928 18880 12940
rect 18932 12928 18938 12980
rect 19886 12968 19892 12980
rect 19847 12940 19892 12968
rect 19886 12928 19892 12940
rect 19944 12928 19950 12980
rect 21266 12968 21272 12980
rect 21227 12940 21272 12968
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 22646 12968 22652 12980
rect 22607 12940 22652 12968
rect 22646 12928 22652 12940
rect 22704 12928 22710 12980
rect 22830 12928 22836 12980
rect 22888 12968 22894 12980
rect 23017 12971 23075 12977
rect 23017 12968 23029 12971
rect 22888 12940 23029 12968
rect 22888 12928 22894 12940
rect 23017 12937 23029 12940
rect 23063 12937 23075 12971
rect 23017 12931 23075 12937
rect 17865 12903 17923 12909
rect 17865 12869 17877 12903
rect 17911 12900 17923 12903
rect 19150 12900 19156 12912
rect 17911 12872 19156 12900
rect 17911 12869 17923 12872
rect 17865 12863 17923 12869
rect 19150 12860 19156 12872
rect 19208 12860 19214 12912
rect 19242 12860 19248 12912
rect 19300 12860 19306 12912
rect 21174 12860 21180 12912
rect 21232 12900 21238 12912
rect 21545 12903 21603 12909
rect 21545 12900 21557 12903
rect 21232 12872 21557 12900
rect 21232 12860 21238 12872
rect 21545 12869 21557 12872
rect 21591 12869 21603 12903
rect 21545 12863 21603 12869
rect 22373 12903 22431 12909
rect 22373 12869 22385 12903
rect 22419 12900 22431 12903
rect 22554 12900 22560 12912
rect 22419 12872 22560 12900
rect 22419 12869 22431 12872
rect 22373 12863 22431 12869
rect 22554 12860 22560 12872
rect 22612 12860 22618 12912
rect 15749 12835 15807 12841
rect 15749 12832 15761 12835
rect 15028 12804 15761 12832
rect 12989 12795 13047 12801
rect 15749 12801 15761 12804
rect 15795 12832 15807 12835
rect 15838 12832 15844 12844
rect 15795 12804 15844 12832
rect 15795 12801 15807 12804
rect 15749 12795 15807 12801
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 16758 12832 16764 12844
rect 16719 12804 16764 12832
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 19260 12832 19288 12860
rect 19429 12835 19487 12841
rect 19429 12832 19441 12835
rect 19260 12804 19441 12832
rect 19429 12801 19441 12804
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 23477 12835 23535 12841
rect 23477 12801 23489 12835
rect 23523 12832 23535 12835
rect 23523 12804 23796 12832
rect 23523 12801 23535 12804
rect 23477 12795 23535 12801
rect 8570 12764 8576 12776
rect 8531 12736 8576 12764
rect 8570 12724 8576 12736
rect 8628 12724 8634 12776
rect 9582 12724 9588 12776
rect 9640 12724 9646 12776
rect 13262 12773 13268 12776
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12764 10747 12767
rect 13256 12764 13268 12773
rect 10735 12736 11468 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 9600 12696 9628 12724
rect 7852 12668 9628 12696
rect 9769 12699 9827 12705
rect 9769 12665 9781 12699
rect 9815 12696 9827 12699
rect 10962 12696 10968 12708
rect 9815 12668 10968 12696
rect 9815 12665 9827 12668
rect 9769 12659 9827 12665
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 11149 12699 11207 12705
rect 11149 12665 11161 12699
rect 11195 12696 11207 12699
rect 11330 12696 11336 12708
rect 11195 12668 11336 12696
rect 11195 12665 11207 12668
rect 11149 12659 11207 12665
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 2498 12588 2504 12640
rect 2556 12628 2562 12640
rect 2685 12631 2743 12637
rect 2685 12628 2697 12631
rect 2556 12600 2697 12628
rect 2556 12588 2562 12600
rect 2685 12597 2697 12600
rect 2731 12597 2743 12631
rect 2685 12591 2743 12597
rect 3142 12588 3148 12640
rect 3200 12628 3206 12640
rect 3200 12600 3245 12628
rect 3200 12588 3206 12600
rect 7834 12588 7840 12640
rect 7892 12628 7898 12640
rect 8389 12631 8447 12637
rect 8389 12628 8401 12631
rect 7892 12600 8401 12628
rect 7892 12588 7898 12600
rect 8389 12597 8401 12600
rect 8435 12628 8447 12631
rect 9950 12628 9956 12640
rect 8435 12600 9956 12628
rect 8435 12597 8447 12600
rect 8389 12591 8447 12597
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10781 12631 10839 12637
rect 10781 12597 10793 12631
rect 10827 12628 10839 12631
rect 11054 12628 11060 12640
rect 10827 12600 11060 12628
rect 10827 12597 10839 12600
rect 10781 12591 10839 12597
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 11241 12631 11299 12637
rect 11241 12597 11253 12631
rect 11287 12628 11299 12631
rect 11440 12628 11468 12736
rect 13188 12736 13268 12764
rect 12253 12699 12311 12705
rect 12253 12665 12265 12699
rect 12299 12696 12311 12699
rect 13188 12696 13216 12736
rect 13256 12727 13268 12736
rect 13262 12724 13268 12727
rect 13320 12724 13326 12776
rect 21266 12724 21272 12776
rect 21324 12764 21330 12776
rect 21361 12767 21419 12773
rect 21361 12764 21373 12767
rect 21324 12736 21373 12764
rect 21324 12724 21330 12736
rect 21361 12733 21373 12736
rect 21407 12733 21419 12767
rect 21910 12764 21916 12776
rect 21871 12736 21916 12764
rect 21361 12727 21419 12733
rect 21910 12724 21916 12736
rect 21968 12724 21974 12776
rect 22465 12767 22523 12773
rect 22465 12733 22477 12767
rect 22511 12764 22523 12767
rect 22830 12764 22836 12776
rect 22511 12736 22836 12764
rect 22511 12733 22523 12736
rect 22465 12727 22523 12733
rect 22830 12724 22836 12736
rect 22888 12724 22894 12776
rect 23106 12724 23112 12776
rect 23164 12764 23170 12776
rect 23658 12764 23664 12776
rect 23164 12736 23664 12764
rect 23164 12724 23170 12736
rect 23658 12724 23664 12736
rect 23716 12724 23722 12776
rect 23768 12764 23796 12804
rect 23928 12767 23986 12773
rect 23928 12764 23940 12767
rect 23768 12736 23940 12764
rect 23928 12733 23940 12736
rect 23974 12764 23986 12767
rect 25038 12764 25044 12776
rect 23974 12736 25044 12764
rect 23974 12733 23986 12736
rect 23928 12727 23986 12733
rect 25038 12724 25044 12736
rect 25096 12724 25102 12776
rect 12299 12668 13216 12696
rect 15565 12699 15623 12705
rect 12299 12665 12311 12668
rect 12253 12659 12311 12665
rect 15565 12665 15577 12699
rect 15611 12696 15623 12699
rect 16114 12696 16120 12708
rect 15611 12668 16120 12696
rect 15611 12665 15623 12668
rect 15565 12659 15623 12665
rect 16114 12656 16120 12668
rect 16172 12696 16178 12708
rect 16577 12699 16635 12705
rect 16577 12696 16589 12699
rect 16172 12668 16589 12696
rect 16172 12656 16178 12668
rect 16577 12665 16589 12668
rect 16623 12665 16635 12699
rect 16577 12659 16635 12665
rect 18417 12699 18475 12705
rect 18417 12665 18429 12699
rect 18463 12696 18475 12699
rect 18506 12696 18512 12708
rect 18463 12668 18512 12696
rect 18463 12665 18475 12668
rect 18417 12659 18475 12665
rect 18506 12656 18512 12668
rect 18564 12696 18570 12708
rect 19245 12699 19303 12705
rect 19245 12696 19257 12699
rect 18564 12668 19257 12696
rect 18564 12656 18570 12668
rect 19245 12665 19257 12668
rect 19291 12665 19303 12699
rect 19245 12659 19303 12665
rect 11514 12628 11520 12640
rect 11287 12600 11520 12628
rect 11287 12597 11299 12600
rect 11241 12591 11299 12597
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12713 12631 12771 12637
rect 12713 12628 12725 12631
rect 12492 12600 12725 12628
rect 12492 12588 12498 12600
rect 12713 12597 12725 12600
rect 12759 12597 12771 12631
rect 12713 12591 12771 12597
rect 13538 12588 13544 12640
rect 13596 12628 13602 12640
rect 14369 12631 14427 12637
rect 14369 12628 14381 12631
rect 13596 12600 14381 12628
rect 13596 12588 13602 12600
rect 14369 12597 14381 12600
rect 14415 12597 14427 12631
rect 14369 12591 14427 12597
rect 15654 12588 15660 12640
rect 15712 12628 15718 12640
rect 16209 12631 16267 12637
rect 16209 12628 16221 12631
rect 15712 12600 16221 12628
rect 15712 12588 15718 12600
rect 16209 12597 16221 12600
rect 16255 12597 16267 12631
rect 18690 12628 18696 12640
rect 18651 12600 18696 12628
rect 16209 12591 16267 12597
rect 18690 12588 18696 12600
rect 18748 12628 18754 12640
rect 19058 12628 19064 12640
rect 18748 12600 19064 12628
rect 18748 12588 18754 12600
rect 19058 12588 19064 12600
rect 19116 12628 19122 12640
rect 19337 12631 19395 12637
rect 19337 12628 19349 12631
rect 19116 12600 19349 12628
rect 19116 12588 19122 12600
rect 19337 12597 19349 12600
rect 19383 12597 19395 12631
rect 19337 12591 19395 12597
rect 25041 12631 25099 12637
rect 25041 12597 25053 12631
rect 25087 12628 25099 12631
rect 25130 12628 25136 12640
rect 25087 12600 25136 12628
rect 25087 12597 25099 12600
rect 25041 12591 25099 12597
rect 25130 12588 25136 12600
rect 25188 12588 25194 12640
rect 25314 12628 25320 12640
rect 25275 12600 25320 12628
rect 25314 12588 25320 12600
rect 25372 12588 25378 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1486 12384 1492 12436
rect 1544 12424 1550 12436
rect 1581 12427 1639 12433
rect 1581 12424 1593 12427
rect 1544 12396 1593 12424
rect 1544 12384 1550 12396
rect 1581 12393 1593 12396
rect 1627 12393 1639 12427
rect 1581 12387 1639 12393
rect 1946 12384 1952 12436
rect 2004 12424 2010 12436
rect 2409 12427 2467 12433
rect 2409 12424 2421 12427
rect 2004 12396 2421 12424
rect 2004 12384 2010 12396
rect 2409 12393 2421 12396
rect 2455 12393 2467 12427
rect 4062 12424 4068 12436
rect 4023 12396 4068 12424
rect 2409 12387 2467 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4338 12384 4344 12436
rect 4396 12424 4402 12436
rect 4525 12427 4583 12433
rect 4525 12424 4537 12427
rect 4396 12396 4537 12424
rect 4396 12384 4402 12396
rect 4525 12393 4537 12396
rect 4571 12393 4583 12427
rect 5166 12424 5172 12436
rect 5127 12396 5172 12424
rect 4525 12387 4583 12393
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 6273 12427 6331 12433
rect 6273 12393 6285 12427
rect 6319 12424 6331 12427
rect 6822 12424 6828 12436
rect 6319 12396 6828 12424
rect 6319 12393 6331 12396
rect 6273 12387 6331 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 6917 12427 6975 12433
rect 6917 12393 6929 12427
rect 6963 12424 6975 12427
rect 7282 12424 7288 12436
rect 6963 12396 7288 12424
rect 6963 12393 6975 12396
rect 6917 12387 6975 12393
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 8021 12427 8079 12433
rect 8021 12393 8033 12427
rect 8067 12424 8079 12427
rect 8202 12424 8208 12436
rect 8067 12396 8208 12424
rect 8067 12393 8079 12396
rect 8021 12387 8079 12393
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 8389 12427 8447 12433
rect 8389 12393 8401 12427
rect 8435 12424 8447 12427
rect 8478 12424 8484 12436
rect 8435 12396 8484 12424
rect 8435 12393 8447 12396
rect 8389 12387 8447 12393
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 8665 12427 8723 12433
rect 8665 12424 8677 12427
rect 8628 12396 8677 12424
rect 8628 12384 8634 12396
rect 8665 12393 8677 12396
rect 8711 12393 8723 12427
rect 8665 12387 8723 12393
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10413 12427 10471 12433
rect 10413 12424 10425 12427
rect 10100 12396 10425 12424
rect 10100 12384 10106 12396
rect 10413 12393 10425 12396
rect 10459 12393 10471 12427
rect 10413 12387 10471 12393
rect 11425 12427 11483 12433
rect 11425 12393 11437 12427
rect 11471 12424 11483 12427
rect 12250 12424 12256 12436
rect 11471 12396 12256 12424
rect 11471 12393 11483 12396
rect 11425 12387 11483 12393
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 12986 12424 12992 12436
rect 12947 12396 12992 12424
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 14645 12427 14703 12433
rect 14645 12393 14657 12427
rect 14691 12424 14703 12427
rect 14734 12424 14740 12436
rect 14691 12396 14740 12424
rect 14691 12393 14703 12396
rect 14645 12387 14703 12393
rect 14734 12384 14740 12396
rect 14792 12424 14798 12436
rect 15013 12427 15071 12433
rect 15013 12424 15025 12427
rect 14792 12396 15025 12424
rect 14792 12384 14798 12396
rect 15013 12393 15025 12396
rect 15059 12393 15071 12427
rect 15013 12387 15071 12393
rect 15289 12427 15347 12433
rect 15289 12393 15301 12427
rect 15335 12424 15347 12427
rect 15746 12424 15752 12436
rect 15335 12396 15752 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 2038 12316 2044 12368
rect 2096 12356 2102 12368
rect 2777 12359 2835 12365
rect 2777 12356 2789 12359
rect 2096 12328 2789 12356
rect 2096 12316 2102 12328
rect 2777 12325 2789 12328
rect 2823 12325 2835 12359
rect 2777 12319 2835 12325
rect 3513 12359 3571 12365
rect 3513 12325 3525 12359
rect 3559 12356 3571 12359
rect 4080 12356 4108 12384
rect 3559 12328 4108 12356
rect 9953 12359 10011 12365
rect 3559 12325 3571 12328
rect 3513 12319 3571 12325
rect 9953 12325 9965 12359
rect 9999 12356 10011 12359
rect 10686 12356 10692 12368
rect 9999 12328 10692 12356
rect 9999 12325 10011 12328
rect 9953 12319 10011 12325
rect 10686 12316 10692 12328
rect 10744 12316 10750 12368
rect 11146 12316 11152 12368
rect 11204 12356 11210 12368
rect 11885 12359 11943 12365
rect 11885 12356 11897 12359
rect 11204 12328 11897 12356
rect 11204 12316 11210 12328
rect 11885 12325 11897 12328
rect 11931 12325 11943 12359
rect 15028 12356 15056 12387
rect 15746 12384 15752 12396
rect 15804 12424 15810 12436
rect 16669 12427 16727 12433
rect 16669 12424 16681 12427
rect 15804 12396 16681 12424
rect 15804 12384 15810 12396
rect 16669 12393 16681 12396
rect 16715 12393 16727 12427
rect 16669 12387 16727 12393
rect 17957 12427 18015 12433
rect 17957 12393 17969 12427
rect 18003 12424 18015 12427
rect 18046 12424 18052 12436
rect 18003 12396 18052 12424
rect 18003 12393 18015 12396
rect 17957 12387 18015 12393
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 18325 12427 18383 12433
rect 18325 12393 18337 12427
rect 18371 12424 18383 12427
rect 18874 12424 18880 12436
rect 18371 12396 18880 12424
rect 18371 12393 18383 12396
rect 18325 12387 18383 12393
rect 18874 12384 18880 12396
rect 18932 12384 18938 12436
rect 19518 12424 19524 12436
rect 19479 12396 19524 12424
rect 19518 12384 19524 12396
rect 19576 12384 19582 12436
rect 21726 12384 21732 12436
rect 21784 12424 21790 12436
rect 21821 12427 21879 12433
rect 21821 12424 21833 12427
rect 21784 12396 21833 12424
rect 21784 12384 21790 12396
rect 21821 12393 21833 12396
rect 21867 12393 21879 12427
rect 21821 12387 21879 12393
rect 22925 12427 22983 12433
rect 22925 12393 22937 12427
rect 22971 12424 22983 12427
rect 23198 12424 23204 12436
rect 22971 12396 23204 12424
rect 22971 12393 22983 12396
rect 22925 12387 22983 12393
rect 23198 12384 23204 12396
rect 23256 12384 23262 12436
rect 23290 12384 23296 12436
rect 23348 12424 23354 12436
rect 23474 12424 23480 12436
rect 23348 12396 23480 12424
rect 23348 12384 23354 12396
rect 23474 12384 23480 12396
rect 23532 12384 23538 12436
rect 24210 12384 24216 12436
rect 24268 12424 24274 12436
rect 24670 12424 24676 12436
rect 24268 12396 24676 12424
rect 24268 12384 24274 12396
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 18601 12359 18659 12365
rect 15028 12328 15792 12356
rect 11885 12319 11943 12325
rect 2130 12248 2136 12300
rect 2188 12288 2194 12300
rect 2866 12288 2872 12300
rect 2188 12260 2872 12288
rect 2188 12248 2194 12260
rect 2866 12248 2872 12260
rect 2924 12248 2930 12300
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12288 4491 12291
rect 4614 12288 4620 12300
rect 4479 12260 4620 12288
rect 4479 12257 4491 12260
rect 4433 12251 4491 12257
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 11054 12248 11060 12300
rect 11112 12288 11118 12300
rect 11422 12288 11428 12300
rect 11112 12260 11428 12288
rect 11112 12248 11118 12260
rect 11422 12248 11428 12260
rect 11480 12288 11486 12300
rect 11793 12291 11851 12297
rect 11793 12288 11805 12291
rect 11480 12260 11805 12288
rect 11480 12248 11486 12260
rect 11793 12257 11805 12260
rect 11839 12257 11851 12291
rect 13354 12288 13360 12300
rect 13315 12260 13360 12288
rect 11793 12251 11851 12257
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12288 13507 12291
rect 13722 12288 13728 12300
rect 13495 12260 13728 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 13722 12248 13728 12260
rect 13780 12288 13786 12300
rect 14274 12288 14280 12300
rect 13780 12260 14280 12288
rect 13780 12248 13786 12260
rect 14274 12248 14280 12260
rect 14332 12248 14338 12300
rect 15286 12248 15292 12300
rect 15344 12288 15350 12300
rect 15562 12288 15568 12300
rect 15344 12260 15568 12288
rect 15344 12248 15350 12260
rect 15562 12248 15568 12260
rect 15620 12288 15626 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15620 12260 15669 12288
rect 15620 12248 15626 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15764 12288 15792 12328
rect 18601 12325 18613 12359
rect 18647 12356 18659 12359
rect 19334 12356 19340 12368
rect 18647 12328 19340 12356
rect 18647 12325 18659 12328
rect 18601 12319 18659 12325
rect 19334 12316 19340 12328
rect 19392 12316 19398 12368
rect 23106 12316 23112 12368
rect 23164 12356 23170 12368
rect 23661 12359 23719 12365
rect 23661 12356 23673 12359
rect 23164 12328 23673 12356
rect 23164 12316 23170 12328
rect 23661 12325 23673 12328
rect 23707 12325 23719 12359
rect 24118 12356 24124 12368
rect 23661 12319 23719 12325
rect 23952 12328 24124 12356
rect 17221 12291 17279 12297
rect 15764 12260 15884 12288
rect 15657 12251 15715 12257
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 3602 12220 3608 12232
rect 3099 12192 3608 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3602 12180 3608 12192
rect 3660 12220 3666 12232
rect 4706 12220 4712 12232
rect 3660 12192 4712 12220
rect 3660 12180 3666 12192
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 5534 12220 5540 12232
rect 5447 12192 5540 12220
rect 5534 12180 5540 12192
rect 5592 12220 5598 12232
rect 5813 12223 5871 12229
rect 5813 12220 5825 12223
rect 5592 12192 5825 12220
rect 5592 12180 5598 12192
rect 5813 12189 5825 12192
rect 5859 12189 5871 12223
rect 11238 12220 11244 12232
rect 11199 12192 11244 12220
rect 5813 12183 5871 12189
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 11974 12220 11980 12232
rect 11935 12192 11980 12220
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 13538 12180 13544 12232
rect 13596 12220 13602 12232
rect 15746 12220 15752 12232
rect 13596 12192 13641 12220
rect 15707 12192 15752 12220
rect 13596 12180 13602 12192
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15856 12229 15884 12260
rect 17221 12257 17233 12291
rect 17267 12288 17279 12291
rect 17494 12288 17500 12300
rect 17267 12260 17500 12288
rect 17267 12257 17279 12260
rect 17221 12251 17279 12257
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 19150 12288 19156 12300
rect 19111 12260 19156 12288
rect 19150 12248 19156 12260
rect 19208 12248 19214 12300
rect 21634 12288 21640 12300
rect 21595 12260 21640 12288
rect 21634 12248 21640 12260
rect 21692 12248 21698 12300
rect 22741 12291 22799 12297
rect 22741 12257 22753 12291
rect 22787 12288 22799 12291
rect 23014 12288 23020 12300
rect 22787 12260 23020 12288
rect 22787 12257 22799 12260
rect 22741 12251 22799 12257
rect 23014 12248 23020 12260
rect 23072 12248 23078 12300
rect 23952 12232 23980 12328
rect 24118 12316 24124 12328
rect 24176 12316 24182 12368
rect 24213 12291 24271 12297
rect 24213 12257 24225 12291
rect 24259 12288 24271 12291
rect 24854 12288 24860 12300
rect 24259 12260 24860 12288
rect 24259 12257 24271 12260
rect 24213 12251 24271 12257
rect 24854 12248 24860 12260
rect 24912 12288 24918 12300
rect 25409 12291 25467 12297
rect 25409 12288 25421 12291
rect 24912 12260 25421 12288
rect 24912 12248 24918 12260
rect 25409 12257 25421 12260
rect 25455 12257 25467 12291
rect 25409 12251 25467 12257
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12220 15899 12223
rect 16298 12220 16304 12232
rect 15887 12192 16304 12220
rect 15887 12189 15899 12192
rect 15841 12183 15899 12189
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 17310 12220 17316 12232
rect 17271 12192 17316 12220
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17402 12180 17408 12232
rect 17460 12220 17466 12232
rect 17460 12192 17505 12220
rect 17460 12180 17466 12192
rect 18506 12180 18512 12232
rect 18564 12220 18570 12232
rect 19242 12220 19248 12232
rect 18564 12192 19248 12220
rect 18564 12180 18570 12192
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 19794 12220 19800 12232
rect 19755 12192 19800 12220
rect 19794 12180 19800 12192
rect 19852 12180 19858 12232
rect 23934 12180 23940 12232
rect 23992 12180 23998 12232
rect 24118 12180 24124 12232
rect 24176 12220 24182 12232
rect 24305 12223 24363 12229
rect 24305 12220 24317 12223
rect 24176 12192 24317 12220
rect 24176 12180 24182 12192
rect 24305 12189 24317 12192
rect 24351 12189 24363 12223
rect 24305 12183 24363 12189
rect 24394 12180 24400 12232
rect 24452 12220 24458 12232
rect 24489 12223 24547 12229
rect 24489 12220 24501 12223
rect 24452 12192 24501 12220
rect 24452 12180 24458 12192
rect 24489 12189 24501 12192
rect 24535 12220 24547 12223
rect 24670 12220 24676 12232
rect 24535 12192 24676 12220
rect 24535 12189 24547 12192
rect 24489 12183 24547 12189
rect 24670 12180 24676 12192
rect 24728 12180 24734 12232
rect 2317 12155 2375 12161
rect 2317 12121 2329 12155
rect 2363 12152 2375 12155
rect 3142 12152 3148 12164
rect 2363 12124 3148 12152
rect 2363 12121 2375 12124
rect 2317 12115 2375 12121
rect 3142 12112 3148 12124
rect 3200 12112 3206 12164
rect 3881 12155 3939 12161
rect 3881 12121 3893 12155
rect 3927 12152 3939 12155
rect 4890 12152 4896 12164
rect 3927 12124 4896 12152
rect 3927 12121 3939 12124
rect 3881 12115 3939 12121
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 10873 12155 10931 12161
rect 10873 12121 10885 12155
rect 10919 12152 10931 12155
rect 11330 12152 11336 12164
rect 10919 12124 11336 12152
rect 10919 12121 10931 12124
rect 10873 12115 10931 12121
rect 11330 12112 11336 12124
rect 11388 12152 11394 12164
rect 12066 12152 12072 12164
rect 11388 12124 12072 12152
rect 11388 12112 11394 12124
rect 12066 12112 12072 12124
rect 12124 12152 12130 12164
rect 13262 12152 13268 12164
rect 12124 12124 13268 12152
rect 12124 12112 12130 12124
rect 13262 12112 13268 12124
rect 13320 12112 13326 12164
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 24026 12152 24032 12164
rect 23891 12124 24032 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 24026 12112 24032 12124
rect 24084 12152 24090 12164
rect 24857 12155 24915 12161
rect 24857 12152 24869 12155
rect 24084 12124 24869 12152
rect 24084 12112 24090 12124
rect 24857 12121 24869 12124
rect 24903 12121 24915 12155
rect 24857 12115 24915 12121
rect 12805 12087 12863 12093
rect 12805 12053 12817 12087
rect 12851 12084 12863 12087
rect 13446 12084 13452 12096
rect 12851 12056 13452 12084
rect 12851 12053 12863 12056
rect 12805 12047 12863 12053
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 14090 12084 14096 12096
rect 14051 12056 14096 12084
rect 14090 12044 14096 12056
rect 14148 12084 14154 12096
rect 14366 12084 14372 12096
rect 14148 12056 14372 12084
rect 14148 12044 14154 12056
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 16850 12084 16856 12096
rect 16811 12056 16856 12084
rect 16850 12044 16856 12056
rect 16908 12044 16914 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1394 11840 1400 11892
rect 1452 11880 1458 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 1452 11852 1593 11880
rect 1452 11840 1458 11852
rect 1581 11849 1593 11852
rect 1627 11849 1639 11883
rect 2038 11880 2044 11892
rect 1999 11852 2044 11880
rect 1581 11843 1639 11849
rect 2038 11840 2044 11852
rect 2096 11840 2102 11892
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 2409 11883 2467 11889
rect 2409 11880 2421 11883
rect 2188 11852 2421 11880
rect 2188 11840 2194 11852
rect 2409 11849 2421 11852
rect 2455 11849 2467 11883
rect 2409 11843 2467 11849
rect 3053 11883 3111 11889
rect 3053 11849 3065 11883
rect 3099 11880 3111 11883
rect 3142 11880 3148 11892
rect 3099 11852 3148 11880
rect 3099 11849 3111 11852
rect 3053 11843 3111 11849
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 4338 11840 4344 11892
rect 4396 11880 4402 11892
rect 4433 11883 4491 11889
rect 4433 11880 4445 11883
rect 4396 11852 4445 11880
rect 4396 11840 4402 11852
rect 4433 11849 4445 11852
rect 4479 11849 4491 11883
rect 4433 11843 4491 11849
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 4801 11883 4859 11889
rect 4801 11880 4813 11883
rect 4764 11852 4813 11880
rect 4764 11840 4770 11852
rect 4801 11849 4813 11852
rect 4847 11849 4859 11883
rect 11146 11880 11152 11892
rect 11107 11852 11152 11880
rect 4801 11843 4859 11849
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 11974 11880 11980 11892
rect 11563 11852 11980 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 11974 11840 11980 11852
rect 12032 11840 12038 11892
rect 12618 11840 12624 11892
rect 12676 11880 12682 11892
rect 12713 11883 12771 11889
rect 12713 11880 12725 11883
rect 12676 11852 12725 11880
rect 12676 11840 12682 11852
rect 12713 11849 12725 11852
rect 12759 11849 12771 11883
rect 14550 11880 14556 11892
rect 14511 11852 14556 11880
rect 12713 11843 12771 11849
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 16114 11880 16120 11892
rect 16075 11852 16120 11880
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 17221 11883 17279 11889
rect 17221 11849 17233 11883
rect 17267 11880 17279 11883
rect 17310 11880 17316 11892
rect 17267 11852 17316 11880
rect 17267 11849 17279 11852
rect 17221 11843 17279 11849
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 17494 11880 17500 11892
rect 17455 11852 17500 11880
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 18230 11880 18236 11892
rect 18191 11852 18236 11880
rect 18230 11840 18236 11852
rect 18288 11880 18294 11892
rect 18601 11883 18659 11889
rect 18601 11880 18613 11883
rect 18288 11852 18613 11880
rect 18288 11840 18294 11852
rect 18601 11849 18613 11852
rect 18647 11849 18659 11883
rect 18601 11843 18659 11849
rect 21634 11840 21640 11892
rect 21692 11880 21698 11892
rect 21913 11883 21971 11889
rect 21913 11880 21925 11883
rect 21692 11852 21925 11880
rect 21692 11840 21698 11852
rect 21913 11849 21925 11852
rect 21959 11849 21971 11883
rect 21913 11843 21971 11849
rect 22278 11840 22284 11892
rect 22336 11880 22342 11892
rect 22649 11883 22707 11889
rect 22649 11880 22661 11883
rect 22336 11852 22661 11880
rect 22336 11840 22342 11852
rect 22649 11849 22661 11852
rect 22695 11849 22707 11883
rect 23014 11880 23020 11892
rect 22975 11852 23020 11880
rect 22649 11843 22707 11849
rect 23014 11840 23020 11852
rect 23072 11840 23078 11892
rect 23477 11883 23535 11889
rect 23477 11849 23489 11883
rect 23523 11880 23535 11883
rect 24854 11880 24860 11892
rect 23523 11852 24860 11880
rect 23523 11849 23535 11852
rect 23477 11843 23535 11849
rect 24854 11840 24860 11852
rect 24912 11840 24918 11892
rect 25038 11880 25044 11892
rect 24999 11852 25044 11880
rect 25038 11840 25044 11852
rect 25096 11840 25102 11892
rect 4157 11815 4215 11821
rect 4157 11781 4169 11815
rect 4203 11812 4215 11815
rect 4614 11812 4620 11824
rect 4203 11784 4620 11812
rect 4203 11781 4215 11784
rect 4157 11775 4215 11781
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 11054 11772 11060 11824
rect 11112 11812 11118 11824
rect 12161 11815 12219 11821
rect 12161 11812 12173 11815
rect 11112 11784 12173 11812
rect 11112 11772 11118 11784
rect 12161 11781 12173 11784
rect 12207 11812 12219 11815
rect 13354 11812 13360 11824
rect 12207 11784 13360 11812
rect 12207 11781 12219 11784
rect 12161 11775 12219 11781
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 16298 11772 16304 11824
rect 16356 11812 16362 11824
rect 25056 11812 25084 11840
rect 16356 11784 16712 11812
rect 16356 11772 16362 11784
rect 3602 11744 3608 11756
rect 3563 11716 3608 11744
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 11793 11747 11851 11753
rect 11793 11744 11805 11747
rect 11296 11716 11805 11744
rect 11296 11704 11302 11716
rect 11793 11713 11805 11716
rect 11839 11744 11851 11747
rect 12342 11744 12348 11756
rect 11839 11716 12348 11744
rect 11839 11713 11851 11716
rect 11793 11707 11851 11713
rect 12342 11704 12348 11716
rect 12400 11744 12406 11756
rect 13265 11747 13323 11753
rect 13265 11744 13277 11747
rect 12400 11716 13277 11744
rect 12400 11704 12406 11716
rect 13265 11713 13277 11716
rect 13311 11744 13323 11747
rect 13538 11744 13544 11756
rect 13311 11716 13544 11744
rect 13311 11713 13323 11716
rect 13265 11707 13323 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 15105 11747 15163 11753
rect 15105 11744 15117 11747
rect 14792 11716 15117 11744
rect 14792 11704 14798 11716
rect 15105 11713 15117 11716
rect 15151 11713 15163 11747
rect 15105 11707 15163 11713
rect 16482 11704 16488 11756
rect 16540 11744 16546 11756
rect 16684 11753 16712 11784
rect 24688 11784 25084 11812
rect 16577 11747 16635 11753
rect 16577 11744 16589 11747
rect 16540 11716 16589 11744
rect 16540 11704 16546 11716
rect 16577 11713 16589 11716
rect 16623 11713 16635 11747
rect 16577 11707 16635 11713
rect 16669 11747 16727 11753
rect 16669 11713 16681 11747
rect 16715 11713 16727 11747
rect 21450 11744 21456 11756
rect 21411 11716 21456 11744
rect 16669 11707 16727 11713
rect 21450 11704 21456 11716
rect 21508 11704 21514 11756
rect 22278 11744 22284 11756
rect 22239 11716 22284 11744
rect 22278 11704 22284 11716
rect 22336 11744 22342 11756
rect 22336 11716 22508 11744
rect 22336 11704 22342 11716
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1670 11676 1676 11688
rect 1443 11648 1676 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 2406 11636 2412 11688
rect 2464 11676 2470 11688
rect 3142 11676 3148 11688
rect 2464 11648 3148 11676
rect 2464 11636 2470 11648
rect 3142 11636 3148 11648
rect 3200 11676 3206 11688
rect 3421 11679 3479 11685
rect 3421 11676 3433 11679
rect 3200 11648 3433 11676
rect 3200 11636 3206 11648
rect 3421 11645 3433 11648
rect 3467 11676 3479 11679
rect 3510 11676 3516 11688
rect 3467 11648 3516 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 13722 11676 13728 11688
rect 13683 11648 13728 11676
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 22480 11685 22508 11716
rect 23842 11704 23848 11756
rect 23900 11744 23906 11756
rect 24026 11744 24032 11756
rect 23900 11716 24032 11744
rect 23900 11704 23906 11716
rect 24026 11704 24032 11716
rect 24084 11704 24090 11756
rect 24688 11753 24716 11784
rect 24673 11747 24731 11753
rect 24673 11713 24685 11747
rect 24719 11713 24731 11747
rect 24673 11707 24731 11713
rect 24946 11704 24952 11756
rect 25004 11744 25010 11756
rect 25593 11747 25651 11753
rect 25593 11744 25605 11747
rect 25004 11716 25605 11744
rect 25004 11704 25010 11716
rect 25593 11713 25605 11716
rect 25639 11713 25651 11747
rect 25593 11707 25651 11713
rect 22465 11679 22523 11685
rect 22465 11645 22477 11679
rect 22511 11645 22523 11679
rect 24397 11679 24455 11685
rect 24397 11676 24409 11679
rect 22465 11639 22523 11645
rect 23860 11648 24409 11676
rect 14734 11568 14740 11620
rect 14792 11608 14798 11620
rect 15013 11611 15071 11617
rect 15013 11608 15025 11611
rect 14792 11580 15025 11608
rect 14792 11568 14798 11580
rect 15013 11577 15025 11580
rect 15059 11577 15071 11611
rect 15013 11571 15071 11577
rect 15657 11611 15715 11617
rect 15657 11577 15669 11611
rect 15703 11608 15715 11611
rect 15746 11608 15752 11620
rect 15703 11580 15752 11608
rect 15703 11577 15715 11580
rect 15657 11571 15715 11577
rect 15746 11568 15752 11580
rect 15804 11568 15810 11620
rect 23860 11552 23888 11648
rect 24397 11645 24409 11648
rect 24443 11645 24455 11679
rect 24397 11639 24455 11645
rect 24118 11608 24124 11620
rect 24031 11580 24124 11608
rect 2961 11543 3019 11549
rect 2961 11509 2973 11543
rect 3007 11540 3019 11543
rect 3234 11540 3240 11552
rect 3007 11512 3240 11540
rect 3007 11509 3019 11512
rect 2961 11503 3019 11509
rect 3234 11500 3240 11512
rect 3292 11540 3298 11552
rect 3513 11543 3571 11549
rect 3513 11540 3525 11543
rect 3292 11512 3525 11540
rect 3292 11500 3298 11512
rect 3513 11509 3525 11512
rect 3559 11540 3571 11543
rect 3970 11540 3976 11552
rect 3559 11512 3976 11540
rect 3559 11509 3571 11512
rect 3513 11503 3571 11509
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 13078 11540 13084 11552
rect 13039 11512 13084 11540
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13173 11543 13231 11549
rect 13173 11509 13185 11543
rect 13219 11540 13231 11543
rect 13446 11540 13452 11552
rect 13219 11512 13452 11540
rect 13219 11509 13231 11512
rect 13173 11503 13231 11509
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 14366 11540 14372 11552
rect 14327 11512 14372 11540
rect 14366 11500 14372 11512
rect 14424 11540 14430 11552
rect 14921 11543 14979 11549
rect 14921 11540 14933 11543
rect 14424 11512 14933 11540
rect 14424 11500 14430 11512
rect 14921 11509 14933 11512
rect 14967 11509 14979 11543
rect 14921 11503 14979 11509
rect 16025 11543 16083 11549
rect 16025 11509 16037 11543
rect 16071 11540 16083 11543
rect 16390 11540 16396 11552
rect 16071 11512 16396 11540
rect 16071 11509 16083 11512
rect 16025 11503 16083 11509
rect 16390 11500 16396 11512
rect 16448 11540 16454 11552
rect 16485 11543 16543 11549
rect 16485 11540 16497 11543
rect 16448 11512 16497 11540
rect 16448 11500 16454 11512
rect 16485 11509 16497 11512
rect 16531 11509 16543 11543
rect 23842 11540 23848 11552
rect 23803 11512 23848 11540
rect 16485 11503 16543 11509
rect 23842 11500 23848 11512
rect 23900 11500 23906 11552
rect 24044 11549 24072 11580
rect 24118 11568 24124 11580
rect 24176 11608 24182 11620
rect 25409 11611 25467 11617
rect 25409 11608 25421 11611
rect 24176 11580 25421 11608
rect 24176 11568 24182 11580
rect 25409 11577 25421 11580
rect 25455 11577 25467 11611
rect 25409 11571 25467 11577
rect 24029 11543 24087 11549
rect 24029 11509 24041 11543
rect 24075 11509 24087 11543
rect 24486 11540 24492 11552
rect 24447 11512 24492 11540
rect 24029 11503 24087 11509
rect 24486 11500 24492 11512
rect 24544 11500 24550 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 2590 11336 2596 11348
rect 2179 11308 2596 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 3142 11336 3148 11348
rect 3103 11308 3148 11336
rect 3142 11296 3148 11308
rect 3200 11296 3206 11348
rect 3513 11339 3571 11345
rect 3513 11305 3525 11339
rect 3559 11336 3571 11339
rect 3602 11336 3608 11348
rect 3559 11308 3608 11336
rect 3559 11305 3571 11308
rect 3513 11299 3571 11305
rect 2501 11271 2559 11277
rect 2501 11237 2513 11271
rect 2547 11268 2559 11271
rect 3528 11268 3556 11299
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 11422 11336 11428 11348
rect 11383 11308 11428 11336
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 12342 11336 12348 11348
rect 12303 11308 12348 11336
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 12989 11339 13047 11345
rect 12989 11336 13001 11339
rect 12584 11308 13001 11336
rect 12584 11296 12590 11308
rect 12989 11305 13001 11308
rect 13035 11305 13047 11339
rect 12989 11299 13047 11305
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 15654 11336 15660 11348
rect 15335 11308 15660 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 16393 11339 16451 11345
rect 16393 11305 16405 11339
rect 16439 11336 16451 11339
rect 16482 11336 16488 11348
rect 16439 11308 16488 11336
rect 16439 11305 16451 11308
rect 16393 11299 16451 11305
rect 16482 11296 16488 11308
rect 16540 11296 16546 11348
rect 16942 11296 16948 11348
rect 17000 11336 17006 11348
rect 17221 11339 17279 11345
rect 17221 11336 17233 11339
rect 17000 11308 17233 11336
rect 17000 11296 17006 11308
rect 17221 11305 17233 11308
rect 17267 11305 17279 11339
rect 17221 11299 17279 11305
rect 22557 11339 22615 11345
rect 22557 11305 22569 11339
rect 22603 11336 22615 11339
rect 22738 11336 22744 11348
rect 22603 11308 22744 11336
rect 22603 11305 22615 11308
rect 22557 11299 22615 11305
rect 22738 11296 22744 11308
rect 22796 11296 22802 11348
rect 23661 11339 23719 11345
rect 23661 11305 23673 11339
rect 23707 11305 23719 11339
rect 23661 11299 23719 11305
rect 24489 11339 24547 11345
rect 24489 11305 24501 11339
rect 24535 11336 24547 11339
rect 24670 11336 24676 11348
rect 24535 11308 24676 11336
rect 24535 11305 24547 11308
rect 24489 11299 24547 11305
rect 2547 11240 3556 11268
rect 12805 11271 12863 11277
rect 2547 11237 2559 11240
rect 2501 11231 2559 11237
rect 12805 11237 12817 11271
rect 12851 11268 12863 11271
rect 13078 11268 13084 11280
rect 12851 11240 13084 11268
rect 12851 11237 12863 11240
rect 12805 11231 12863 11237
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 13357 11271 13415 11277
rect 13357 11237 13369 11271
rect 13403 11268 13415 11271
rect 13446 11268 13452 11280
rect 13403 11240 13452 11268
rect 13403 11237 13415 11240
rect 13357 11231 13415 11237
rect 13446 11228 13452 11240
rect 13504 11228 13510 11280
rect 15105 11271 15163 11277
rect 15105 11237 15117 11271
rect 15151 11268 15163 11271
rect 15562 11268 15568 11280
rect 15151 11240 15568 11268
rect 15151 11237 15163 11240
rect 15105 11231 15163 11237
rect 15562 11228 15568 11240
rect 15620 11228 15626 11280
rect 15749 11271 15807 11277
rect 15749 11237 15761 11271
rect 15795 11268 15807 11271
rect 16114 11268 16120 11280
rect 15795 11240 16120 11268
rect 15795 11237 15807 11240
rect 15749 11231 15807 11237
rect 16114 11228 16120 11240
rect 16172 11268 16178 11280
rect 16850 11268 16856 11280
rect 16172 11240 16856 11268
rect 16172 11228 16178 11240
rect 16850 11228 16856 11240
rect 16908 11228 16914 11280
rect 23676 11268 23704 11299
rect 24670 11296 24676 11308
rect 24728 11296 24734 11348
rect 26326 11268 26332 11280
rect 23676 11240 26332 11268
rect 26326 11228 26332 11240
rect 26384 11228 26390 11280
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11200 14703 11203
rect 14734 11200 14740 11212
rect 14691 11172 14740 11200
rect 14691 11169 14703 11172
rect 14645 11163 14703 11169
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 15378 11160 15384 11212
rect 15436 11200 15442 11212
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 15436 11172 15669 11200
rect 15436 11160 15442 11172
rect 15657 11169 15669 11172
rect 15703 11200 15715 11203
rect 16022 11200 16028 11212
rect 15703 11172 16028 11200
rect 15703 11169 15715 11172
rect 15657 11163 15715 11169
rect 16022 11160 16028 11172
rect 16080 11160 16086 11212
rect 22370 11200 22376 11212
rect 22331 11172 22376 11200
rect 22370 11160 22376 11172
rect 22428 11160 22434 11212
rect 23474 11200 23480 11212
rect 23435 11172 23480 11200
rect 23474 11160 23480 11172
rect 23532 11160 23538 11212
rect 24578 11200 24584 11212
rect 24539 11172 24584 11200
rect 24578 11160 24584 11172
rect 24636 11200 24642 11212
rect 24854 11200 24860 11212
rect 24636 11172 24860 11200
rect 24636 11160 24642 11172
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 13449 11135 13507 11141
rect 13449 11132 13461 11135
rect 13228 11104 13461 11132
rect 13228 11092 13234 11104
rect 13449 11101 13461 11104
rect 13495 11101 13507 11135
rect 13449 11095 13507 11101
rect 13633 11135 13691 11141
rect 13633 11101 13645 11135
rect 13679 11132 13691 11135
rect 13722 11132 13728 11144
rect 13679 11104 13728 11132
rect 13679 11101 13691 11104
rect 13633 11095 13691 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 15746 11092 15752 11144
rect 15804 11132 15810 11144
rect 15933 11135 15991 11141
rect 15933 11132 15945 11135
rect 15804 11104 15945 11132
rect 15804 11092 15810 11104
rect 15933 11101 15945 11104
rect 15979 11132 15991 11135
rect 16298 11132 16304 11144
rect 15979 11104 16304 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16298 11092 16304 11104
rect 16356 11092 16362 11144
rect 24118 11132 24124 11144
rect 24079 11104 24124 11132
rect 24118 11092 24124 11104
rect 24176 11132 24182 11144
rect 24486 11132 24492 11144
rect 24176 11104 24492 11132
rect 24176 11092 24182 11104
rect 24486 11092 24492 11104
rect 24544 11092 24550 11144
rect 14090 11024 14096 11076
rect 14148 11064 14154 11076
rect 14277 11067 14335 11073
rect 14277 11064 14289 11067
rect 14148 11036 14289 11064
rect 14148 11024 14154 11036
rect 14277 11033 14289 11036
rect 14323 11064 14335 11067
rect 14642 11064 14648 11076
rect 14323 11036 14648 11064
rect 14323 11033 14335 11036
rect 14277 11027 14335 11033
rect 14642 11024 14648 11036
rect 14700 11024 14706 11076
rect 16850 11064 16856 11076
rect 16811 11036 16856 11064
rect 16850 11024 16856 11036
rect 16908 11064 16914 11076
rect 17402 11064 17408 11076
rect 16908 11036 17408 11064
rect 16908 11024 16914 11036
rect 17402 11024 17408 11036
rect 17460 11024 17466 11076
rect 23750 11024 23756 11076
rect 23808 11064 23814 11076
rect 24765 11067 24823 11073
rect 24765 11064 24777 11067
rect 23808 11036 24777 11064
rect 23808 11024 23814 11036
rect 24765 11033 24777 11036
rect 24811 11033 24823 11067
rect 24765 11027 24823 11033
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2498 10792 2504 10804
rect 2459 10764 2504 10792
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 13722 10792 13728 10804
rect 13683 10764 13728 10792
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 15378 10792 15384 10804
rect 15339 10764 15384 10792
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 15746 10792 15752 10804
rect 15707 10764 15752 10792
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 16114 10792 16120 10804
rect 16075 10764 16120 10792
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 22370 10792 22376 10804
rect 22331 10764 22376 10792
rect 22370 10752 22376 10764
rect 22428 10752 22434 10804
rect 23474 10752 23480 10804
rect 23532 10792 23538 10804
rect 23845 10795 23903 10801
rect 23845 10792 23857 10795
rect 23532 10764 23857 10792
rect 23532 10752 23538 10764
rect 23845 10761 23857 10764
rect 23891 10761 23903 10795
rect 23845 10755 23903 10761
rect 23934 10752 23940 10804
rect 23992 10792 23998 10804
rect 24765 10795 24823 10801
rect 24765 10792 24777 10795
rect 23992 10764 24777 10792
rect 23992 10752 23998 10764
rect 24765 10761 24777 10764
rect 24811 10761 24823 10795
rect 24765 10755 24823 10761
rect 24854 10752 24860 10804
rect 24912 10792 24918 10804
rect 25133 10795 25191 10801
rect 25133 10792 25145 10795
rect 24912 10764 25145 10792
rect 24912 10752 24918 10764
rect 25133 10761 25145 10764
rect 25179 10792 25191 10795
rect 25774 10792 25780 10804
rect 25179 10764 25780 10792
rect 25179 10761 25191 10764
rect 25133 10755 25191 10761
rect 25774 10752 25780 10764
rect 25832 10752 25838 10804
rect 24394 10656 24400 10668
rect 24355 10628 24400 10656
rect 24394 10616 24400 10628
rect 24452 10616 24458 10668
rect 1394 10588 1400 10600
rect 1355 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10588 1458 10600
rect 1949 10591 2007 10597
rect 1949 10588 1961 10591
rect 1452 10560 1961 10588
rect 1452 10548 1458 10560
rect 1949 10557 1961 10560
rect 1995 10557 2007 10591
rect 24412 10588 24440 10616
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 24412 10560 24593 10588
rect 1949 10551 2007 10557
rect 24581 10557 24593 10560
rect 24627 10557 24639 10591
rect 24581 10551 24639 10557
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 13078 10452 13084 10464
rect 13039 10424 13084 10452
rect 13078 10412 13084 10424
rect 13136 10412 13142 10464
rect 13446 10452 13452 10464
rect 13407 10424 13452 10452
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 14642 10452 14648 10464
rect 14603 10424 14648 10452
rect 14642 10412 14648 10424
rect 14700 10412 14706 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 24762 10248 24768 10260
rect 24723 10220 24768 10248
rect 24762 10208 24768 10220
rect 24820 10208 24826 10260
rect 24581 10115 24639 10121
rect 24581 10081 24593 10115
rect 24627 10112 24639 10115
rect 24670 10112 24676 10124
rect 24627 10084 24676 10112
rect 24627 10081 24639 10084
rect 24581 10075 24639 10081
rect 24670 10072 24676 10084
rect 24728 10072 24734 10124
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 24210 9596 24216 9648
rect 24268 9636 24274 9648
rect 24397 9639 24455 9645
rect 24397 9636 24409 9639
rect 24268 9608 24409 9636
rect 24268 9596 24274 9608
rect 24397 9605 24409 9608
rect 24443 9605 24455 9639
rect 24397 9599 24455 9605
rect 24412 9500 24440 9599
rect 24581 9503 24639 9509
rect 24581 9500 24593 9503
rect 24412 9472 24593 9500
rect 24581 9469 24593 9472
rect 24627 9469 24639 9503
rect 25130 9500 25136 9512
rect 25091 9472 25136 9500
rect 24581 9463 24639 9469
rect 25130 9460 25136 9472
rect 25188 9460 25194 9512
rect 19334 9392 19340 9444
rect 19392 9432 19398 9444
rect 25958 9432 25964 9444
rect 19392 9404 25964 9432
rect 19392 9392 19398 9404
rect 25958 9392 25964 9404
rect 26016 9392 26022 9444
rect 24026 9324 24032 9376
rect 24084 9364 24090 9376
rect 24765 9367 24823 9373
rect 24765 9364 24777 9367
rect 24084 9336 24777 9364
rect 24084 9324 24090 9336
rect 24765 9333 24777 9336
rect 24811 9333 24823 9367
rect 24765 9327 24823 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 9582 8616 9588 8628
rect 1627 8588 9588 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8412 1458 8424
rect 1949 8415 2007 8421
rect 1949 8412 1961 8415
rect 1452 8384 1961 8412
rect 1452 8372 1458 8384
rect 1949 8381 1961 8384
rect 1995 8381 2007 8415
rect 1949 8375 2007 8381
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 9582 5896 9588 5908
rect 1627 5868 9588 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1452 5324 1593 5352
rect 1452 5312 1458 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 1581 5315 1639 5321
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 566 2796 572 2848
rect 624 2836 630 2848
rect 3326 2836 3332 2848
rect 624 2808 3332 2836
rect 624 2796 630 2808
rect 3326 2796 3332 2808
rect 3384 2796 3390 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 12434 2632 12440 2644
rect 12395 2604 12440 2632
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 14090 2632 14096 2644
rect 14051 2604 14096 2632
rect 14090 2592 14096 2604
rect 14148 2592 14154 2644
rect 12452 2564 12480 2592
rect 12958 2567 13016 2573
rect 12958 2564 12970 2567
rect 12452 2536 12970 2564
rect 12958 2533 12970 2536
rect 13004 2533 13016 2567
rect 12958 2527 13016 2533
rect 12069 2499 12127 2505
rect 12069 2465 12081 2499
rect 12115 2496 12127 2499
rect 12710 2496 12716 2508
rect 12115 2468 12716 2496
rect 12115 2465 12127 2468
rect 12069 2459 12127 2465
rect 12710 2456 12716 2468
rect 12768 2456 12774 2508
rect 24213 2295 24271 2301
rect 24213 2261 24225 2295
rect 24259 2292 24271 2295
rect 25130 2292 25136 2304
rect 24259 2264 25136 2292
rect 24259 2261 24271 2264
rect 24213 2255 24271 2261
rect 25130 2252 25136 2264
rect 25188 2252 25194 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 9220 27412 9272 27464
rect 9404 27412 9456 27464
rect 26424 27412 26476 27464
rect 26516 27412 26568 27464
rect 3516 27276 3568 27328
rect 4896 27276 4948 27328
rect 11612 26188 11664 26240
rect 18144 26188 18196 26240
rect 13452 26120 13504 26172
rect 22744 26120 22796 26172
rect 10968 25984 11020 26036
rect 24584 25984 24636 26036
rect 4620 25916 4672 25968
rect 19340 25916 19392 25968
rect 12624 25848 12676 25900
rect 25872 25848 25924 25900
rect 10692 25780 10744 25832
rect 18696 25780 18748 25832
rect 1952 25712 2004 25764
rect 20812 25712 20864 25764
rect 8760 25644 8812 25696
rect 19248 25644 19300 25696
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 2780 25440 2832 25492
rect 8760 25483 8812 25492
rect 8760 25449 8769 25483
rect 8769 25449 8803 25483
rect 8803 25449 8812 25483
rect 8760 25440 8812 25449
rect 10692 25440 10744 25492
rect 11612 25483 11664 25492
rect 11612 25449 11621 25483
rect 11621 25449 11655 25483
rect 11655 25449 11664 25483
rect 11612 25440 11664 25449
rect 24768 25483 24820 25492
rect 2320 25304 2372 25356
rect 2596 25304 2648 25356
rect 4344 25304 4396 25356
rect 6000 25304 6052 25356
rect 11244 25372 11296 25424
rect 9956 25304 10008 25356
rect 296 25168 348 25220
rect 1584 25143 1636 25152
rect 1584 25109 1593 25143
rect 1593 25109 1627 25143
rect 1627 25109 1636 25143
rect 1584 25100 1636 25109
rect 6276 25143 6328 25152
rect 6276 25109 6285 25143
rect 6285 25109 6319 25143
rect 6319 25109 6328 25143
rect 6276 25100 6328 25109
rect 7196 25143 7248 25152
rect 7196 25109 7205 25143
rect 7205 25109 7239 25143
rect 7239 25109 7248 25143
rect 7196 25100 7248 25109
rect 9312 25100 9364 25152
rect 11336 25100 11388 25152
rect 12900 25304 12952 25356
rect 13268 25304 13320 25356
rect 14188 25304 14240 25356
rect 16580 25304 16632 25356
rect 18788 25304 18840 25356
rect 22192 25372 22244 25424
rect 22744 25415 22796 25424
rect 22744 25381 22753 25415
rect 22753 25381 22787 25415
rect 22787 25381 22796 25415
rect 22744 25372 22796 25381
rect 24768 25449 24777 25483
rect 24777 25449 24811 25483
rect 24811 25449 24820 25483
rect 24768 25440 24820 25449
rect 27068 25372 27120 25424
rect 20904 25304 20956 25356
rect 21180 25347 21232 25356
rect 21180 25313 21189 25347
rect 21189 25313 21223 25347
rect 21223 25313 21232 25347
rect 21180 25304 21232 25313
rect 22468 25347 22520 25356
rect 22468 25313 22477 25347
rect 22477 25313 22511 25347
rect 22511 25313 22520 25347
rect 22468 25304 22520 25313
rect 24124 25304 24176 25356
rect 24584 25347 24636 25356
rect 24584 25313 24593 25347
rect 24593 25313 24627 25347
rect 24627 25313 24636 25347
rect 24584 25304 24636 25313
rect 12164 25236 12216 25288
rect 15568 25236 15620 25288
rect 16396 25236 16448 25288
rect 17040 25236 17092 25288
rect 18052 25236 18104 25288
rect 19156 25279 19208 25288
rect 19156 25245 19165 25279
rect 19165 25245 19199 25279
rect 19199 25245 19208 25279
rect 19156 25236 19208 25245
rect 21456 25279 21508 25288
rect 21456 25245 21465 25279
rect 21465 25245 21499 25279
rect 21499 25245 21508 25279
rect 21456 25236 21508 25245
rect 12624 25211 12676 25220
rect 12624 25177 12633 25211
rect 12633 25177 12667 25211
rect 12667 25177 12676 25211
rect 12624 25168 12676 25177
rect 17224 25168 17276 25220
rect 25044 25168 25096 25220
rect 12440 25100 12492 25152
rect 14096 25100 14148 25152
rect 15384 25100 15436 25152
rect 15660 25143 15712 25152
rect 15660 25109 15669 25143
rect 15669 25109 15703 25143
rect 15703 25109 15712 25143
rect 15660 25100 15712 25109
rect 16672 25143 16724 25152
rect 16672 25109 16681 25143
rect 16681 25109 16715 25143
rect 16715 25109 16724 25143
rect 16672 25100 16724 25109
rect 18604 25100 18656 25152
rect 19524 25143 19576 25152
rect 19524 25109 19533 25143
rect 19533 25109 19567 25143
rect 19567 25109 19576 25143
rect 19524 25100 19576 25109
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 2688 24939 2740 24948
rect 2688 24905 2697 24939
rect 2697 24905 2731 24939
rect 2731 24905 2740 24939
rect 2688 24896 2740 24905
rect 3792 24939 3844 24948
rect 3792 24905 3801 24939
rect 3801 24905 3835 24939
rect 3835 24905 3844 24939
rect 3792 24896 3844 24905
rect 4896 24939 4948 24948
rect 4896 24905 4905 24939
rect 4905 24905 4939 24939
rect 4939 24905 4948 24939
rect 4896 24896 4948 24905
rect 9312 24896 9364 24948
rect 17224 24896 17276 24948
rect 7196 24760 7248 24812
rect 13360 24828 13412 24880
rect 14924 24828 14976 24880
rect 18052 24896 18104 24948
rect 22468 24896 22520 24948
rect 24124 24896 24176 24948
rect 8392 24760 8444 24812
rect 9496 24803 9548 24812
rect 9496 24769 9505 24803
rect 9505 24769 9539 24803
rect 9539 24769 9548 24803
rect 9496 24760 9548 24769
rect 11244 24803 11296 24812
rect 11244 24769 11253 24803
rect 11253 24769 11287 24803
rect 11287 24769 11296 24803
rect 11244 24760 11296 24769
rect 2320 24692 2372 24744
rect 3148 24735 3200 24744
rect 3148 24701 3157 24735
rect 3157 24701 3191 24735
rect 3191 24701 3200 24735
rect 3148 24692 3200 24701
rect 1584 24599 1636 24608
rect 1584 24565 1593 24599
rect 1593 24565 1627 24599
rect 1627 24565 1636 24599
rect 1584 24556 1636 24565
rect 2412 24599 2464 24608
rect 2412 24565 2421 24599
rect 2421 24565 2455 24599
rect 2455 24565 2464 24599
rect 2412 24556 2464 24565
rect 4344 24692 4396 24744
rect 6000 24624 6052 24676
rect 6368 24624 6420 24676
rect 3700 24556 3752 24608
rect 4252 24556 4304 24608
rect 4712 24556 4764 24608
rect 5448 24556 5500 24608
rect 6920 24599 6972 24608
rect 6920 24565 6929 24599
rect 6929 24565 6963 24599
rect 6963 24565 6972 24599
rect 6920 24556 6972 24565
rect 7932 24692 7984 24744
rect 8300 24735 8352 24744
rect 8300 24701 8309 24735
rect 8309 24701 8343 24735
rect 8343 24701 8352 24735
rect 8300 24692 8352 24701
rect 9128 24692 9180 24744
rect 10876 24624 10928 24676
rect 12992 24692 13044 24744
rect 7748 24556 7800 24608
rect 8484 24599 8536 24608
rect 8484 24565 8493 24599
rect 8493 24565 8527 24599
rect 8527 24565 8536 24599
rect 8484 24556 8536 24565
rect 8944 24599 8996 24608
rect 8944 24565 8953 24599
rect 8953 24565 8987 24599
rect 8987 24565 8996 24599
rect 9956 24599 10008 24608
rect 8944 24556 8996 24565
rect 9956 24565 9965 24599
rect 9965 24565 9999 24599
rect 9999 24565 10008 24599
rect 9956 24556 10008 24565
rect 10784 24556 10836 24608
rect 10968 24599 11020 24608
rect 10968 24565 10977 24599
rect 10977 24565 11011 24599
rect 11011 24565 11020 24599
rect 10968 24556 11020 24565
rect 11888 24556 11940 24608
rect 12164 24599 12216 24608
rect 12164 24565 12173 24599
rect 12173 24565 12207 24599
rect 12207 24565 12216 24599
rect 12164 24556 12216 24565
rect 12808 24599 12860 24608
rect 12808 24565 12817 24599
rect 12817 24565 12851 24599
rect 12851 24565 12860 24599
rect 12808 24556 12860 24565
rect 13268 24556 13320 24608
rect 16488 24692 16540 24744
rect 14372 24667 14424 24676
rect 14372 24633 14381 24667
rect 14381 24633 14415 24667
rect 14415 24633 14424 24667
rect 14372 24624 14424 24633
rect 14280 24556 14332 24608
rect 15108 24556 15160 24608
rect 15568 24599 15620 24608
rect 15568 24565 15577 24599
rect 15577 24565 15611 24599
rect 15611 24565 15620 24599
rect 15568 24556 15620 24565
rect 15936 24556 15988 24608
rect 16028 24556 16080 24608
rect 16396 24556 16448 24608
rect 17040 24556 17092 24608
rect 18604 24803 18656 24812
rect 18604 24769 18613 24803
rect 18613 24769 18647 24803
rect 18647 24769 18656 24803
rect 18604 24760 18656 24769
rect 20076 24828 20128 24880
rect 24768 24828 24820 24880
rect 19340 24760 19392 24812
rect 20444 24760 20496 24812
rect 20536 24760 20588 24812
rect 24860 24760 24912 24812
rect 26056 24760 26108 24812
rect 20168 24624 20220 24676
rect 18604 24556 18656 24608
rect 18788 24556 18840 24608
rect 19984 24599 20036 24608
rect 19984 24565 19993 24599
rect 19993 24565 20027 24599
rect 20027 24565 20036 24599
rect 19984 24556 20036 24565
rect 20720 24556 20772 24608
rect 21180 24556 21232 24608
rect 24032 24692 24084 24744
rect 23112 24624 23164 24676
rect 23388 24556 23440 24608
rect 24676 24556 24728 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 4160 24352 4212 24404
rect 7196 24352 7248 24404
rect 8484 24352 8536 24404
rect 6552 24284 6604 24336
rect 9036 24284 9088 24336
rect 9772 24352 9824 24404
rect 11336 24352 11388 24404
rect 13636 24395 13688 24404
rect 13636 24361 13645 24395
rect 13645 24361 13679 24395
rect 13679 24361 13688 24395
rect 13636 24352 13688 24361
rect 14096 24352 14148 24404
rect 14832 24352 14884 24404
rect 15476 24395 15528 24404
rect 15476 24361 15485 24395
rect 15485 24361 15519 24395
rect 15519 24361 15528 24395
rect 15476 24352 15528 24361
rect 16580 24395 16632 24404
rect 16580 24361 16589 24395
rect 16589 24361 16623 24395
rect 16623 24361 16632 24395
rect 16580 24352 16632 24361
rect 19248 24352 19300 24404
rect 19524 24395 19576 24404
rect 19524 24361 19533 24395
rect 19533 24361 19567 24395
rect 19567 24361 19576 24395
rect 19524 24352 19576 24361
rect 20076 24352 20128 24404
rect 20168 24352 20220 24404
rect 25504 24395 25556 24404
rect 25504 24361 25513 24395
rect 25513 24361 25547 24395
rect 25547 24361 25556 24395
rect 25504 24352 25556 24361
rect 9864 24284 9916 24336
rect 16396 24284 16448 24336
rect 16672 24284 16724 24336
rect 1768 24216 1820 24268
rect 3240 24216 3292 24268
rect 4620 24216 4672 24268
rect 5540 24216 5592 24268
rect 6276 24216 6328 24268
rect 12072 24259 12124 24268
rect 12072 24225 12081 24259
rect 12081 24225 12115 24259
rect 12115 24225 12124 24259
rect 12072 24216 12124 24225
rect 14096 24216 14148 24268
rect 15292 24216 15344 24268
rect 15660 24216 15712 24268
rect 18052 24216 18104 24268
rect 19340 24216 19392 24268
rect 21088 24216 21140 24268
rect 22836 24259 22888 24268
rect 22836 24225 22845 24259
rect 22845 24225 22879 24259
rect 22879 24225 22888 24259
rect 22836 24216 22888 24225
rect 23940 24216 23992 24268
rect 24860 24216 24912 24268
rect 25780 24216 25832 24268
rect 2780 24148 2832 24200
rect 4344 24148 4396 24200
rect 4804 24148 4856 24200
rect 6920 24080 6972 24132
rect 9496 24148 9548 24200
rect 11428 24148 11480 24200
rect 11060 24080 11112 24132
rect 12256 24191 12308 24200
rect 12256 24157 12265 24191
rect 12265 24157 12299 24191
rect 12299 24157 12308 24191
rect 12256 24148 12308 24157
rect 14188 24148 14240 24200
rect 14648 24148 14700 24200
rect 15936 24191 15988 24200
rect 15936 24157 15945 24191
rect 15945 24157 15979 24191
rect 15979 24157 15988 24191
rect 15936 24148 15988 24157
rect 14740 24080 14792 24132
rect 15844 24080 15896 24132
rect 17868 24148 17920 24200
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 18696 24191 18748 24200
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 20812 24148 20864 24200
rect 19248 24080 19300 24132
rect 19524 24080 19576 24132
rect 20352 24080 20404 24132
rect 21640 24080 21692 24132
rect 22284 24148 22336 24200
rect 23020 24191 23072 24200
rect 23020 24157 23029 24191
rect 23029 24157 23063 24191
rect 23063 24157 23072 24191
rect 23020 24148 23072 24157
rect 23480 24148 23532 24200
rect 1400 24012 1452 24064
rect 1768 24012 1820 24064
rect 2780 24012 2832 24064
rect 4896 24055 4948 24064
rect 4896 24021 4905 24055
rect 4905 24021 4939 24055
rect 4939 24021 4948 24055
rect 4896 24012 4948 24021
rect 5264 24055 5316 24064
rect 5264 24021 5273 24055
rect 5273 24021 5307 24055
rect 5307 24021 5316 24055
rect 5264 24012 5316 24021
rect 7012 24055 7064 24064
rect 7012 24021 7021 24055
rect 7021 24021 7055 24055
rect 7055 24021 7064 24055
rect 7012 24012 7064 24021
rect 7656 24012 7708 24064
rect 8116 24012 8168 24064
rect 8944 24055 8996 24064
rect 8944 24021 8953 24055
rect 8953 24021 8987 24055
rect 8987 24021 8996 24055
rect 8944 24012 8996 24021
rect 10692 24055 10744 24064
rect 10692 24021 10701 24055
rect 10701 24021 10735 24055
rect 10735 24021 10744 24055
rect 10692 24012 10744 24021
rect 12348 24012 12400 24064
rect 12992 24055 13044 24064
rect 12992 24021 13001 24055
rect 13001 24021 13035 24055
rect 13035 24021 13044 24055
rect 12992 24012 13044 24021
rect 13728 24012 13780 24064
rect 15476 24012 15528 24064
rect 18604 24012 18656 24064
rect 19156 24055 19208 24064
rect 19156 24021 19165 24055
rect 19165 24021 19199 24055
rect 19199 24021 19208 24055
rect 19156 24012 19208 24021
rect 20720 24012 20772 24064
rect 22376 24080 22428 24132
rect 23572 24012 23624 24064
rect 24124 24012 24176 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2136 23808 2188 23860
rect 2688 23808 2740 23860
rect 3240 23808 3292 23860
rect 3792 23851 3844 23860
rect 3792 23817 3801 23851
rect 3801 23817 3835 23851
rect 3835 23817 3844 23851
rect 3792 23808 3844 23817
rect 4620 23851 4672 23860
rect 4620 23817 4629 23851
rect 4629 23817 4663 23851
rect 4663 23817 4672 23851
rect 4620 23808 4672 23817
rect 5080 23808 5132 23860
rect 8300 23851 8352 23860
rect 8300 23817 8309 23851
rect 8309 23817 8343 23851
rect 8343 23817 8352 23851
rect 8300 23808 8352 23817
rect 8852 23808 8904 23860
rect 9772 23808 9824 23860
rect 11428 23851 11480 23860
rect 11428 23817 11437 23851
rect 11437 23817 11471 23851
rect 11471 23817 11480 23851
rect 11428 23808 11480 23817
rect 12256 23851 12308 23860
rect 12256 23817 12265 23851
rect 12265 23817 12299 23851
rect 12299 23817 12308 23851
rect 12256 23808 12308 23817
rect 15844 23808 15896 23860
rect 15936 23808 15988 23860
rect 18696 23808 18748 23860
rect 22376 23808 22428 23860
rect 5264 23672 5316 23724
rect 10876 23740 10928 23792
rect 2504 23647 2556 23656
rect 2504 23613 2513 23647
rect 2513 23613 2547 23647
rect 2547 23613 2556 23647
rect 2504 23604 2556 23613
rect 4528 23604 4580 23656
rect 4896 23604 4948 23656
rect 7012 23672 7064 23724
rect 7288 23715 7340 23724
rect 7288 23681 7297 23715
rect 7297 23681 7331 23715
rect 7331 23681 7340 23715
rect 7288 23672 7340 23681
rect 6552 23604 6604 23656
rect 8300 23672 8352 23724
rect 8944 23715 8996 23724
rect 8944 23681 8953 23715
rect 8953 23681 8987 23715
rect 8987 23681 8996 23715
rect 8944 23672 8996 23681
rect 9956 23672 10008 23724
rect 10692 23715 10744 23724
rect 10692 23681 10701 23715
rect 10701 23681 10735 23715
rect 10735 23681 10744 23715
rect 10692 23672 10744 23681
rect 14832 23672 14884 23724
rect 20352 23715 20404 23724
rect 20352 23681 20361 23715
rect 20361 23681 20395 23715
rect 20395 23681 20404 23715
rect 20352 23672 20404 23681
rect 24032 23808 24084 23860
rect 25596 23808 25648 23860
rect 25780 23851 25832 23860
rect 25780 23817 25789 23851
rect 25789 23817 25823 23851
rect 25823 23817 25832 23851
rect 25780 23808 25832 23817
rect 25228 23740 25280 23792
rect 10048 23604 10100 23656
rect 10140 23604 10192 23656
rect 10784 23604 10836 23656
rect 11336 23604 11388 23656
rect 19248 23604 19300 23656
rect 21916 23604 21968 23656
rect 8852 23579 8904 23588
rect 8852 23545 8861 23579
rect 8861 23545 8895 23579
rect 8895 23545 8904 23579
rect 8852 23536 8904 23545
rect 10600 23536 10652 23588
rect 12256 23536 12308 23588
rect 12716 23579 12768 23588
rect 12716 23545 12728 23579
rect 12728 23545 12768 23579
rect 15476 23579 15528 23588
rect 12716 23536 12768 23545
rect 15476 23545 15510 23579
rect 15510 23545 15528 23579
rect 15476 23536 15528 23545
rect 1676 23468 1728 23520
rect 1952 23511 2004 23520
rect 1952 23477 1961 23511
rect 1961 23477 1995 23511
rect 1995 23477 2004 23511
rect 1952 23468 2004 23477
rect 2688 23511 2740 23520
rect 2688 23477 2697 23511
rect 2697 23477 2731 23511
rect 2731 23477 2740 23511
rect 2688 23468 2740 23477
rect 3516 23511 3568 23520
rect 3516 23477 3525 23511
rect 3525 23477 3559 23511
rect 3559 23477 3568 23511
rect 3516 23468 3568 23477
rect 5172 23511 5224 23520
rect 5172 23477 5181 23511
rect 5181 23477 5215 23511
rect 5215 23477 5224 23511
rect 5172 23468 5224 23477
rect 6552 23511 6604 23520
rect 6552 23477 6561 23511
rect 6561 23477 6595 23511
rect 6595 23477 6604 23511
rect 6552 23468 6604 23477
rect 6920 23468 6972 23520
rect 9772 23468 9824 23520
rect 20536 23536 20588 23588
rect 22100 23536 22152 23588
rect 22652 23604 22704 23656
rect 22468 23536 22520 23588
rect 22836 23536 22888 23588
rect 10784 23468 10836 23520
rect 13820 23511 13872 23520
rect 13820 23477 13829 23511
rect 13829 23477 13863 23511
rect 13863 23477 13872 23511
rect 13820 23468 13872 23477
rect 14188 23511 14240 23520
rect 14188 23477 14197 23511
rect 14197 23477 14231 23511
rect 14231 23477 14240 23511
rect 14188 23468 14240 23477
rect 14740 23468 14792 23520
rect 15844 23468 15896 23520
rect 16580 23511 16632 23520
rect 16580 23477 16589 23511
rect 16589 23477 16623 23511
rect 16623 23477 16632 23511
rect 16580 23468 16632 23477
rect 17500 23511 17552 23520
rect 17500 23477 17509 23511
rect 17509 23477 17543 23511
rect 17543 23477 17552 23511
rect 17500 23468 17552 23477
rect 19340 23468 19392 23520
rect 20352 23468 20404 23520
rect 20812 23468 20864 23520
rect 21732 23511 21784 23520
rect 21732 23477 21741 23511
rect 21741 23477 21775 23511
rect 21775 23477 21784 23511
rect 21732 23468 21784 23477
rect 22284 23468 22336 23520
rect 22560 23511 22612 23520
rect 22560 23477 22569 23511
rect 22569 23477 22603 23511
rect 22603 23477 22612 23511
rect 22560 23468 22612 23477
rect 23388 23468 23440 23520
rect 24032 23511 24084 23520
rect 24032 23477 24041 23511
rect 24041 23477 24075 23511
rect 24075 23477 24084 23511
rect 24032 23468 24084 23477
rect 24124 23511 24176 23520
rect 24124 23477 24133 23511
rect 24133 23477 24167 23511
rect 24167 23477 24176 23511
rect 24124 23468 24176 23477
rect 24952 23468 25004 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 2596 23264 2648 23316
rect 4068 23264 4120 23316
rect 2228 23196 2280 23248
rect 3516 23239 3568 23248
rect 3516 23205 3525 23239
rect 3525 23205 3559 23239
rect 3559 23205 3568 23239
rect 3516 23196 3568 23205
rect 3976 23196 4028 23248
rect 5448 23264 5500 23316
rect 7288 23307 7340 23316
rect 7288 23273 7297 23307
rect 7297 23273 7331 23307
rect 7331 23273 7340 23307
rect 7288 23264 7340 23273
rect 9036 23307 9088 23316
rect 9036 23273 9045 23307
rect 9045 23273 9079 23307
rect 9079 23273 9088 23307
rect 9036 23264 9088 23273
rect 9588 23264 9640 23316
rect 9772 23264 9824 23316
rect 11244 23307 11296 23316
rect 11244 23273 11253 23307
rect 11253 23273 11287 23307
rect 11287 23273 11296 23307
rect 11244 23264 11296 23273
rect 12072 23264 12124 23316
rect 12716 23307 12768 23316
rect 12716 23273 12725 23307
rect 12725 23273 12759 23307
rect 12759 23273 12768 23307
rect 12716 23264 12768 23273
rect 13636 23264 13688 23316
rect 13728 23264 13780 23316
rect 15108 23307 15160 23316
rect 15108 23273 15117 23307
rect 15117 23273 15151 23307
rect 15151 23273 15160 23307
rect 15108 23264 15160 23273
rect 15476 23264 15528 23316
rect 16488 23264 16540 23316
rect 17500 23264 17552 23316
rect 18328 23264 18380 23316
rect 18512 23307 18564 23316
rect 18512 23273 18521 23307
rect 18521 23273 18555 23307
rect 18555 23273 18564 23307
rect 18512 23264 18564 23273
rect 20536 23264 20588 23316
rect 23020 23264 23072 23316
rect 23572 23307 23624 23316
rect 23572 23273 23581 23307
rect 23581 23273 23615 23307
rect 23615 23273 23624 23307
rect 23572 23264 23624 23273
rect 24860 23307 24912 23316
rect 24860 23273 24869 23307
rect 24869 23273 24903 23307
rect 24903 23273 24912 23307
rect 24860 23264 24912 23273
rect 25504 23307 25556 23316
rect 25504 23273 25513 23307
rect 25513 23273 25547 23307
rect 25547 23273 25556 23307
rect 25504 23264 25556 23273
rect 12440 23196 12492 23248
rect 16120 23196 16172 23248
rect 16580 23239 16632 23248
rect 16580 23205 16614 23239
rect 16614 23205 16632 23239
rect 16580 23196 16632 23205
rect 18696 23196 18748 23248
rect 21732 23196 21784 23248
rect 6184 23128 6236 23180
rect 7656 23171 7708 23180
rect 7656 23137 7690 23171
rect 7690 23137 7708 23171
rect 7656 23128 7708 23137
rect 10048 23171 10100 23180
rect 10048 23137 10057 23171
rect 10057 23137 10091 23171
rect 10091 23137 10100 23171
rect 10048 23128 10100 23137
rect 11612 23171 11664 23180
rect 11612 23137 11646 23171
rect 11646 23137 11664 23171
rect 11612 23128 11664 23137
rect 12624 23128 12676 23180
rect 15936 23128 15988 23180
rect 16396 23128 16448 23180
rect 19248 23128 19300 23180
rect 21640 23128 21692 23180
rect 23848 23128 23900 23180
rect 25320 23171 25372 23180
rect 25320 23137 25329 23171
rect 25329 23137 25363 23171
rect 25363 23137 25372 23171
rect 25320 23128 25372 23137
rect 4988 23060 5040 23112
rect 7380 23103 7432 23112
rect 7380 23069 7389 23103
rect 7389 23069 7423 23103
rect 7423 23069 7432 23103
rect 7380 23060 7432 23069
rect 9496 23060 9548 23112
rect 3884 22992 3936 23044
rect 9772 22992 9824 23044
rect 10600 23060 10652 23112
rect 10784 23060 10836 23112
rect 11336 23103 11388 23112
rect 11336 23069 11345 23103
rect 11345 23069 11379 23103
rect 11379 23069 11388 23103
rect 11336 23060 11388 23069
rect 12532 23060 12584 23112
rect 13636 23060 13688 23112
rect 14096 23103 14148 23112
rect 14096 23069 14105 23103
rect 14105 23069 14139 23103
rect 14139 23069 14148 23103
rect 15292 23103 15344 23112
rect 14096 23060 14148 23069
rect 15292 23069 15301 23103
rect 15301 23069 15335 23103
rect 15335 23069 15344 23103
rect 15292 23060 15344 23069
rect 23940 23060 23992 23112
rect 23480 22992 23532 23044
rect 5080 22967 5132 22976
rect 5080 22933 5089 22967
rect 5089 22933 5123 22967
rect 5123 22933 5132 22967
rect 5080 22924 5132 22933
rect 6552 22967 6604 22976
rect 6552 22933 6561 22967
rect 6561 22933 6595 22967
rect 6595 22933 6604 22967
rect 6552 22924 6604 22933
rect 7196 22924 7248 22976
rect 8392 22924 8444 22976
rect 10784 22967 10836 22976
rect 10784 22933 10793 22967
rect 10793 22933 10827 22967
rect 10827 22933 10836 22967
rect 10784 22924 10836 22933
rect 12808 22924 12860 22976
rect 14372 22924 14424 22976
rect 16672 22924 16724 22976
rect 21088 22967 21140 22976
rect 21088 22933 21097 22967
rect 21097 22933 21131 22967
rect 21131 22933 21140 22967
rect 21088 22924 21140 22933
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2228 22763 2280 22772
rect 2228 22729 2237 22763
rect 2237 22729 2271 22763
rect 2271 22729 2280 22763
rect 2228 22720 2280 22729
rect 4896 22720 4948 22772
rect 7012 22720 7064 22772
rect 4988 22695 5040 22704
rect 4988 22661 4997 22695
rect 4997 22661 5031 22695
rect 5031 22661 5040 22695
rect 4988 22652 5040 22661
rect 2596 22584 2648 22636
rect 2136 22516 2188 22568
rect 3976 22516 4028 22568
rect 5080 22584 5132 22636
rect 8944 22720 8996 22772
rect 9496 22763 9548 22772
rect 9496 22729 9505 22763
rect 9505 22729 9539 22763
rect 9539 22729 9548 22763
rect 9496 22720 9548 22729
rect 10968 22720 11020 22772
rect 12716 22720 12768 22772
rect 14096 22720 14148 22772
rect 15844 22763 15896 22772
rect 15844 22729 15853 22763
rect 15853 22729 15887 22763
rect 15887 22729 15896 22763
rect 15844 22720 15896 22729
rect 18052 22763 18104 22772
rect 18052 22729 18061 22763
rect 18061 22729 18095 22763
rect 18095 22729 18104 22763
rect 18052 22720 18104 22729
rect 18696 22720 18748 22772
rect 19984 22720 20036 22772
rect 20628 22720 20680 22772
rect 5816 22627 5868 22636
rect 5816 22593 5825 22627
rect 5825 22593 5859 22627
rect 5859 22593 5868 22627
rect 5816 22584 5868 22593
rect 6552 22584 6604 22636
rect 7472 22627 7524 22636
rect 7472 22593 7481 22627
rect 7481 22593 7515 22627
rect 7515 22593 7524 22627
rect 7472 22584 7524 22593
rect 8208 22584 8260 22636
rect 9036 22627 9088 22636
rect 9036 22593 9045 22627
rect 9045 22593 9079 22627
rect 9079 22593 9088 22627
rect 9036 22584 9088 22593
rect 9772 22652 9824 22704
rect 6184 22516 6236 22568
rect 10600 22516 10652 22568
rect 11612 22584 11664 22636
rect 4160 22448 4212 22500
rect 11336 22516 11388 22568
rect 12440 22584 12492 22636
rect 15660 22652 15712 22704
rect 16396 22652 16448 22704
rect 13820 22584 13872 22636
rect 12532 22516 12584 22568
rect 12808 22559 12860 22568
rect 12808 22525 12817 22559
rect 12817 22525 12851 22559
rect 12851 22525 12860 22559
rect 12808 22516 12860 22525
rect 14096 22559 14148 22568
rect 14096 22525 14105 22559
rect 14105 22525 14139 22559
rect 14139 22525 14148 22559
rect 14096 22516 14148 22525
rect 7288 22491 7340 22500
rect 4068 22423 4120 22432
rect 4068 22389 4077 22423
rect 4077 22389 4111 22423
rect 4111 22389 4120 22423
rect 4068 22380 4120 22389
rect 5356 22380 5408 22432
rect 7288 22457 7297 22491
rect 7297 22457 7331 22491
rect 7331 22457 7340 22491
rect 7288 22448 7340 22457
rect 10784 22448 10836 22500
rect 13452 22448 13504 22500
rect 13820 22448 13872 22500
rect 15384 22448 15436 22500
rect 7196 22423 7248 22432
rect 7196 22389 7205 22423
rect 7205 22389 7239 22423
rect 7239 22389 7248 22423
rect 7196 22380 7248 22389
rect 8392 22423 8444 22432
rect 8392 22389 8401 22423
rect 8401 22389 8435 22423
rect 8435 22389 8444 22423
rect 8392 22380 8444 22389
rect 12440 22423 12492 22432
rect 12440 22389 12449 22423
rect 12449 22389 12483 22423
rect 12483 22389 12492 22423
rect 12440 22380 12492 22389
rect 14740 22380 14792 22432
rect 15844 22380 15896 22432
rect 18328 22584 18380 22636
rect 18880 22584 18932 22636
rect 19248 22584 19300 22636
rect 21732 22720 21784 22772
rect 22008 22763 22060 22772
rect 22008 22729 22017 22763
rect 22017 22729 22051 22763
rect 22051 22729 22060 22763
rect 22008 22720 22060 22729
rect 22560 22720 22612 22772
rect 21824 22652 21876 22704
rect 19984 22516 20036 22568
rect 21088 22516 21140 22568
rect 21732 22516 21784 22568
rect 22192 22516 22244 22568
rect 22928 22584 22980 22636
rect 22560 22516 22612 22568
rect 25320 22720 25372 22772
rect 24308 22627 24360 22636
rect 24308 22593 24317 22627
rect 24317 22593 24351 22627
rect 24351 22593 24360 22627
rect 24308 22584 24360 22593
rect 17408 22491 17460 22500
rect 17408 22457 17417 22491
rect 17417 22457 17451 22491
rect 17451 22457 17460 22491
rect 17408 22448 17460 22457
rect 20904 22448 20956 22500
rect 16488 22380 16540 22432
rect 16672 22423 16724 22432
rect 16672 22389 16681 22423
rect 16681 22389 16715 22423
rect 16715 22389 16724 22423
rect 16672 22380 16724 22389
rect 18052 22380 18104 22432
rect 22652 22380 22704 22432
rect 23664 22380 23716 22432
rect 23940 22448 23992 22500
rect 25228 22448 25280 22500
rect 24952 22380 25004 22432
rect 25136 22423 25188 22432
rect 25136 22389 25145 22423
rect 25145 22389 25179 22423
rect 25179 22389 25188 22423
rect 25136 22380 25188 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2780 22219 2832 22228
rect 2780 22185 2789 22219
rect 2789 22185 2823 22219
rect 2823 22185 2832 22219
rect 2780 22176 2832 22185
rect 5816 22219 5868 22228
rect 4068 22108 4120 22160
rect 5816 22185 5825 22219
rect 5825 22185 5859 22219
rect 5859 22185 5868 22219
rect 5816 22176 5868 22185
rect 7104 22176 7156 22228
rect 7656 22219 7708 22228
rect 7656 22185 7665 22219
rect 7665 22185 7699 22219
rect 7699 22185 7708 22219
rect 7656 22176 7708 22185
rect 10784 22176 10836 22228
rect 11796 22176 11848 22228
rect 13268 22176 13320 22228
rect 6184 22108 6236 22160
rect 11336 22151 11388 22160
rect 11336 22117 11370 22151
rect 11370 22117 11388 22151
rect 11336 22108 11388 22117
rect 12900 22108 12952 22160
rect 13084 22108 13136 22160
rect 13820 22176 13872 22228
rect 18052 22219 18104 22228
rect 18052 22185 18061 22219
rect 18061 22185 18095 22219
rect 18095 22185 18104 22219
rect 18052 22176 18104 22185
rect 18328 22176 18380 22228
rect 9128 22040 9180 22092
rect 9588 22040 9640 22092
rect 10968 22040 11020 22092
rect 11612 22040 11664 22092
rect 13544 22108 13596 22160
rect 18512 22176 18564 22228
rect 20076 22176 20128 22228
rect 20904 22219 20956 22228
rect 2596 21972 2648 22024
rect 3516 21972 3568 22024
rect 3976 21972 4028 22024
rect 6736 21972 6788 22024
rect 7472 21972 7524 22024
rect 9496 21972 9548 22024
rect 12624 21972 12676 22024
rect 6092 21947 6144 21956
rect 6092 21913 6101 21947
rect 6101 21913 6135 21947
rect 6135 21913 6144 21947
rect 6092 21904 6144 21913
rect 6828 21904 6880 21956
rect 9036 21947 9088 21956
rect 9036 21913 9045 21947
rect 9045 21913 9079 21947
rect 9079 21913 9088 21947
rect 9036 21904 9088 21913
rect 13176 21972 13228 22024
rect 13912 22015 13964 22024
rect 13912 21981 13921 22015
rect 13921 21981 13955 22015
rect 13955 21981 13964 22015
rect 13912 21972 13964 21981
rect 14004 21972 14056 22024
rect 1492 21836 1544 21888
rect 2412 21879 2464 21888
rect 2412 21845 2421 21879
rect 2421 21845 2455 21879
rect 2455 21845 2464 21879
rect 2412 21836 2464 21845
rect 3424 21879 3476 21888
rect 3424 21845 3433 21879
rect 3433 21845 3467 21879
rect 3467 21845 3476 21879
rect 3424 21836 3476 21845
rect 3792 21879 3844 21888
rect 3792 21845 3801 21879
rect 3801 21845 3835 21879
rect 3835 21845 3844 21879
rect 3792 21836 3844 21845
rect 6276 21836 6328 21888
rect 7380 21836 7432 21888
rect 9772 21836 9824 21888
rect 10048 21836 10100 21888
rect 10968 21836 11020 21888
rect 12992 21836 13044 21888
rect 13912 21836 13964 21888
rect 14372 22040 14424 22092
rect 14280 21904 14332 21956
rect 14832 21904 14884 21956
rect 14740 21836 14792 21888
rect 17040 22040 17092 22092
rect 18972 22083 19024 22092
rect 18972 22049 18981 22083
rect 18981 22049 19015 22083
rect 19015 22049 19024 22083
rect 18972 22040 19024 22049
rect 20536 22108 20588 22160
rect 20904 22185 20913 22219
rect 20913 22185 20947 22219
rect 20947 22185 20956 22219
rect 20904 22176 20956 22185
rect 21272 22219 21324 22228
rect 21272 22185 21281 22219
rect 21281 22185 21315 22219
rect 21315 22185 21324 22219
rect 21272 22176 21324 22185
rect 22192 22176 22244 22228
rect 23848 22176 23900 22228
rect 23940 22176 23992 22228
rect 21640 22108 21692 22160
rect 15660 21972 15712 22024
rect 15936 21972 15988 22024
rect 17776 21972 17828 22024
rect 21364 22015 21416 22024
rect 21364 21981 21373 22015
rect 21373 21981 21407 22015
rect 21407 21981 21416 22015
rect 21364 21972 21416 21981
rect 21548 22040 21600 22092
rect 21824 22040 21876 22092
rect 22928 22108 22980 22160
rect 22744 22083 22796 22092
rect 22744 22049 22753 22083
rect 22753 22049 22787 22083
rect 22787 22049 22796 22083
rect 22744 22040 22796 22049
rect 24308 22040 24360 22092
rect 22192 21972 22244 22024
rect 24400 21972 24452 22024
rect 16304 21904 16356 21956
rect 20536 21904 20588 21956
rect 21916 21904 21968 21956
rect 15936 21836 15988 21888
rect 16580 21836 16632 21888
rect 19984 21879 20036 21888
rect 19984 21845 19993 21879
rect 19993 21845 20027 21879
rect 20027 21845 20036 21879
rect 19984 21836 20036 21845
rect 21548 21836 21600 21888
rect 23848 21836 23900 21888
rect 26148 21972 26200 22024
rect 24860 21904 24912 21956
rect 24952 21836 25004 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 2504 21675 2556 21684
rect 2504 21641 2513 21675
rect 2513 21641 2547 21675
rect 2547 21641 2556 21675
rect 2504 21632 2556 21641
rect 4160 21675 4212 21684
rect 4160 21641 4169 21675
rect 4169 21641 4203 21675
rect 4203 21641 4212 21675
rect 4160 21632 4212 21641
rect 4620 21632 4672 21684
rect 6184 21675 6236 21684
rect 4068 21564 4120 21616
rect 6184 21641 6193 21675
rect 6193 21641 6227 21675
rect 6227 21641 6236 21675
rect 6184 21632 6236 21641
rect 8760 21675 8812 21684
rect 8760 21641 8769 21675
rect 8769 21641 8803 21675
rect 8803 21641 8812 21675
rect 8760 21632 8812 21641
rect 9128 21675 9180 21684
rect 9128 21641 9137 21675
rect 9137 21641 9171 21675
rect 9171 21641 9180 21675
rect 9128 21632 9180 21641
rect 9680 21632 9732 21684
rect 11336 21675 11388 21684
rect 11336 21641 11345 21675
rect 11345 21641 11379 21675
rect 11379 21641 11388 21675
rect 11336 21632 11388 21641
rect 12348 21632 12400 21684
rect 14832 21632 14884 21684
rect 15936 21632 15988 21684
rect 16304 21632 16356 21684
rect 19340 21632 19392 21684
rect 21180 21675 21232 21684
rect 21180 21641 21189 21675
rect 21189 21641 21223 21675
rect 21223 21641 21232 21675
rect 21180 21632 21232 21641
rect 22192 21675 22244 21684
rect 22192 21641 22201 21675
rect 22201 21641 22235 21675
rect 22235 21641 22244 21675
rect 22192 21632 22244 21641
rect 22928 21632 22980 21684
rect 1768 21539 1820 21548
rect 1768 21505 1777 21539
rect 1777 21505 1811 21539
rect 1811 21505 1820 21539
rect 1768 21496 1820 21505
rect 5448 21539 5500 21548
rect 5448 21505 5457 21539
rect 5457 21505 5491 21539
rect 5491 21505 5500 21539
rect 5448 21496 5500 21505
rect 9128 21496 9180 21548
rect 9404 21496 9456 21548
rect 10048 21496 10100 21548
rect 12348 21496 12400 21548
rect 13728 21496 13780 21548
rect 1492 21471 1544 21480
rect 1492 21437 1501 21471
rect 1501 21437 1535 21471
rect 1535 21437 1544 21471
rect 1492 21428 1544 21437
rect 3976 21428 4028 21480
rect 5264 21428 5316 21480
rect 7380 21471 7432 21480
rect 7380 21437 7389 21471
rect 7389 21437 7423 21471
rect 7423 21437 7432 21471
rect 7380 21428 7432 21437
rect 7656 21471 7708 21480
rect 7656 21437 7690 21471
rect 7690 21437 7708 21471
rect 7656 21428 7708 21437
rect 8208 21428 8260 21480
rect 11060 21428 11112 21480
rect 12164 21428 12216 21480
rect 3516 21360 3568 21412
rect 14648 21428 14700 21480
rect 15844 21564 15896 21616
rect 17776 21607 17828 21616
rect 17776 21573 17785 21607
rect 17785 21573 17819 21607
rect 17819 21573 17828 21607
rect 17776 21564 17828 21573
rect 18512 21564 18564 21616
rect 18972 21564 19024 21616
rect 16672 21428 16724 21480
rect 20536 21496 20588 21548
rect 21732 21539 21784 21548
rect 21732 21505 21741 21539
rect 21741 21505 21775 21539
rect 21775 21505 21784 21539
rect 21732 21496 21784 21505
rect 22468 21496 22520 21548
rect 22836 21496 22888 21548
rect 19432 21428 19484 21480
rect 22744 21428 22796 21480
rect 23940 21471 23992 21480
rect 23940 21437 23974 21471
rect 23974 21437 23992 21471
rect 23940 21428 23992 21437
rect 14280 21360 14332 21412
rect 15292 21360 15344 21412
rect 15476 21360 15528 21412
rect 2872 21292 2924 21344
rect 6644 21335 6696 21344
rect 6644 21301 6653 21335
rect 6653 21301 6687 21335
rect 6687 21301 6696 21335
rect 6644 21292 6696 21301
rect 7104 21335 7156 21344
rect 7104 21301 7113 21335
rect 7113 21301 7147 21335
rect 7147 21301 7156 21335
rect 7104 21292 7156 21301
rect 9680 21335 9732 21344
rect 9680 21301 9689 21335
rect 9689 21301 9723 21335
rect 9723 21301 9732 21335
rect 9680 21292 9732 21301
rect 10048 21335 10100 21344
rect 10048 21301 10057 21335
rect 10057 21301 10091 21335
rect 10091 21301 10100 21335
rect 10048 21292 10100 21301
rect 10968 21292 11020 21344
rect 13176 21292 13228 21344
rect 14004 21292 14056 21344
rect 14096 21292 14148 21344
rect 15844 21292 15896 21344
rect 17592 21360 17644 21412
rect 20720 21360 20772 21412
rect 24860 21360 24912 21412
rect 16120 21335 16172 21344
rect 16120 21301 16129 21335
rect 16129 21301 16163 21335
rect 16163 21301 16172 21335
rect 16120 21292 16172 21301
rect 16304 21292 16356 21344
rect 16948 21292 17000 21344
rect 18420 21335 18472 21344
rect 18420 21301 18429 21335
rect 18429 21301 18463 21335
rect 18463 21301 18472 21335
rect 18420 21292 18472 21301
rect 19064 21292 19116 21344
rect 21364 21292 21416 21344
rect 21548 21335 21600 21344
rect 21548 21301 21557 21335
rect 21557 21301 21591 21335
rect 21591 21301 21600 21335
rect 21548 21292 21600 21301
rect 24952 21292 25004 21344
rect 25688 21335 25740 21344
rect 25688 21301 25697 21335
rect 25697 21301 25731 21335
rect 25731 21301 25740 21335
rect 25688 21292 25740 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1492 21088 1544 21140
rect 5448 21088 5500 21140
rect 6276 21088 6328 21140
rect 7656 21088 7708 21140
rect 8024 21131 8076 21140
rect 8024 21097 8033 21131
rect 8033 21097 8067 21131
rect 8067 21097 8076 21131
rect 8024 21088 8076 21097
rect 8300 21088 8352 21140
rect 8576 21088 8628 21140
rect 11244 21088 11296 21140
rect 12624 21088 12676 21140
rect 13452 21131 13504 21140
rect 13452 21097 13461 21131
rect 13461 21097 13495 21131
rect 13495 21097 13504 21131
rect 13452 21088 13504 21097
rect 16120 21088 16172 21140
rect 18420 21088 18472 21140
rect 19340 21088 19392 21140
rect 20076 21088 20128 21140
rect 20720 21131 20772 21140
rect 20720 21097 20729 21131
rect 20729 21097 20763 21131
rect 20763 21097 20772 21131
rect 20720 21088 20772 21097
rect 21272 21088 21324 21140
rect 2872 21063 2924 21072
rect 2872 21029 2881 21063
rect 2881 21029 2915 21063
rect 2915 21029 2924 21063
rect 2872 21020 2924 21029
rect 3608 21020 3660 21072
rect 4160 21020 4212 21072
rect 8116 21020 8168 21072
rect 2596 20952 2648 21004
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 2872 20884 2924 20936
rect 4068 20884 4120 20936
rect 2504 20816 2556 20868
rect 5264 20952 5316 21004
rect 6092 20952 6144 21004
rect 6552 20952 6604 21004
rect 8300 20952 8352 21004
rect 9772 20952 9824 21004
rect 11612 21020 11664 21072
rect 12164 21063 12216 21072
rect 12164 21029 12173 21063
rect 12173 21029 12207 21063
rect 12207 21029 12216 21063
rect 12164 21020 12216 21029
rect 13820 21020 13872 21072
rect 16948 21020 17000 21072
rect 17592 21063 17644 21072
rect 17592 21029 17601 21063
rect 17601 21029 17635 21063
rect 17635 21029 17644 21063
rect 17592 21020 17644 21029
rect 19156 21020 19208 21072
rect 20812 21020 20864 21072
rect 21732 21088 21784 21140
rect 22008 21088 22060 21140
rect 22744 21088 22796 21140
rect 23940 21088 23992 21140
rect 10324 20995 10376 21004
rect 4620 20927 4672 20936
rect 4620 20893 4629 20927
rect 4629 20893 4663 20927
rect 4663 20893 4672 20927
rect 4620 20884 4672 20893
rect 6920 20927 6972 20936
rect 6920 20893 6929 20927
rect 6929 20893 6963 20927
rect 6963 20893 6972 20927
rect 6920 20884 6972 20893
rect 6736 20816 6788 20868
rect 7564 20884 7616 20936
rect 8668 20927 8720 20936
rect 8668 20893 8677 20927
rect 8677 20893 8711 20927
rect 8711 20893 8720 20927
rect 10324 20961 10358 20995
rect 10358 20961 10376 20995
rect 10324 20952 10376 20961
rect 13360 20952 13412 21004
rect 8668 20884 8720 20893
rect 13452 20884 13504 20936
rect 13820 20884 13872 20936
rect 14280 20884 14332 20936
rect 3516 20748 3568 20800
rect 6092 20791 6144 20800
rect 6092 20757 6101 20791
rect 6101 20757 6135 20791
rect 6135 20757 6144 20791
rect 6092 20748 6144 20757
rect 6920 20748 6972 20800
rect 9404 20748 9456 20800
rect 9680 20748 9732 20800
rect 10048 20748 10100 20800
rect 12348 20748 12400 20800
rect 13912 20748 13964 20800
rect 17040 20952 17092 21004
rect 20168 20995 20220 21004
rect 15476 20884 15528 20936
rect 16120 20884 16172 20936
rect 15844 20816 15896 20868
rect 14832 20748 14884 20800
rect 20168 20961 20177 20995
rect 20177 20961 20211 20995
rect 20211 20961 20220 20995
rect 20168 20952 20220 20961
rect 24952 20952 25004 21004
rect 22192 20884 22244 20936
rect 23020 20884 23072 20936
rect 17960 20748 18012 20800
rect 19432 20748 19484 20800
rect 21824 20791 21876 20800
rect 21824 20757 21833 20791
rect 21833 20757 21867 20791
rect 21867 20757 21876 20791
rect 21824 20748 21876 20757
rect 25044 20791 25096 20800
rect 25044 20757 25053 20791
rect 25053 20757 25087 20791
rect 25087 20757 25096 20791
rect 25044 20748 25096 20757
rect 25688 20748 25740 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2504 20587 2556 20596
rect 2504 20553 2513 20587
rect 2513 20553 2547 20587
rect 2547 20553 2556 20587
rect 2504 20544 2556 20553
rect 4068 20544 4120 20596
rect 6000 20544 6052 20596
rect 6552 20587 6604 20596
rect 6552 20553 6561 20587
rect 6561 20553 6595 20587
rect 6595 20553 6604 20587
rect 6552 20544 6604 20553
rect 7012 20544 7064 20596
rect 7564 20587 7616 20596
rect 7564 20553 7573 20587
rect 7573 20553 7607 20587
rect 7607 20553 7616 20587
rect 7564 20544 7616 20553
rect 10784 20544 10836 20596
rect 11796 20544 11848 20596
rect 13820 20587 13872 20596
rect 13820 20553 13829 20587
rect 13829 20553 13863 20587
rect 13863 20553 13872 20587
rect 13820 20544 13872 20553
rect 14832 20544 14884 20596
rect 12808 20476 12860 20528
rect 15384 20476 15436 20528
rect 3148 20451 3200 20460
rect 3148 20417 3157 20451
rect 3157 20417 3191 20451
rect 3191 20417 3200 20451
rect 3148 20408 3200 20417
rect 3608 20408 3660 20460
rect 3976 20408 4028 20460
rect 4528 20451 4580 20460
rect 4528 20417 4537 20451
rect 4537 20417 4571 20451
rect 4571 20417 4580 20451
rect 4528 20408 4580 20417
rect 9772 20408 9824 20460
rect 11704 20408 11756 20460
rect 12992 20451 13044 20460
rect 2412 20383 2464 20392
rect 2412 20349 2421 20383
rect 2421 20349 2455 20383
rect 2455 20349 2464 20383
rect 2412 20340 2464 20349
rect 7380 20340 7432 20392
rect 9404 20340 9456 20392
rect 11980 20340 12032 20392
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 2044 20247 2096 20256
rect 2044 20213 2053 20247
rect 2053 20213 2087 20247
rect 2087 20213 2096 20247
rect 2044 20204 2096 20213
rect 2872 20247 2924 20256
rect 2872 20213 2881 20247
rect 2881 20213 2915 20247
rect 2915 20213 2924 20247
rect 2872 20204 2924 20213
rect 3608 20204 3660 20256
rect 5540 20272 5592 20324
rect 8116 20272 8168 20324
rect 10048 20272 10100 20324
rect 10324 20272 10376 20324
rect 11612 20272 11664 20324
rect 12992 20417 13001 20451
rect 13001 20417 13035 20451
rect 13035 20417 13044 20451
rect 12992 20408 13044 20417
rect 17960 20408 18012 20460
rect 19248 20544 19300 20596
rect 24768 20544 24820 20596
rect 20076 20408 20128 20460
rect 24124 20451 24176 20460
rect 24124 20417 24133 20451
rect 24133 20417 24167 20451
rect 24167 20417 24176 20451
rect 24124 20408 24176 20417
rect 24308 20451 24360 20460
rect 24308 20417 24317 20451
rect 24317 20417 24351 20451
rect 24351 20417 24360 20451
rect 24308 20408 24360 20417
rect 25136 20408 25188 20460
rect 12348 20340 12400 20392
rect 12808 20383 12860 20392
rect 12808 20349 12817 20383
rect 12817 20349 12851 20383
rect 12851 20349 12860 20383
rect 12808 20340 12860 20349
rect 14096 20383 14148 20392
rect 14096 20349 14105 20383
rect 14105 20349 14139 20383
rect 14139 20349 14148 20383
rect 14096 20340 14148 20349
rect 14648 20340 14700 20392
rect 16580 20340 16632 20392
rect 20628 20340 20680 20392
rect 8024 20204 8076 20256
rect 8852 20204 8904 20256
rect 9404 20247 9456 20256
rect 9404 20213 9413 20247
rect 9413 20213 9447 20247
rect 9447 20213 9456 20247
rect 9404 20204 9456 20213
rect 13820 20272 13872 20324
rect 15384 20272 15436 20324
rect 15660 20272 15712 20324
rect 16948 20272 17000 20324
rect 19156 20272 19208 20324
rect 23388 20340 23440 20392
rect 23664 20340 23716 20392
rect 23756 20340 23808 20392
rect 25320 20340 25372 20392
rect 25136 20272 25188 20324
rect 26240 20272 26292 20324
rect 12164 20204 12216 20256
rect 12440 20247 12492 20256
rect 12440 20213 12449 20247
rect 12449 20213 12483 20247
rect 12483 20213 12492 20247
rect 13452 20247 13504 20256
rect 12440 20204 12492 20213
rect 13452 20213 13461 20247
rect 13461 20213 13495 20247
rect 13495 20213 13504 20247
rect 13452 20204 13504 20213
rect 16120 20204 16172 20256
rect 18052 20247 18104 20256
rect 18052 20213 18061 20247
rect 18061 20213 18095 20247
rect 18095 20213 18104 20247
rect 18052 20204 18104 20213
rect 18420 20204 18472 20256
rect 20444 20247 20496 20256
rect 20444 20213 20453 20247
rect 20453 20213 20487 20247
rect 20487 20213 20496 20247
rect 20444 20204 20496 20213
rect 21088 20247 21140 20256
rect 21088 20213 21097 20247
rect 21097 20213 21131 20247
rect 21131 20213 21140 20247
rect 21088 20204 21140 20213
rect 21824 20204 21876 20256
rect 22192 20204 22244 20256
rect 22376 20204 22428 20256
rect 22652 20247 22704 20256
rect 22652 20213 22661 20247
rect 22661 20213 22695 20247
rect 22695 20213 22704 20247
rect 22652 20204 22704 20213
rect 23020 20247 23072 20256
rect 23020 20213 23029 20247
rect 23029 20213 23063 20247
rect 23063 20213 23072 20247
rect 23020 20204 23072 20213
rect 23572 20204 23624 20256
rect 23940 20204 23992 20256
rect 24308 20204 24360 20256
rect 25044 20247 25096 20256
rect 25044 20213 25053 20247
rect 25053 20213 25087 20247
rect 25087 20213 25096 20247
rect 25044 20204 25096 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2872 20000 2924 20052
rect 3516 20043 3568 20052
rect 3516 20009 3525 20043
rect 3525 20009 3559 20043
rect 3559 20009 3568 20043
rect 3516 20000 3568 20009
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 2872 19839 2924 19848
rect 2872 19805 2881 19839
rect 2881 19805 2915 19839
rect 2915 19805 2924 19839
rect 2872 19796 2924 19805
rect 3148 19932 3200 19984
rect 4068 20000 4120 20052
rect 4620 20000 4672 20052
rect 4436 19932 4488 19984
rect 6736 20000 6788 20052
rect 6920 20000 6972 20052
rect 7840 20000 7892 20052
rect 8208 20000 8260 20052
rect 8668 20000 8720 20052
rect 10140 20000 10192 20052
rect 10784 20043 10836 20052
rect 10784 20009 10793 20043
rect 10793 20009 10827 20043
rect 10827 20009 10836 20043
rect 10784 20000 10836 20009
rect 11060 20000 11112 20052
rect 12256 20000 12308 20052
rect 12624 20000 12676 20052
rect 13728 20000 13780 20052
rect 14648 20000 14700 20052
rect 16672 20043 16724 20052
rect 16672 20009 16681 20043
rect 16681 20009 16715 20043
rect 16715 20009 16724 20043
rect 16672 20000 16724 20009
rect 17776 20000 17828 20052
rect 18236 20000 18288 20052
rect 19524 20000 19576 20052
rect 21088 20000 21140 20052
rect 21824 20000 21876 20052
rect 23020 20000 23072 20052
rect 23756 20000 23808 20052
rect 24860 20043 24912 20052
rect 24860 20009 24869 20043
rect 24869 20009 24903 20043
rect 24903 20009 24912 20043
rect 24860 20000 24912 20009
rect 13360 19932 13412 19984
rect 16304 19932 16356 19984
rect 18420 19932 18472 19984
rect 20168 19932 20220 19984
rect 22008 19975 22060 19984
rect 22008 19941 22017 19975
rect 22017 19941 22051 19975
rect 22051 19941 22060 19975
rect 22008 19932 22060 19941
rect 24768 19932 24820 19984
rect 25044 19932 25096 19984
rect 4528 19864 4580 19916
rect 7288 19907 7340 19916
rect 7288 19873 7297 19907
rect 7297 19873 7331 19907
rect 7331 19873 7340 19907
rect 7288 19864 7340 19873
rect 9864 19864 9916 19916
rect 10968 19864 11020 19916
rect 12256 19907 12308 19916
rect 12256 19873 12265 19907
rect 12265 19873 12299 19907
rect 12299 19873 12308 19907
rect 12256 19864 12308 19873
rect 14096 19864 14148 19916
rect 15384 19864 15436 19916
rect 15844 19864 15896 19916
rect 17868 19864 17920 19916
rect 19524 19864 19576 19916
rect 21272 19907 21324 19916
rect 21272 19873 21281 19907
rect 21281 19873 21315 19907
rect 21315 19873 21324 19907
rect 21272 19864 21324 19873
rect 22376 19864 22428 19916
rect 22744 19864 22796 19916
rect 22928 19907 22980 19916
rect 22928 19873 22962 19907
rect 22962 19873 22980 19907
rect 22928 19864 22980 19873
rect 25688 19864 25740 19916
rect 6276 19796 6328 19848
rect 8576 19839 8628 19848
rect 8576 19805 8585 19839
rect 8585 19805 8619 19839
rect 8619 19805 8628 19839
rect 8576 19796 8628 19805
rect 10048 19796 10100 19848
rect 11980 19796 12032 19848
rect 12992 19796 13044 19848
rect 14004 19839 14056 19848
rect 14004 19805 14013 19839
rect 14013 19805 14047 19839
rect 14047 19805 14056 19839
rect 14004 19796 14056 19805
rect 6920 19771 6972 19780
rect 6920 19737 6929 19771
rect 6929 19737 6963 19771
rect 6963 19737 6972 19771
rect 6920 19728 6972 19737
rect 16764 19728 16816 19780
rect 19340 19796 19392 19848
rect 1860 19703 1912 19712
rect 1860 19669 1869 19703
rect 1869 19669 1903 19703
rect 1903 19669 1912 19703
rect 1860 19660 1912 19669
rect 2872 19660 2924 19712
rect 3700 19660 3752 19712
rect 7196 19660 7248 19712
rect 8944 19660 8996 19712
rect 9404 19660 9456 19712
rect 11428 19703 11480 19712
rect 11428 19669 11437 19703
rect 11437 19669 11471 19703
rect 11471 19669 11480 19703
rect 11428 19660 11480 19669
rect 14648 19660 14700 19712
rect 15476 19660 15528 19712
rect 17776 19660 17828 19712
rect 20536 19796 20588 19848
rect 20904 19796 20956 19848
rect 25320 19839 25372 19848
rect 25320 19805 25329 19839
rect 25329 19805 25363 19839
rect 25363 19805 25372 19839
rect 25320 19796 25372 19805
rect 25596 19796 25648 19848
rect 19984 19728 20036 19780
rect 23664 19728 23716 19780
rect 18328 19660 18380 19712
rect 19248 19703 19300 19712
rect 19248 19669 19257 19703
rect 19257 19669 19291 19703
rect 19291 19669 19300 19703
rect 19248 19660 19300 19669
rect 20444 19660 20496 19712
rect 21916 19660 21968 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2780 19499 2832 19508
rect 2780 19465 2789 19499
rect 2789 19465 2823 19499
rect 2823 19465 2832 19499
rect 2780 19456 2832 19465
rect 3976 19456 4028 19508
rect 4436 19499 4488 19508
rect 4436 19465 4445 19499
rect 4445 19465 4479 19499
rect 4479 19465 4488 19499
rect 4436 19456 4488 19465
rect 6828 19499 6880 19508
rect 6828 19465 6837 19499
rect 6837 19465 6871 19499
rect 6871 19465 6880 19499
rect 6828 19456 6880 19465
rect 7288 19456 7340 19508
rect 9128 19456 9180 19508
rect 10048 19456 10100 19508
rect 12256 19456 12308 19508
rect 2872 19388 2924 19440
rect 3148 19388 3200 19440
rect 9312 19388 9364 19440
rect 12164 19388 12216 19440
rect 1860 19320 1912 19372
rect 3516 19363 3568 19372
rect 3516 19329 3525 19363
rect 3525 19329 3559 19363
rect 3559 19329 3568 19363
rect 3516 19320 3568 19329
rect 4528 19363 4580 19372
rect 4528 19329 4537 19363
rect 4537 19329 4571 19363
rect 4571 19329 4580 19363
rect 4528 19320 4580 19329
rect 6736 19320 6788 19372
rect 7472 19320 7524 19372
rect 9128 19363 9180 19372
rect 9128 19329 9137 19363
rect 9137 19329 9171 19363
rect 9171 19329 9180 19363
rect 9128 19320 9180 19329
rect 9680 19320 9732 19372
rect 2228 19252 2280 19304
rect 3792 19252 3844 19304
rect 8668 19252 8720 19304
rect 9956 19295 10008 19304
rect 9956 19261 9965 19295
rect 9965 19261 9999 19295
rect 9999 19261 10008 19295
rect 9956 19252 10008 19261
rect 11336 19252 11388 19304
rect 12532 19252 12584 19304
rect 13084 19252 13136 19304
rect 13360 19295 13412 19304
rect 13360 19261 13369 19295
rect 13369 19261 13403 19295
rect 13403 19261 13412 19295
rect 13360 19252 13412 19261
rect 13820 19456 13872 19508
rect 17592 19499 17644 19508
rect 17592 19465 17601 19499
rect 17601 19465 17635 19499
rect 17635 19465 17644 19499
rect 17592 19456 17644 19465
rect 17868 19456 17920 19508
rect 19340 19456 19392 19508
rect 20628 19456 20680 19508
rect 21272 19456 21324 19508
rect 22928 19456 22980 19508
rect 17500 19388 17552 19440
rect 17960 19388 18012 19440
rect 16948 19363 17000 19372
rect 16948 19329 16957 19363
rect 16957 19329 16991 19363
rect 16991 19329 17000 19363
rect 16948 19320 17000 19329
rect 21088 19320 21140 19372
rect 21916 19363 21968 19372
rect 21916 19329 21925 19363
rect 21925 19329 21959 19363
rect 21959 19329 21968 19363
rect 21916 19320 21968 19329
rect 2872 19184 2924 19236
rect 3424 19227 3476 19236
rect 3424 19193 3433 19227
rect 3433 19193 3467 19227
rect 3467 19193 3476 19227
rect 3424 19184 3476 19193
rect 4804 19227 4856 19236
rect 4804 19193 4838 19227
rect 4838 19193 4856 19227
rect 4804 19184 4856 19193
rect 1676 19116 1728 19168
rect 2964 19159 3016 19168
rect 2964 19125 2973 19159
rect 2973 19125 3007 19159
rect 3007 19125 3016 19159
rect 2964 19116 3016 19125
rect 5540 19116 5592 19168
rect 6000 19116 6052 19168
rect 7196 19159 7248 19168
rect 7196 19125 7205 19159
rect 7205 19125 7239 19159
rect 7239 19125 7248 19159
rect 7196 19116 7248 19125
rect 7288 19159 7340 19168
rect 7288 19125 7297 19159
rect 7297 19125 7331 19159
rect 7331 19125 7340 19159
rect 8576 19159 8628 19168
rect 7288 19116 7340 19125
rect 8576 19125 8585 19159
rect 8585 19125 8619 19159
rect 8619 19125 8628 19159
rect 8576 19116 8628 19125
rect 8668 19116 8720 19168
rect 9864 19184 9916 19236
rect 13820 19227 13872 19236
rect 13820 19193 13854 19227
rect 13854 19193 13872 19227
rect 13820 19184 13872 19193
rect 9220 19116 9272 19168
rect 10140 19159 10192 19168
rect 10140 19125 10149 19159
rect 10149 19125 10183 19159
rect 10183 19125 10192 19159
rect 10140 19116 10192 19125
rect 10968 19116 11020 19168
rect 11244 19159 11296 19168
rect 11244 19125 11253 19159
rect 11253 19125 11287 19159
rect 11287 19125 11296 19159
rect 11244 19116 11296 19125
rect 12900 19116 12952 19168
rect 13084 19159 13136 19168
rect 13084 19125 13093 19159
rect 13093 19125 13127 19159
rect 13127 19125 13136 19159
rect 13084 19116 13136 19125
rect 15844 19252 15896 19304
rect 16304 19252 16356 19304
rect 16764 19295 16816 19304
rect 16764 19261 16773 19295
rect 16773 19261 16807 19295
rect 16807 19261 16816 19295
rect 16764 19252 16816 19261
rect 18328 19252 18380 19304
rect 18972 19252 19024 19304
rect 19892 19252 19944 19304
rect 20536 19252 20588 19304
rect 21732 19295 21784 19304
rect 21732 19261 21741 19295
rect 21741 19261 21775 19295
rect 21775 19261 21784 19295
rect 21732 19252 21784 19261
rect 24768 19252 24820 19304
rect 18144 19184 18196 19236
rect 19064 19184 19116 19236
rect 20076 19184 20128 19236
rect 15476 19116 15528 19168
rect 15660 19116 15712 19168
rect 16396 19159 16448 19168
rect 16396 19125 16405 19159
rect 16405 19125 16439 19159
rect 16439 19125 16448 19159
rect 16396 19116 16448 19125
rect 16856 19159 16908 19168
rect 16856 19125 16865 19159
rect 16865 19125 16899 19159
rect 16899 19125 16908 19159
rect 16856 19116 16908 19125
rect 17960 19116 18012 19168
rect 20720 19116 20772 19168
rect 25320 19184 25372 19236
rect 25780 19184 25832 19236
rect 21364 19159 21416 19168
rect 21364 19125 21373 19159
rect 21373 19125 21407 19159
rect 21407 19125 21416 19159
rect 21364 19116 21416 19125
rect 22376 19159 22428 19168
rect 22376 19125 22385 19159
rect 22385 19125 22419 19159
rect 22419 19125 22428 19159
rect 22376 19116 22428 19125
rect 23480 19159 23532 19168
rect 23480 19125 23489 19159
rect 23489 19125 23523 19159
rect 23523 19125 23532 19159
rect 23480 19116 23532 19125
rect 25044 19159 25096 19168
rect 25044 19125 25053 19159
rect 25053 19125 25087 19159
rect 25087 19125 25096 19159
rect 25044 19116 25096 19125
rect 25228 19116 25280 19168
rect 25688 19159 25740 19168
rect 25688 19125 25697 19159
rect 25697 19125 25731 19159
rect 25731 19125 25740 19159
rect 25688 19116 25740 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1400 18912 1452 18964
rect 3516 18912 3568 18964
rect 3792 18912 3844 18964
rect 6828 18912 6880 18964
rect 7472 18955 7524 18964
rect 7472 18921 7481 18955
rect 7481 18921 7515 18955
rect 7515 18921 7524 18955
rect 7472 18912 7524 18921
rect 7840 18955 7892 18964
rect 7840 18921 7849 18955
rect 7849 18921 7883 18955
rect 7883 18921 7892 18955
rect 7840 18912 7892 18921
rect 9680 18912 9732 18964
rect 11980 18955 12032 18964
rect 11980 18921 11989 18955
rect 11989 18921 12023 18955
rect 12023 18921 12032 18955
rect 11980 18912 12032 18921
rect 12532 18912 12584 18964
rect 13820 18955 13872 18964
rect 13820 18921 13829 18955
rect 13829 18921 13863 18955
rect 13863 18921 13872 18955
rect 13820 18912 13872 18921
rect 14648 18912 14700 18964
rect 16856 18912 16908 18964
rect 19064 18912 19116 18964
rect 19524 18912 19576 18964
rect 20076 18912 20128 18964
rect 20904 18912 20956 18964
rect 21088 18912 21140 18964
rect 21732 18912 21784 18964
rect 23296 18912 23348 18964
rect 4804 18844 4856 18896
rect 6276 18887 6328 18896
rect 5264 18819 5316 18828
rect 5264 18785 5273 18819
rect 5273 18785 5307 18819
rect 5307 18785 5316 18819
rect 5264 18776 5316 18785
rect 6276 18853 6285 18887
rect 6285 18853 6319 18887
rect 6319 18853 6328 18887
rect 6276 18844 6328 18853
rect 9404 18844 9456 18896
rect 10692 18844 10744 18896
rect 2044 18708 2096 18760
rect 2412 18751 2464 18760
rect 2412 18717 2421 18751
rect 2421 18717 2455 18751
rect 2455 18717 2464 18751
rect 2412 18708 2464 18717
rect 5172 18708 5224 18760
rect 6368 18776 6420 18828
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 12808 18844 12860 18896
rect 12992 18844 13044 18896
rect 16028 18844 16080 18896
rect 18236 18844 18288 18896
rect 18696 18887 18748 18896
rect 18696 18853 18705 18887
rect 18705 18853 18739 18887
rect 18739 18853 18748 18887
rect 18696 18844 18748 18853
rect 19340 18887 19392 18896
rect 19340 18853 19349 18887
rect 19349 18853 19383 18887
rect 19383 18853 19392 18887
rect 19340 18844 19392 18853
rect 12532 18776 12584 18828
rect 13728 18776 13780 18828
rect 14464 18819 14516 18828
rect 14464 18785 14473 18819
rect 14473 18785 14507 18819
rect 14507 18785 14516 18819
rect 14464 18776 14516 18785
rect 15384 18819 15436 18828
rect 15384 18785 15393 18819
rect 15393 18785 15427 18819
rect 15427 18785 15436 18819
rect 15384 18776 15436 18785
rect 16948 18819 17000 18828
rect 16948 18785 16982 18819
rect 16982 18785 17000 18819
rect 16948 18776 17000 18785
rect 17960 18776 18012 18828
rect 19156 18776 19208 18828
rect 6092 18708 6144 18760
rect 8484 18751 8536 18760
rect 6552 18640 6604 18692
rect 8484 18717 8493 18751
rect 8493 18717 8527 18751
rect 8527 18717 8536 18751
rect 8484 18708 8536 18717
rect 7656 18640 7708 18692
rect 10692 18708 10744 18760
rect 15660 18708 15712 18760
rect 16396 18708 16448 18760
rect 19984 18776 20036 18828
rect 21364 18751 21416 18760
rect 21364 18717 21373 18751
rect 21373 18717 21407 18751
rect 21407 18717 21416 18751
rect 21364 18708 21416 18717
rect 21548 18844 21600 18896
rect 22284 18844 22336 18896
rect 24952 18887 25004 18896
rect 24952 18853 24961 18887
rect 24961 18853 24995 18887
rect 24995 18853 25004 18887
rect 24952 18844 25004 18853
rect 25596 18887 25648 18896
rect 25596 18853 25605 18887
rect 25605 18853 25639 18887
rect 25639 18853 25648 18887
rect 25596 18844 25648 18853
rect 23020 18776 23072 18828
rect 21732 18708 21784 18760
rect 24768 18776 24820 18828
rect 23480 18751 23532 18760
rect 23480 18717 23489 18751
rect 23489 18717 23523 18751
rect 23523 18717 23532 18751
rect 23480 18708 23532 18717
rect 25044 18751 25096 18760
rect 25044 18717 25053 18751
rect 25053 18717 25087 18751
rect 25087 18717 25096 18751
rect 25044 18708 25096 18717
rect 9128 18640 9180 18692
rect 9588 18640 9640 18692
rect 22192 18640 22244 18692
rect 23572 18640 23624 18692
rect 25872 18640 25924 18692
rect 1860 18615 1912 18624
rect 1860 18581 1869 18615
rect 1869 18581 1903 18615
rect 1903 18581 1912 18615
rect 1860 18572 1912 18581
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 2228 18572 2280 18624
rect 3424 18615 3476 18624
rect 3424 18581 3433 18615
rect 3433 18581 3467 18615
rect 3467 18581 3476 18615
rect 3424 18572 3476 18581
rect 6460 18615 6512 18624
rect 6460 18581 6469 18615
rect 6469 18581 6503 18615
rect 6503 18581 6512 18615
rect 6460 18572 6512 18581
rect 8024 18615 8076 18624
rect 8024 18581 8033 18615
rect 8033 18581 8067 18615
rect 8067 18581 8076 18615
rect 8024 18572 8076 18581
rect 11060 18615 11112 18624
rect 11060 18581 11069 18615
rect 11069 18581 11103 18615
rect 11103 18581 11112 18615
rect 11060 18572 11112 18581
rect 11428 18615 11480 18624
rect 11428 18581 11437 18615
rect 11437 18581 11471 18615
rect 11471 18581 11480 18615
rect 11428 18572 11480 18581
rect 12348 18572 12400 18624
rect 14004 18572 14056 18624
rect 18144 18572 18196 18624
rect 20352 18615 20404 18624
rect 20352 18581 20361 18615
rect 20361 18581 20395 18615
rect 20395 18581 20404 18615
rect 20352 18572 20404 18581
rect 22928 18615 22980 18624
rect 22928 18581 22937 18615
rect 22937 18581 22971 18615
rect 22971 18581 22980 18615
rect 22928 18572 22980 18581
rect 23848 18572 23900 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1400 18368 1452 18420
rect 6552 18411 6604 18420
rect 6552 18377 6561 18411
rect 6561 18377 6595 18411
rect 6595 18377 6604 18411
rect 6552 18368 6604 18377
rect 8484 18368 8536 18420
rect 12072 18368 12124 18420
rect 12532 18368 12584 18420
rect 13268 18368 13320 18420
rect 13820 18411 13872 18420
rect 13820 18377 13829 18411
rect 13829 18377 13863 18411
rect 13863 18377 13872 18411
rect 13820 18368 13872 18377
rect 14372 18411 14424 18420
rect 14372 18377 14381 18411
rect 14381 18377 14415 18411
rect 14415 18377 14424 18411
rect 14372 18368 14424 18377
rect 15568 18368 15620 18420
rect 16948 18368 17000 18420
rect 19524 18411 19576 18420
rect 19524 18377 19533 18411
rect 19533 18377 19567 18411
rect 19567 18377 19576 18411
rect 19524 18368 19576 18377
rect 20352 18368 20404 18420
rect 21364 18368 21416 18420
rect 23296 18411 23348 18420
rect 23296 18377 23305 18411
rect 23305 18377 23339 18411
rect 23339 18377 23348 18411
rect 23296 18368 23348 18377
rect 23480 18368 23532 18420
rect 25872 18368 25924 18420
rect 5908 18300 5960 18352
rect 6736 18300 6788 18352
rect 9588 18300 9640 18352
rect 9956 18343 10008 18352
rect 9956 18309 9965 18343
rect 9965 18309 9999 18343
rect 9999 18309 10008 18343
rect 9956 18300 10008 18309
rect 1768 18164 1820 18216
rect 4160 18232 4212 18284
rect 11060 18275 11112 18284
rect 3516 18164 3568 18216
rect 3700 18164 3752 18216
rect 6092 18207 6144 18216
rect 6092 18173 6101 18207
rect 6101 18173 6135 18207
rect 6135 18173 6144 18207
rect 6092 18164 6144 18173
rect 6828 18207 6880 18216
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 8116 18164 8168 18216
rect 8944 18164 8996 18216
rect 11060 18241 11069 18275
rect 11069 18241 11103 18275
rect 11103 18241 11112 18275
rect 11060 18232 11112 18241
rect 12256 18275 12308 18284
rect 12256 18241 12265 18275
rect 12265 18241 12299 18275
rect 12299 18241 12308 18275
rect 12256 18232 12308 18241
rect 14004 18232 14056 18284
rect 14188 18232 14240 18284
rect 14464 18164 14516 18216
rect 21088 18300 21140 18352
rect 21548 18300 21600 18352
rect 16948 18232 17000 18284
rect 17500 18232 17552 18284
rect 18144 18232 18196 18284
rect 18972 18232 19024 18284
rect 19524 18232 19576 18284
rect 21916 18232 21968 18284
rect 25044 18232 25096 18284
rect 17776 18164 17828 18216
rect 18696 18164 18748 18216
rect 19248 18164 19300 18216
rect 22284 18207 22336 18216
rect 22284 18173 22293 18207
rect 22293 18173 22327 18207
rect 22327 18173 22336 18207
rect 22284 18164 22336 18173
rect 24860 18164 24912 18216
rect 2412 18139 2464 18148
rect 2412 18105 2446 18139
rect 2446 18105 2464 18139
rect 2412 18096 2464 18105
rect 3148 18096 3200 18148
rect 2044 18071 2096 18080
rect 2044 18037 2053 18071
rect 2053 18037 2087 18071
rect 2087 18037 2096 18071
rect 2044 18028 2096 18037
rect 2780 18028 2832 18080
rect 7104 18139 7156 18148
rect 7104 18105 7113 18139
rect 7113 18105 7147 18139
rect 7147 18105 7156 18139
rect 7104 18096 7156 18105
rect 10048 18096 10100 18148
rect 10876 18139 10928 18148
rect 3792 18071 3844 18080
rect 3792 18037 3801 18071
rect 3801 18037 3835 18071
rect 3835 18037 3844 18071
rect 3792 18028 3844 18037
rect 7656 18028 7708 18080
rect 9956 18028 10008 18080
rect 10876 18105 10885 18139
rect 10885 18105 10919 18139
rect 10919 18105 10928 18139
rect 10876 18096 10928 18105
rect 13452 18096 13504 18148
rect 12624 18071 12676 18080
rect 12624 18037 12633 18071
rect 12633 18037 12667 18071
rect 12667 18037 12676 18071
rect 12624 18028 12676 18037
rect 12808 18028 12860 18080
rect 14188 18071 14240 18080
rect 14188 18037 14197 18071
rect 14197 18037 14231 18071
rect 14231 18037 14240 18071
rect 14188 18028 14240 18037
rect 14372 18028 14424 18080
rect 17868 18096 17920 18148
rect 19984 18096 20036 18148
rect 22192 18139 22244 18148
rect 22192 18105 22201 18139
rect 22201 18105 22235 18139
rect 22235 18105 22244 18139
rect 22192 18096 22244 18105
rect 23848 18096 23900 18148
rect 25596 18096 25648 18148
rect 16856 18071 16908 18080
rect 16856 18037 16865 18071
rect 16865 18037 16899 18071
rect 16899 18037 16908 18071
rect 16856 18028 16908 18037
rect 17500 18071 17552 18080
rect 17500 18037 17509 18071
rect 17509 18037 17543 18071
rect 17543 18037 17552 18071
rect 17500 18028 17552 18037
rect 18236 18028 18288 18080
rect 20720 18028 20772 18080
rect 23020 18071 23072 18080
rect 23020 18037 23029 18071
rect 23029 18037 23063 18071
rect 23063 18037 23072 18071
rect 23020 18028 23072 18037
rect 23296 18028 23348 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 3148 17867 3200 17876
rect 3148 17833 3157 17867
rect 3157 17833 3191 17867
rect 3191 17833 3200 17867
rect 3148 17824 3200 17833
rect 3792 17824 3844 17876
rect 4252 17867 4304 17876
rect 4252 17833 4261 17867
rect 4261 17833 4295 17867
rect 4295 17833 4304 17867
rect 4252 17824 4304 17833
rect 4804 17824 4856 17876
rect 5264 17867 5316 17876
rect 5264 17833 5273 17867
rect 5273 17833 5307 17867
rect 5307 17833 5316 17867
rect 5264 17824 5316 17833
rect 8484 17824 8536 17876
rect 9404 17867 9456 17876
rect 9404 17833 9413 17867
rect 9413 17833 9447 17867
rect 9447 17833 9456 17867
rect 9404 17824 9456 17833
rect 10048 17824 10100 17876
rect 10876 17824 10928 17876
rect 12348 17824 12400 17876
rect 14372 17867 14424 17876
rect 14372 17833 14381 17867
rect 14381 17833 14415 17867
rect 14415 17833 14424 17867
rect 14372 17824 14424 17833
rect 15752 17824 15804 17876
rect 17500 17824 17552 17876
rect 17960 17824 18012 17876
rect 19984 17824 20036 17876
rect 20904 17867 20956 17876
rect 20904 17833 20913 17867
rect 20913 17833 20947 17867
rect 20947 17833 20956 17867
rect 20904 17824 20956 17833
rect 21364 17867 21416 17876
rect 21364 17833 21373 17867
rect 21373 17833 21407 17867
rect 21407 17833 21416 17867
rect 21364 17824 21416 17833
rect 22284 17867 22336 17876
rect 22284 17833 22293 17867
rect 22293 17833 22327 17867
rect 22327 17833 22336 17867
rect 22284 17824 22336 17833
rect 24952 17824 25004 17876
rect 25596 17824 25648 17876
rect 1768 17731 1820 17740
rect 1768 17697 1777 17731
rect 1777 17697 1811 17731
rect 1811 17697 1820 17731
rect 1768 17688 1820 17697
rect 1860 17688 1912 17740
rect 2596 17688 2648 17740
rect 4068 17731 4120 17740
rect 4068 17697 4077 17731
rect 4077 17697 4111 17731
rect 4111 17697 4120 17731
rect 4068 17688 4120 17697
rect 6276 17688 6328 17740
rect 6920 17688 6972 17740
rect 8116 17756 8168 17808
rect 10784 17756 10836 17808
rect 13820 17799 13872 17808
rect 13820 17765 13829 17799
rect 13829 17765 13863 17799
rect 13863 17765 13872 17799
rect 13820 17756 13872 17765
rect 14740 17756 14792 17808
rect 18052 17756 18104 17808
rect 19156 17756 19208 17808
rect 20720 17756 20772 17808
rect 21916 17799 21968 17808
rect 21916 17765 21925 17799
rect 21925 17765 21959 17799
rect 21959 17765 21968 17799
rect 21916 17756 21968 17765
rect 23756 17756 23808 17808
rect 7656 17731 7708 17740
rect 7656 17697 7690 17731
rect 7690 17697 7708 17731
rect 7656 17688 7708 17697
rect 9864 17731 9916 17740
rect 9864 17697 9873 17731
rect 9873 17697 9907 17731
rect 9907 17697 9916 17731
rect 9864 17688 9916 17697
rect 11428 17731 11480 17740
rect 11428 17697 11462 17731
rect 11462 17697 11480 17731
rect 11428 17688 11480 17697
rect 12256 17688 12308 17740
rect 13452 17688 13504 17740
rect 15568 17688 15620 17740
rect 16304 17731 16356 17740
rect 16304 17697 16313 17731
rect 16313 17697 16347 17731
rect 16347 17697 16356 17731
rect 16304 17688 16356 17697
rect 17684 17688 17736 17740
rect 4436 17620 4488 17672
rect 5908 17663 5960 17672
rect 5908 17629 5917 17663
rect 5917 17629 5951 17663
rect 5951 17629 5960 17663
rect 5908 17620 5960 17629
rect 10692 17620 10744 17672
rect 11060 17620 11112 17672
rect 13268 17620 13320 17672
rect 16396 17620 16448 17672
rect 18788 17620 18840 17672
rect 21548 17688 21600 17740
rect 24400 17731 24452 17740
rect 24400 17697 24409 17731
rect 24409 17697 24443 17731
rect 24443 17697 24452 17731
rect 24400 17688 24452 17697
rect 24768 17688 24820 17740
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 22192 17620 22244 17672
rect 22928 17663 22980 17672
rect 22928 17629 22937 17663
rect 22937 17629 22971 17663
rect 22971 17629 22980 17663
rect 22928 17620 22980 17629
rect 23020 17663 23072 17672
rect 23020 17629 23029 17663
rect 23029 17629 23063 17663
rect 23063 17629 23072 17663
rect 23020 17620 23072 17629
rect 23848 17620 23900 17672
rect 24676 17663 24728 17672
rect 24676 17629 24685 17663
rect 24685 17629 24719 17663
rect 24719 17629 24728 17663
rect 24676 17620 24728 17629
rect 8760 17595 8812 17604
rect 8760 17561 8769 17595
rect 8769 17561 8803 17595
rect 8803 17561 8812 17595
rect 8760 17552 8812 17561
rect 12808 17595 12860 17604
rect 12808 17561 12817 17595
rect 12817 17561 12851 17595
rect 12851 17561 12860 17595
rect 12808 17552 12860 17561
rect 13360 17595 13412 17604
rect 13360 17561 13369 17595
rect 13369 17561 13403 17595
rect 13403 17561 13412 17595
rect 13360 17552 13412 17561
rect 22008 17552 22060 17604
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 3240 17484 3292 17536
rect 6368 17484 6420 17536
rect 7196 17484 7248 17536
rect 9128 17484 9180 17536
rect 11152 17484 11204 17536
rect 12072 17484 12124 17536
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 14832 17527 14884 17536
rect 14832 17493 14841 17527
rect 14841 17493 14875 17527
rect 14875 17493 14884 17527
rect 14832 17484 14884 17493
rect 19064 17484 19116 17536
rect 23848 17484 23900 17536
rect 24032 17527 24084 17536
rect 24032 17493 24041 17527
rect 24041 17493 24075 17527
rect 24075 17493 24084 17527
rect 24032 17484 24084 17493
rect 25872 17484 25924 17536
rect 26148 17484 26200 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 3608 17323 3660 17332
rect 3608 17289 3617 17323
rect 3617 17289 3651 17323
rect 3651 17289 3660 17323
rect 3608 17280 3660 17289
rect 2596 17212 2648 17264
rect 6552 17280 6604 17332
rect 6736 17280 6788 17332
rect 7656 17280 7708 17332
rect 9864 17280 9916 17332
rect 11612 17323 11664 17332
rect 11612 17289 11621 17323
rect 11621 17289 11655 17323
rect 11655 17289 11664 17323
rect 11612 17280 11664 17289
rect 13452 17280 13504 17332
rect 14096 17323 14148 17332
rect 14096 17289 14105 17323
rect 14105 17289 14139 17323
rect 14139 17289 14148 17323
rect 14096 17280 14148 17289
rect 14740 17280 14792 17332
rect 17776 17323 17828 17332
rect 17776 17289 17785 17323
rect 17785 17289 17819 17323
rect 17819 17289 17828 17323
rect 17776 17280 17828 17289
rect 18052 17280 18104 17332
rect 18788 17323 18840 17332
rect 18788 17289 18797 17323
rect 18797 17289 18831 17323
rect 18831 17289 18840 17323
rect 18788 17280 18840 17289
rect 18880 17280 18932 17332
rect 23664 17323 23716 17332
rect 4436 17255 4488 17264
rect 4436 17221 4445 17255
rect 4445 17221 4479 17255
rect 4479 17221 4488 17255
rect 4436 17212 4488 17221
rect 11428 17212 11480 17264
rect 2688 17144 2740 17196
rect 4160 17144 4212 17196
rect 4344 17144 4396 17196
rect 6092 17144 6144 17196
rect 6552 17144 6604 17196
rect 7748 17144 7800 17196
rect 3240 17076 3292 17128
rect 8024 17119 8076 17128
rect 2964 17008 3016 17060
rect 8024 17085 8033 17119
rect 8033 17085 8067 17119
rect 8067 17085 8076 17119
rect 8024 17076 8076 17085
rect 10692 17187 10744 17196
rect 10692 17153 10701 17187
rect 10701 17153 10735 17187
rect 10735 17153 10744 17187
rect 10692 17144 10744 17153
rect 10876 17187 10928 17196
rect 10876 17153 10885 17187
rect 10885 17153 10919 17187
rect 10919 17153 10928 17187
rect 10876 17144 10928 17153
rect 14832 17144 14884 17196
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 8760 17076 8812 17128
rect 11060 17076 11112 17128
rect 12992 17076 13044 17128
rect 14648 17076 14700 17128
rect 17684 17212 17736 17264
rect 22928 17212 22980 17264
rect 15844 17144 15896 17196
rect 18972 17119 19024 17128
rect 18972 17085 18981 17119
rect 18981 17085 19015 17119
rect 19015 17085 19024 17119
rect 18972 17076 19024 17085
rect 19064 17076 19116 17128
rect 19248 17119 19300 17128
rect 19248 17085 19271 17119
rect 19271 17085 19300 17119
rect 19248 17076 19300 17085
rect 4988 17008 5040 17060
rect 10784 17008 10836 17060
rect 15016 17051 15068 17060
rect 1952 16940 2004 16992
rect 2228 16983 2280 16992
rect 2228 16949 2237 16983
rect 2237 16949 2271 16983
rect 2271 16949 2280 16983
rect 2228 16940 2280 16949
rect 4068 16983 4120 16992
rect 4068 16949 4077 16983
rect 4077 16949 4111 16983
rect 4111 16949 4120 16983
rect 4068 16940 4120 16949
rect 6276 16983 6328 16992
rect 6276 16949 6285 16983
rect 6285 16949 6319 16983
rect 6319 16949 6328 16983
rect 6276 16940 6328 16949
rect 9404 16983 9456 16992
rect 9404 16949 9413 16983
rect 9413 16949 9447 16983
rect 9447 16949 9456 16983
rect 9404 16940 9456 16949
rect 10140 16940 10192 16992
rect 12164 16983 12216 16992
rect 12164 16949 12173 16983
rect 12173 16949 12207 16983
rect 12207 16949 12216 16983
rect 12164 16940 12216 16949
rect 12532 16940 12584 16992
rect 15016 17017 15025 17051
rect 15025 17017 15059 17051
rect 15059 17017 15068 17051
rect 15016 17008 15068 17017
rect 16304 17008 16356 17060
rect 21732 17076 21784 17128
rect 22652 17076 22704 17128
rect 22928 17076 22980 17128
rect 23664 17289 23673 17323
rect 23673 17289 23707 17323
rect 23707 17289 23716 17323
rect 23664 17280 23716 17289
rect 25412 17212 25464 17264
rect 26148 17212 26200 17264
rect 24676 17144 24728 17196
rect 25228 17119 25280 17128
rect 25228 17085 25237 17119
rect 25237 17085 25271 17119
rect 25271 17085 25280 17119
rect 25228 17076 25280 17085
rect 19524 17008 19576 17060
rect 21456 17051 21508 17060
rect 21456 17017 21490 17051
rect 21490 17017 21508 17051
rect 14004 16940 14056 16992
rect 16212 16983 16264 16992
rect 16212 16949 16221 16983
rect 16221 16949 16255 16983
rect 16255 16949 16264 16983
rect 16212 16940 16264 16949
rect 21456 17008 21508 17017
rect 21916 17008 21968 17060
rect 25412 17008 25464 17060
rect 22652 16940 22704 16992
rect 23848 16940 23900 16992
rect 24032 16983 24084 16992
rect 24032 16949 24041 16983
rect 24041 16949 24075 16983
rect 24075 16949 24084 16983
rect 24032 16940 24084 16949
rect 24676 16983 24728 16992
rect 24676 16949 24685 16983
rect 24685 16949 24719 16983
rect 24719 16949 24728 16983
rect 24676 16940 24728 16949
rect 25596 16940 25648 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2228 16736 2280 16788
rect 3700 16736 3752 16788
rect 5172 16779 5224 16788
rect 5172 16745 5181 16779
rect 5181 16745 5215 16779
rect 5215 16745 5224 16779
rect 5172 16736 5224 16745
rect 5356 16736 5408 16788
rect 6184 16736 6236 16788
rect 6920 16779 6972 16788
rect 6920 16745 6929 16779
rect 6929 16745 6963 16779
rect 6963 16745 6972 16779
rect 6920 16736 6972 16745
rect 8392 16736 8444 16788
rect 10140 16736 10192 16788
rect 10876 16736 10928 16788
rect 13728 16736 13780 16788
rect 14648 16779 14700 16788
rect 14648 16745 14657 16779
rect 14657 16745 14691 16779
rect 14691 16745 14700 16779
rect 14648 16736 14700 16745
rect 15016 16779 15068 16788
rect 15016 16745 15025 16779
rect 15025 16745 15059 16779
rect 15059 16745 15068 16779
rect 15016 16736 15068 16745
rect 16856 16736 16908 16788
rect 19064 16736 19116 16788
rect 19248 16736 19300 16788
rect 19984 16736 20036 16788
rect 2872 16711 2924 16720
rect 2872 16677 2881 16711
rect 2881 16677 2915 16711
rect 2915 16677 2924 16711
rect 2872 16668 2924 16677
rect 3332 16711 3384 16720
rect 3332 16677 3341 16711
rect 3341 16677 3375 16711
rect 3375 16677 3384 16711
rect 3332 16668 3384 16677
rect 6460 16668 6512 16720
rect 7656 16711 7708 16720
rect 7656 16677 7665 16711
rect 7665 16677 7699 16711
rect 7699 16677 7708 16711
rect 7656 16668 7708 16677
rect 8760 16668 8812 16720
rect 1768 16600 1820 16652
rect 3056 16600 3108 16652
rect 3608 16600 3660 16652
rect 2228 16575 2280 16584
rect 2228 16541 2237 16575
rect 2237 16541 2271 16575
rect 2271 16541 2280 16575
rect 2228 16532 2280 16541
rect 2412 16575 2464 16584
rect 2412 16541 2421 16575
rect 2421 16541 2455 16575
rect 2455 16541 2464 16575
rect 2412 16532 2464 16541
rect 6184 16600 6236 16652
rect 6552 16643 6604 16652
rect 4160 16532 4212 16584
rect 6000 16532 6052 16584
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 6736 16643 6788 16652
rect 6736 16609 6745 16643
rect 6745 16609 6779 16643
rect 6779 16609 6788 16643
rect 6736 16600 6788 16609
rect 8208 16643 8260 16652
rect 8208 16609 8217 16643
rect 8217 16609 8251 16643
rect 8251 16609 8260 16643
rect 8208 16600 8260 16609
rect 9864 16643 9916 16652
rect 9864 16609 9873 16643
rect 9873 16609 9907 16643
rect 9907 16609 9916 16643
rect 9864 16600 9916 16609
rect 10968 16600 11020 16652
rect 11060 16600 11112 16652
rect 11428 16643 11480 16652
rect 11428 16609 11462 16643
rect 11462 16609 11480 16643
rect 11428 16600 11480 16609
rect 11796 16600 11848 16652
rect 13268 16600 13320 16652
rect 13544 16600 13596 16652
rect 16304 16668 16356 16720
rect 16764 16668 16816 16720
rect 21272 16736 21324 16788
rect 21916 16779 21968 16788
rect 21916 16745 21925 16779
rect 21925 16745 21959 16779
rect 21959 16745 21968 16779
rect 21916 16736 21968 16745
rect 23020 16736 23072 16788
rect 24860 16779 24912 16788
rect 24860 16745 24869 16779
rect 24869 16745 24903 16779
rect 24903 16745 24912 16779
rect 24860 16736 24912 16745
rect 25136 16779 25188 16788
rect 25136 16745 25145 16779
rect 25145 16745 25179 16779
rect 25179 16745 25188 16779
rect 25136 16736 25188 16745
rect 15752 16643 15804 16652
rect 15752 16609 15786 16643
rect 15786 16609 15804 16643
rect 15752 16600 15804 16609
rect 4804 16464 4856 16516
rect 8944 16532 8996 16584
rect 12900 16532 12952 16584
rect 13912 16575 13964 16584
rect 13912 16541 13921 16575
rect 13921 16541 13955 16575
rect 13955 16541 13964 16575
rect 13912 16532 13964 16541
rect 17224 16532 17276 16584
rect 17776 16532 17828 16584
rect 20628 16600 20680 16652
rect 21732 16600 21784 16652
rect 22376 16600 22428 16652
rect 25596 16668 25648 16720
rect 23020 16643 23072 16652
rect 23020 16609 23054 16643
rect 23054 16609 23072 16643
rect 23020 16600 23072 16609
rect 24952 16643 25004 16652
rect 24952 16609 24961 16643
rect 24961 16609 24995 16643
rect 24995 16609 25004 16643
rect 24952 16600 25004 16609
rect 8208 16464 8260 16516
rect 17040 16464 17092 16516
rect 18512 16532 18564 16584
rect 19708 16575 19760 16584
rect 19708 16541 19717 16575
rect 19717 16541 19751 16575
rect 19751 16541 19760 16575
rect 19708 16532 19760 16541
rect 19156 16464 19208 16516
rect 19340 16464 19392 16516
rect 21088 16532 21140 16584
rect 22008 16532 22060 16584
rect 22468 16532 22520 16584
rect 23848 16464 23900 16516
rect 24124 16464 24176 16516
rect 1768 16396 1820 16448
rect 4988 16396 5040 16448
rect 5172 16396 5224 16448
rect 6276 16439 6328 16448
rect 6276 16405 6285 16439
rect 6285 16405 6319 16439
rect 6319 16405 6328 16439
rect 6276 16396 6328 16405
rect 7012 16396 7064 16448
rect 7104 16396 7156 16448
rect 11060 16439 11112 16448
rect 11060 16405 11069 16439
rect 11069 16405 11103 16439
rect 11103 16405 11112 16439
rect 11060 16396 11112 16405
rect 12532 16439 12584 16448
rect 12532 16405 12541 16439
rect 12541 16405 12575 16439
rect 12575 16405 12584 16439
rect 12532 16396 12584 16405
rect 13452 16396 13504 16448
rect 17408 16396 17460 16448
rect 20628 16439 20680 16448
rect 20628 16405 20637 16439
rect 20637 16405 20671 16439
rect 20671 16405 20680 16439
rect 20628 16396 20680 16405
rect 22468 16396 22520 16448
rect 24860 16396 24912 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2412 16192 2464 16244
rect 2688 16235 2740 16244
rect 2688 16201 2697 16235
rect 2697 16201 2731 16235
rect 2731 16201 2740 16235
rect 2688 16192 2740 16201
rect 4344 16192 4396 16244
rect 5356 16192 5408 16244
rect 6000 16192 6052 16244
rect 8116 16192 8168 16244
rect 8944 16192 8996 16244
rect 9680 16235 9732 16244
rect 9680 16201 9689 16235
rect 9689 16201 9723 16235
rect 9723 16201 9732 16235
rect 9680 16192 9732 16201
rect 11428 16192 11480 16244
rect 13544 16235 13596 16244
rect 13544 16201 13553 16235
rect 13553 16201 13587 16235
rect 13587 16201 13596 16235
rect 13544 16192 13596 16201
rect 13820 16192 13872 16244
rect 17040 16235 17092 16244
rect 17040 16201 17049 16235
rect 17049 16201 17083 16235
rect 17083 16201 17092 16235
rect 17040 16192 17092 16201
rect 19708 16192 19760 16244
rect 21272 16192 21324 16244
rect 22192 16192 22244 16244
rect 2964 16124 3016 16176
rect 5448 16124 5500 16176
rect 6184 16167 6236 16176
rect 6184 16133 6193 16167
rect 6193 16133 6227 16167
rect 6227 16133 6236 16167
rect 6184 16124 6236 16133
rect 2780 16056 2832 16108
rect 6000 16056 6052 16108
rect 11060 16056 11112 16108
rect 12164 16124 12216 16176
rect 12532 16124 12584 16176
rect 19984 16167 20036 16176
rect 19984 16133 19993 16167
rect 19993 16133 20027 16167
rect 20027 16133 20036 16167
rect 19984 16124 20036 16133
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 13544 16056 13596 16108
rect 13912 16056 13964 16108
rect 14372 16056 14424 16108
rect 15752 16056 15804 16108
rect 16672 16056 16724 16108
rect 21088 16099 21140 16108
rect 21088 16065 21097 16099
rect 21097 16065 21131 16099
rect 21131 16065 21140 16099
rect 21088 16056 21140 16065
rect 1768 15988 1820 16040
rect 2872 15988 2924 16040
rect 4804 15988 4856 16040
rect 5172 15988 5224 16040
rect 7104 15988 7156 16040
rect 7932 16031 7984 16040
rect 7932 15997 7941 16031
rect 7941 15997 7975 16031
rect 7975 15997 7984 16031
rect 7932 15988 7984 15997
rect 14464 16031 14516 16040
rect 14464 15997 14473 16031
rect 14473 15997 14507 16031
rect 14507 15997 14516 16031
rect 14464 15988 14516 15997
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 1492 15920 1544 15972
rect 2412 15920 2464 15972
rect 3332 15852 3384 15904
rect 4160 15895 4212 15904
rect 4160 15861 4169 15895
rect 4169 15861 4203 15895
rect 4203 15861 4212 15895
rect 4160 15852 4212 15861
rect 5264 15852 5316 15904
rect 6276 15852 6328 15904
rect 6644 15852 6696 15904
rect 9404 15920 9456 15972
rect 10140 15920 10192 15972
rect 11336 15920 11388 15972
rect 12624 15920 12676 15972
rect 9036 15852 9088 15904
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 12440 15895 12492 15904
rect 12440 15861 12449 15895
rect 12449 15861 12483 15895
rect 12483 15861 12492 15895
rect 13084 15920 13136 15972
rect 14556 15920 14608 15972
rect 17224 15920 17276 15972
rect 18144 15920 18196 15972
rect 21088 15920 21140 15972
rect 12440 15852 12492 15861
rect 12992 15852 13044 15904
rect 13360 15852 13412 15904
rect 13636 15852 13688 15904
rect 15568 15895 15620 15904
rect 15568 15861 15577 15895
rect 15577 15861 15611 15895
rect 15611 15861 15620 15895
rect 15568 15852 15620 15861
rect 15936 15895 15988 15904
rect 15936 15861 15945 15895
rect 15945 15861 15979 15895
rect 15979 15861 15988 15895
rect 15936 15852 15988 15861
rect 16120 15852 16172 15904
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 17776 15895 17828 15904
rect 17776 15861 17785 15895
rect 17785 15861 17819 15895
rect 17819 15861 17828 15895
rect 17776 15852 17828 15861
rect 20260 15852 20312 15904
rect 20904 15895 20956 15904
rect 20904 15861 20913 15895
rect 20913 15861 20947 15895
rect 20947 15861 20956 15895
rect 20904 15852 20956 15861
rect 23020 16124 23072 16176
rect 23756 16192 23808 16244
rect 24952 16235 25004 16244
rect 24952 16201 24961 16235
rect 24961 16201 24995 16235
rect 24995 16201 25004 16235
rect 24952 16192 25004 16201
rect 25504 16192 25556 16244
rect 25596 16192 25648 16244
rect 26240 16124 26292 16176
rect 22560 16099 22612 16108
rect 22560 16065 22569 16099
rect 22569 16065 22603 16099
rect 22603 16065 22612 16099
rect 22560 16056 22612 16065
rect 22744 16056 22796 16108
rect 24216 16099 24268 16108
rect 24216 16065 24225 16099
rect 24225 16065 24259 16099
rect 24259 16065 24268 16099
rect 24216 16056 24268 16065
rect 22192 15988 22244 16040
rect 25228 16031 25280 16040
rect 22468 15895 22520 15904
rect 22468 15861 22477 15895
rect 22477 15861 22511 15895
rect 22511 15861 22520 15895
rect 22468 15852 22520 15861
rect 23112 15852 23164 15904
rect 25228 15997 25237 16031
rect 25237 15997 25271 16031
rect 25271 15997 25280 16031
rect 25228 15988 25280 15997
rect 24768 15852 24820 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2228 15648 2280 15700
rect 4344 15648 4396 15700
rect 8208 15648 8260 15700
rect 8484 15648 8536 15700
rect 9312 15648 9364 15700
rect 11060 15648 11112 15700
rect 13452 15691 13504 15700
rect 13452 15657 13461 15691
rect 13461 15657 13495 15691
rect 13495 15657 13504 15691
rect 13452 15648 13504 15657
rect 14372 15691 14424 15700
rect 14372 15657 14381 15691
rect 14381 15657 14415 15691
rect 14415 15657 14424 15691
rect 14372 15648 14424 15657
rect 16672 15691 16724 15700
rect 16672 15657 16681 15691
rect 16681 15657 16715 15691
rect 16715 15657 16724 15691
rect 16672 15648 16724 15657
rect 17408 15691 17460 15700
rect 17408 15657 17417 15691
rect 17417 15657 17451 15691
rect 17451 15657 17460 15691
rect 17408 15648 17460 15657
rect 17684 15691 17736 15700
rect 17684 15657 17693 15691
rect 17693 15657 17727 15691
rect 17727 15657 17736 15691
rect 17684 15648 17736 15657
rect 18144 15691 18196 15700
rect 18144 15657 18153 15691
rect 18153 15657 18187 15691
rect 18187 15657 18196 15691
rect 18144 15648 18196 15657
rect 18512 15691 18564 15700
rect 18512 15657 18521 15691
rect 18521 15657 18555 15691
rect 18555 15657 18564 15691
rect 18512 15648 18564 15657
rect 19340 15648 19392 15700
rect 19984 15691 20036 15700
rect 19984 15657 19993 15691
rect 19993 15657 20027 15691
rect 20027 15657 20036 15691
rect 19984 15648 20036 15657
rect 20812 15648 20864 15700
rect 2412 15623 2464 15632
rect 2412 15589 2421 15623
rect 2421 15589 2455 15623
rect 2455 15589 2464 15623
rect 2412 15580 2464 15589
rect 2320 15555 2372 15564
rect 2320 15521 2329 15555
rect 2329 15521 2363 15555
rect 2363 15521 2372 15555
rect 2320 15512 2372 15521
rect 2780 15512 2832 15564
rect 7656 15580 7708 15632
rect 8944 15580 8996 15632
rect 11152 15580 11204 15632
rect 12348 15580 12400 15632
rect 12440 15580 12492 15632
rect 16396 15580 16448 15632
rect 20720 15580 20772 15632
rect 22560 15648 22612 15700
rect 24216 15648 24268 15700
rect 25044 15648 25096 15700
rect 21456 15580 21508 15632
rect 22652 15580 22704 15632
rect 4160 15512 4212 15564
rect 6460 15512 6512 15564
rect 8392 15512 8444 15564
rect 11060 15555 11112 15564
rect 11060 15521 11094 15555
rect 11094 15521 11112 15555
rect 11060 15512 11112 15521
rect 11888 15512 11940 15564
rect 12900 15555 12952 15564
rect 12900 15521 12909 15555
rect 12909 15521 12943 15555
rect 12943 15521 12952 15555
rect 12900 15512 12952 15521
rect 14464 15512 14516 15564
rect 15844 15512 15896 15564
rect 17316 15512 17368 15564
rect 18880 15555 18932 15564
rect 18880 15521 18914 15555
rect 18914 15521 18932 15555
rect 18880 15512 18932 15521
rect 20536 15512 20588 15564
rect 22376 15512 22428 15564
rect 23296 15512 23348 15564
rect 25044 15555 25096 15564
rect 25044 15521 25053 15555
rect 25053 15521 25087 15555
rect 25087 15521 25096 15555
rect 25044 15512 25096 15521
rect 2228 15376 2280 15428
rect 2596 15444 2648 15496
rect 3884 15487 3936 15496
rect 3884 15453 3893 15487
rect 3893 15453 3927 15487
rect 3927 15453 3936 15487
rect 3884 15444 3936 15453
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 5540 15376 5592 15428
rect 1676 15351 1728 15360
rect 1676 15317 1685 15351
rect 1685 15317 1719 15351
rect 1719 15317 1728 15351
rect 1676 15308 1728 15317
rect 3056 15351 3108 15360
rect 3056 15317 3065 15351
rect 3065 15317 3099 15351
rect 3099 15317 3108 15351
rect 3056 15308 3108 15317
rect 4804 15308 4856 15360
rect 4988 15308 5040 15360
rect 6000 15308 6052 15360
rect 9404 15444 9456 15496
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 9864 15444 9916 15496
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 10692 15444 10744 15496
rect 12440 15444 12492 15496
rect 13452 15444 13504 15496
rect 13636 15487 13688 15496
rect 13636 15453 13645 15487
rect 13645 15453 13679 15487
rect 13679 15453 13688 15487
rect 13636 15444 13688 15453
rect 15292 15487 15344 15496
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 7564 15308 7616 15360
rect 7932 15308 7984 15360
rect 9680 15308 9732 15360
rect 11428 15308 11480 15360
rect 12164 15351 12216 15360
rect 12164 15317 12173 15351
rect 12173 15317 12207 15351
rect 12207 15317 12216 15351
rect 12164 15308 12216 15317
rect 13084 15308 13136 15360
rect 15936 15308 15988 15360
rect 20260 15444 20312 15496
rect 23756 15444 23808 15496
rect 24860 15444 24912 15496
rect 25320 15487 25372 15496
rect 25320 15453 25329 15487
rect 25329 15453 25363 15487
rect 25363 15453 25372 15487
rect 25320 15444 25372 15453
rect 24124 15376 24176 15428
rect 18972 15308 19024 15360
rect 19248 15308 19300 15360
rect 20720 15308 20772 15360
rect 20812 15308 20864 15360
rect 22744 15308 22796 15360
rect 23664 15308 23716 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2320 15104 2372 15156
rect 5172 15147 5224 15156
rect 5172 15113 5181 15147
rect 5181 15113 5215 15147
rect 5215 15113 5224 15147
rect 5172 15104 5224 15113
rect 6276 15104 6328 15156
rect 7012 15147 7064 15156
rect 7012 15113 7021 15147
rect 7021 15113 7055 15147
rect 7055 15113 7064 15147
rect 7012 15104 7064 15113
rect 8484 15147 8536 15156
rect 8484 15113 8493 15147
rect 8493 15113 8527 15147
rect 8527 15113 8536 15147
rect 8484 15104 8536 15113
rect 9404 15104 9456 15156
rect 11060 15104 11112 15156
rect 12164 15147 12216 15156
rect 12164 15113 12173 15147
rect 12173 15113 12207 15147
rect 12207 15113 12216 15147
rect 12164 15104 12216 15113
rect 12348 15104 12400 15156
rect 13544 15147 13596 15156
rect 13544 15113 13553 15147
rect 13553 15113 13587 15147
rect 13587 15113 13596 15147
rect 13544 15104 13596 15113
rect 13636 15104 13688 15156
rect 17040 15147 17092 15156
rect 17040 15113 17049 15147
rect 17049 15113 17083 15147
rect 17083 15113 17092 15147
rect 17040 15104 17092 15113
rect 17868 15147 17920 15156
rect 17868 15113 17877 15147
rect 17877 15113 17911 15147
rect 17911 15113 17920 15147
rect 17868 15104 17920 15113
rect 18880 15104 18932 15156
rect 20260 15147 20312 15156
rect 20260 15113 20269 15147
rect 20269 15113 20303 15147
rect 20303 15113 20312 15147
rect 20260 15104 20312 15113
rect 22008 15104 22060 15156
rect 22376 15104 22428 15156
rect 22652 15147 22704 15156
rect 22652 15113 22661 15147
rect 22661 15113 22695 15147
rect 22695 15113 22704 15147
rect 22652 15104 22704 15113
rect 23940 15104 23992 15156
rect 24768 15147 24820 15156
rect 24768 15113 24777 15147
rect 24777 15113 24811 15147
rect 24811 15113 24820 15147
rect 24768 15104 24820 15113
rect 25320 15104 25372 15156
rect 2412 15036 2464 15088
rect 8392 15036 8444 15088
rect 1676 14968 1728 15020
rect 2780 15011 2832 15020
rect 2780 14977 2789 15011
rect 2789 14977 2823 15011
rect 2823 14977 2832 15011
rect 2780 14968 2832 14977
rect 6552 14968 6604 15020
rect 7656 15011 7708 15020
rect 7656 14977 7665 15011
rect 7665 14977 7699 15011
rect 7699 14977 7708 15011
rect 7656 14968 7708 14977
rect 8576 15011 8628 15020
rect 8576 14977 8585 15011
rect 8585 14977 8619 15011
rect 8619 14977 8628 15011
rect 8576 14968 8628 14977
rect 12440 14968 12492 15020
rect 22192 15036 22244 15088
rect 22560 15036 22612 15088
rect 24676 15036 24728 15088
rect 17224 14968 17276 15020
rect 1676 14875 1728 14884
rect 1676 14841 1685 14875
rect 1685 14841 1719 14875
rect 1719 14841 1728 14875
rect 1676 14832 1728 14841
rect 3056 14943 3108 14952
rect 3056 14909 3090 14943
rect 3090 14909 3108 14943
rect 3056 14900 3108 14909
rect 5540 14943 5592 14952
rect 5540 14909 5549 14943
rect 5549 14909 5583 14943
rect 5583 14909 5592 14943
rect 5540 14900 5592 14909
rect 6276 14943 6328 14952
rect 6276 14909 6285 14943
rect 6285 14909 6319 14943
rect 6319 14909 6328 14943
rect 9772 14943 9824 14952
rect 6276 14900 6328 14909
rect 9772 14909 9781 14943
rect 9781 14909 9815 14943
rect 9815 14909 9824 14943
rect 9772 14900 9824 14909
rect 13728 14900 13780 14952
rect 14372 14900 14424 14952
rect 15292 14900 15344 14952
rect 2964 14832 3016 14884
rect 7380 14875 7432 14884
rect 7380 14841 7389 14875
rect 7389 14841 7423 14875
rect 7423 14841 7432 14875
rect 7380 14832 7432 14841
rect 10140 14832 10192 14884
rect 10692 14832 10744 14884
rect 14740 14832 14792 14884
rect 17776 14900 17828 14952
rect 18052 14900 18104 14952
rect 20812 15011 20864 15020
rect 20812 14977 20821 15011
rect 20821 14977 20855 15011
rect 20855 14977 20864 15011
rect 20812 14968 20864 14977
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 20168 14900 20220 14952
rect 20536 14900 20588 14952
rect 21916 14943 21968 14952
rect 21916 14909 21925 14943
rect 21925 14909 21959 14943
rect 21959 14909 21968 14943
rect 21916 14900 21968 14909
rect 23664 14900 23716 14952
rect 19248 14832 19300 14884
rect 19984 14832 20036 14884
rect 20812 14832 20864 14884
rect 21456 14832 21508 14884
rect 22192 14875 22244 14884
rect 22192 14841 22201 14875
rect 22201 14841 22235 14875
rect 22235 14841 22244 14875
rect 22192 14832 22244 14841
rect 23480 14875 23532 14884
rect 23480 14841 23489 14875
rect 23489 14841 23523 14875
rect 23523 14841 23532 14875
rect 23480 14832 23532 14841
rect 2780 14764 2832 14816
rect 4160 14807 4212 14816
rect 4160 14773 4169 14807
rect 4169 14773 4203 14807
rect 4203 14773 4212 14807
rect 4160 14764 4212 14773
rect 5632 14807 5684 14816
rect 5632 14773 5641 14807
rect 5641 14773 5675 14807
rect 5675 14773 5684 14807
rect 5632 14764 5684 14773
rect 7564 14764 7616 14816
rect 12808 14807 12860 14816
rect 12808 14773 12817 14807
rect 12817 14773 12851 14807
rect 12851 14773 12860 14807
rect 12808 14764 12860 14773
rect 15844 14764 15896 14816
rect 16120 14764 16172 14816
rect 16672 14807 16724 14816
rect 16672 14773 16681 14807
rect 16681 14773 16715 14807
rect 16715 14773 16724 14807
rect 16672 14764 16724 14773
rect 20352 14807 20404 14816
rect 20352 14773 20361 14807
rect 20361 14773 20395 14807
rect 20395 14773 20404 14807
rect 20352 14764 20404 14773
rect 21824 14764 21876 14816
rect 22652 14764 22704 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2228 14560 2280 14612
rect 2504 14560 2556 14612
rect 3608 14560 3660 14612
rect 3884 14603 3936 14612
rect 3884 14569 3893 14603
rect 3893 14569 3927 14603
rect 3927 14569 3936 14603
rect 3884 14560 3936 14569
rect 6736 14560 6788 14612
rect 8024 14603 8076 14612
rect 8024 14569 8033 14603
rect 8033 14569 8067 14603
rect 8067 14569 8076 14603
rect 8024 14560 8076 14569
rect 8484 14560 8536 14612
rect 8760 14560 8812 14612
rect 9772 14560 9824 14612
rect 4896 14492 4948 14544
rect 5356 14535 5408 14544
rect 5356 14501 5365 14535
rect 5365 14501 5399 14535
rect 5399 14501 5408 14535
rect 5356 14492 5408 14501
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 4712 14467 4764 14476
rect 2780 14424 2832 14433
rect 4712 14433 4721 14467
rect 4721 14433 4755 14467
rect 4755 14433 4764 14467
rect 4712 14424 4764 14433
rect 5448 14424 5500 14476
rect 2044 14356 2096 14408
rect 4804 14356 4856 14408
rect 6276 14492 6328 14544
rect 10784 14560 10836 14612
rect 10968 14603 11020 14612
rect 10968 14569 10977 14603
rect 10977 14569 11011 14603
rect 11011 14569 11020 14603
rect 10968 14560 11020 14569
rect 12624 14560 12676 14612
rect 6828 14424 6880 14476
rect 8392 14424 8444 14476
rect 11980 14492 12032 14544
rect 12808 14560 12860 14612
rect 16396 14560 16448 14612
rect 16580 14560 16632 14612
rect 17316 14560 17368 14612
rect 19248 14603 19300 14612
rect 19248 14569 19257 14603
rect 19257 14569 19291 14603
rect 19291 14569 19300 14603
rect 19248 14560 19300 14569
rect 20904 14560 20956 14612
rect 20996 14560 21048 14612
rect 21548 14603 21600 14612
rect 21548 14569 21557 14603
rect 21557 14569 21591 14603
rect 21591 14569 21600 14603
rect 21548 14560 21600 14569
rect 22008 14603 22060 14612
rect 22008 14569 22017 14603
rect 22017 14569 22051 14603
rect 22051 14569 22060 14603
rect 22008 14560 22060 14569
rect 22468 14560 22520 14612
rect 22928 14560 22980 14612
rect 23112 14560 23164 14612
rect 23296 14560 23348 14612
rect 25136 14560 25188 14612
rect 13728 14535 13780 14544
rect 13728 14501 13737 14535
rect 13737 14501 13771 14535
rect 13771 14501 13780 14535
rect 13728 14492 13780 14501
rect 15384 14492 15436 14544
rect 16488 14492 16540 14544
rect 17592 14492 17644 14544
rect 19616 14492 19668 14544
rect 20260 14492 20312 14544
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 10692 14424 10744 14476
rect 13544 14424 13596 14476
rect 7472 14399 7524 14408
rect 1952 14288 2004 14340
rect 3884 14288 3936 14340
rect 7472 14365 7481 14399
rect 7481 14365 7515 14399
rect 7515 14365 7524 14399
rect 7472 14356 7524 14365
rect 10140 14356 10192 14408
rect 12808 14356 12860 14408
rect 13728 14356 13780 14408
rect 20536 14424 20588 14476
rect 20996 14424 21048 14476
rect 21364 14424 21416 14476
rect 22376 14424 22428 14476
rect 23388 14424 23440 14476
rect 24216 14467 24268 14476
rect 24216 14433 24225 14467
rect 24225 14433 24259 14467
rect 24259 14433 24268 14467
rect 24216 14424 24268 14433
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 16764 14356 16816 14408
rect 17592 14356 17644 14408
rect 17776 14356 17828 14408
rect 19984 14399 20036 14408
rect 19984 14365 19993 14399
rect 19993 14365 20027 14399
rect 20027 14365 20036 14399
rect 19984 14356 20036 14365
rect 20168 14356 20220 14408
rect 23112 14399 23164 14408
rect 23112 14365 23121 14399
rect 23121 14365 23155 14399
rect 23155 14365 23164 14399
rect 23112 14356 23164 14365
rect 16304 14331 16356 14340
rect 16304 14297 16313 14331
rect 16313 14297 16347 14331
rect 16347 14297 16356 14331
rect 16304 14288 16356 14297
rect 20904 14288 20956 14340
rect 21640 14288 21692 14340
rect 21824 14288 21876 14340
rect 24676 14356 24728 14408
rect 3240 14263 3292 14272
rect 3240 14229 3249 14263
rect 3249 14229 3283 14263
rect 3283 14229 3292 14263
rect 3240 14220 3292 14229
rect 6000 14220 6052 14272
rect 9680 14220 9732 14272
rect 11796 14220 11848 14272
rect 12164 14220 12216 14272
rect 14004 14220 14056 14272
rect 14648 14263 14700 14272
rect 14648 14229 14657 14263
rect 14657 14229 14691 14263
rect 14691 14229 14700 14263
rect 14648 14220 14700 14229
rect 15844 14263 15896 14272
rect 15844 14229 15853 14263
rect 15853 14229 15887 14263
rect 15887 14229 15896 14263
rect 15844 14220 15896 14229
rect 19340 14220 19392 14272
rect 19524 14220 19576 14272
rect 22284 14220 22336 14272
rect 22560 14220 22612 14272
rect 23664 14263 23716 14272
rect 23664 14229 23673 14263
rect 23673 14229 23707 14263
rect 23707 14229 23716 14263
rect 23664 14220 23716 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1860 13880 1912 13932
rect 1952 13812 2004 13864
rect 3056 14016 3108 14068
rect 4712 14016 4764 14068
rect 4896 14059 4948 14068
rect 4896 14025 4905 14059
rect 4905 14025 4939 14059
rect 4939 14025 4948 14059
rect 4896 14016 4948 14025
rect 5172 14059 5224 14068
rect 5172 14025 5181 14059
rect 5181 14025 5215 14059
rect 5215 14025 5224 14059
rect 5172 14016 5224 14025
rect 6276 14059 6328 14068
rect 6276 14025 6285 14059
rect 6285 14025 6319 14059
rect 6319 14025 6328 14059
rect 6276 14016 6328 14025
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 8484 14016 8536 14068
rect 10140 14016 10192 14068
rect 14740 14016 14792 14068
rect 16028 14016 16080 14068
rect 16488 14016 16540 14068
rect 17592 14016 17644 14068
rect 17868 14059 17920 14068
rect 17868 14025 17877 14059
rect 17877 14025 17911 14059
rect 17911 14025 17920 14059
rect 17868 14016 17920 14025
rect 2964 13812 3016 13864
rect 5540 13880 5592 13932
rect 5632 13880 5684 13932
rect 12440 13991 12492 14000
rect 12440 13957 12449 13991
rect 12449 13957 12483 13991
rect 12483 13957 12492 13991
rect 12440 13948 12492 13957
rect 17408 13948 17460 14000
rect 5356 13812 5408 13864
rect 6828 13855 6880 13864
rect 3608 13744 3660 13796
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 8392 13880 8444 13932
rect 12164 13923 12216 13932
rect 7104 13855 7156 13864
rect 7104 13821 7127 13855
rect 7127 13821 7156 13855
rect 7104 13812 7156 13821
rect 9772 13812 9824 13864
rect 11888 13855 11940 13864
rect 11888 13821 11897 13855
rect 11897 13821 11931 13855
rect 11931 13821 11940 13855
rect 11888 13812 11940 13821
rect 12164 13889 12173 13923
rect 12173 13889 12207 13923
rect 12207 13889 12216 13923
rect 12164 13880 12216 13889
rect 14004 13923 14056 13932
rect 14004 13889 14013 13923
rect 14013 13889 14047 13923
rect 14047 13889 14056 13923
rect 14004 13880 14056 13889
rect 16948 13923 17000 13932
rect 16948 13889 16957 13923
rect 16957 13889 16991 13923
rect 16991 13889 17000 13923
rect 16948 13880 17000 13889
rect 20352 14016 20404 14068
rect 20996 14059 21048 14068
rect 20996 14025 21005 14059
rect 21005 14025 21039 14059
rect 21039 14025 21048 14059
rect 20996 14016 21048 14025
rect 21824 14059 21876 14068
rect 21824 14025 21833 14059
rect 21833 14025 21867 14059
rect 21867 14025 21876 14059
rect 21824 14016 21876 14025
rect 22100 14059 22152 14068
rect 22100 14025 22109 14059
rect 22109 14025 22143 14059
rect 22143 14025 22152 14059
rect 23112 14059 23164 14068
rect 22100 14016 22152 14025
rect 23112 14025 23121 14059
rect 23121 14025 23155 14059
rect 23155 14025 23164 14059
rect 23112 14016 23164 14025
rect 23480 14059 23532 14068
rect 23480 14025 23489 14059
rect 23489 14025 23523 14059
rect 23523 14025 23532 14059
rect 23480 14016 23532 14025
rect 21916 13948 21968 14000
rect 12440 13812 12492 13864
rect 9128 13744 9180 13796
rect 11244 13787 11296 13796
rect 11244 13753 11253 13787
rect 11253 13753 11287 13787
rect 11287 13753 11296 13787
rect 11244 13744 11296 13753
rect 12256 13744 12308 13796
rect 14372 13855 14424 13864
rect 14372 13821 14381 13855
rect 14381 13821 14415 13855
rect 14415 13821 14424 13855
rect 14372 13812 14424 13821
rect 14648 13855 14700 13864
rect 14648 13821 14682 13855
rect 14682 13821 14700 13855
rect 14648 13812 14700 13821
rect 17408 13812 17460 13864
rect 17868 13812 17920 13864
rect 19248 13880 19300 13932
rect 19616 13880 19668 13932
rect 12624 13744 12676 13796
rect 18604 13744 18656 13796
rect 20260 13812 20312 13864
rect 22008 13812 22060 13864
rect 23388 13812 23440 13864
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 19340 13744 19392 13796
rect 3240 13676 3292 13728
rect 4436 13676 4488 13728
rect 5172 13676 5224 13728
rect 8484 13676 8536 13728
rect 11980 13676 12032 13728
rect 12532 13676 12584 13728
rect 13820 13719 13872 13728
rect 13820 13685 13829 13719
rect 13829 13685 13863 13719
rect 13863 13685 13872 13719
rect 13820 13676 13872 13685
rect 18236 13676 18288 13728
rect 18696 13676 18748 13728
rect 25044 13719 25096 13728
rect 25044 13685 25053 13719
rect 25053 13685 25087 13719
rect 25087 13685 25096 13719
rect 25044 13676 25096 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1768 13472 1820 13524
rect 2596 13472 2648 13524
rect 3792 13472 3844 13524
rect 4896 13472 4948 13524
rect 5172 13515 5224 13524
rect 5172 13481 5181 13515
rect 5181 13481 5215 13515
rect 5215 13481 5224 13515
rect 5172 13472 5224 13481
rect 5632 13515 5684 13524
rect 5632 13481 5641 13515
rect 5641 13481 5675 13515
rect 5675 13481 5684 13515
rect 5632 13472 5684 13481
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 9128 13515 9180 13524
rect 9128 13481 9137 13515
rect 9137 13481 9171 13515
rect 9171 13481 9180 13515
rect 9128 13472 9180 13481
rect 9772 13472 9824 13524
rect 2688 13404 2740 13456
rect 3884 13447 3936 13456
rect 3884 13413 3893 13447
rect 3893 13413 3927 13447
rect 3927 13413 3936 13447
rect 3884 13404 3936 13413
rect 3976 13404 4028 13456
rect 4252 13404 4304 13456
rect 2504 13336 2556 13388
rect 6828 13404 6880 13456
rect 8024 13404 8076 13456
rect 10692 13472 10744 13524
rect 11980 13472 12032 13524
rect 12624 13515 12676 13524
rect 12624 13481 12633 13515
rect 12633 13481 12667 13515
rect 12667 13481 12676 13515
rect 12624 13472 12676 13481
rect 6000 13379 6052 13388
rect 6000 13345 6034 13379
rect 6034 13345 6052 13379
rect 6000 13336 6052 13345
rect 12440 13336 12492 13388
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 4160 13268 4212 13320
rect 4896 13268 4948 13320
rect 8300 13268 8352 13320
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 10140 13311 10192 13320
rect 8484 13268 8536 13277
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 4068 13243 4120 13252
rect 4068 13209 4077 13243
rect 4077 13209 4111 13243
rect 4111 13209 4120 13243
rect 4068 13200 4120 13209
rect 6828 13200 6880 13252
rect 7840 13243 7892 13252
rect 7840 13209 7849 13243
rect 7849 13209 7883 13243
rect 7883 13209 7892 13243
rect 7840 13200 7892 13209
rect 9772 13200 9824 13252
rect 10048 13200 10100 13252
rect 12624 13268 12676 13320
rect 15936 13472 15988 13524
rect 16488 13472 16540 13524
rect 16764 13515 16816 13524
rect 16764 13481 16773 13515
rect 16773 13481 16807 13515
rect 16807 13481 16816 13515
rect 16764 13472 16816 13481
rect 16856 13515 16908 13524
rect 16856 13481 16865 13515
rect 16865 13481 16899 13515
rect 16899 13481 16908 13515
rect 17408 13515 17460 13524
rect 16856 13472 16908 13481
rect 17408 13481 17417 13515
rect 17417 13481 17451 13515
rect 17451 13481 17460 13515
rect 17408 13472 17460 13481
rect 18236 13515 18288 13524
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 18328 13472 18380 13524
rect 18696 13472 18748 13524
rect 20628 13472 20680 13524
rect 21640 13515 21692 13524
rect 21640 13481 21649 13515
rect 21649 13481 21683 13515
rect 21683 13481 21692 13515
rect 21640 13472 21692 13481
rect 23204 13472 23256 13524
rect 23296 13472 23348 13524
rect 23664 13515 23716 13524
rect 23664 13481 23673 13515
rect 23673 13481 23707 13515
rect 23707 13481 23716 13515
rect 23664 13472 23716 13481
rect 24860 13515 24912 13524
rect 24860 13481 24869 13515
rect 24869 13481 24903 13515
rect 24903 13481 24912 13515
rect 24860 13472 24912 13481
rect 26056 13472 26108 13524
rect 14280 13404 14332 13456
rect 14556 13404 14608 13456
rect 15752 13404 15804 13456
rect 18052 13379 18104 13388
rect 18052 13345 18061 13379
rect 18061 13345 18095 13379
rect 18095 13345 18104 13379
rect 18052 13336 18104 13345
rect 18420 13336 18472 13388
rect 20536 13379 20588 13388
rect 20536 13345 20545 13379
rect 20545 13345 20579 13379
rect 20579 13345 20588 13379
rect 20536 13336 20588 13345
rect 21916 13336 21968 13388
rect 22560 13379 22612 13388
rect 22560 13345 22569 13379
rect 22569 13345 22603 13379
rect 22603 13345 22612 13379
rect 22560 13336 22612 13345
rect 22652 13336 22704 13388
rect 23204 13336 23256 13388
rect 24032 13379 24084 13388
rect 24032 13345 24041 13379
rect 24041 13345 24075 13379
rect 24075 13345 24084 13379
rect 24032 13336 24084 13345
rect 25320 13379 25372 13388
rect 25320 13345 25329 13379
rect 25329 13345 25363 13379
rect 25363 13345 25372 13379
rect 25320 13336 25372 13345
rect 13820 13200 13872 13252
rect 1952 13175 2004 13184
rect 1952 13141 1961 13175
rect 1961 13141 1995 13175
rect 1995 13141 2004 13175
rect 1952 13132 2004 13141
rect 3608 13132 3660 13184
rect 7932 13175 7984 13184
rect 7932 13141 7941 13175
rect 7941 13141 7975 13175
rect 7975 13141 7984 13175
rect 7932 13132 7984 13141
rect 11152 13132 11204 13184
rect 12256 13175 12308 13184
rect 12256 13141 12265 13175
rect 12265 13141 12299 13175
rect 12299 13141 12308 13175
rect 12256 13132 12308 13141
rect 14556 13132 14608 13184
rect 15844 13311 15896 13320
rect 15844 13277 15853 13311
rect 15853 13277 15887 13311
rect 15887 13277 15896 13311
rect 18696 13311 18748 13320
rect 15844 13268 15896 13277
rect 18696 13277 18705 13311
rect 18705 13277 18739 13311
rect 18739 13277 18748 13311
rect 18696 13268 18748 13277
rect 19156 13268 19208 13320
rect 24216 13311 24268 13320
rect 24216 13277 24225 13311
rect 24225 13277 24259 13311
rect 24259 13277 24268 13311
rect 24216 13268 24268 13277
rect 17776 13200 17828 13252
rect 18236 13200 18288 13252
rect 19892 13200 19944 13252
rect 19340 13132 19392 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 2780 12928 2832 12980
rect 6000 12928 6052 12980
rect 6092 12928 6144 12980
rect 8024 12971 8076 12980
rect 8024 12937 8033 12971
rect 8033 12937 8067 12971
rect 8067 12937 8076 12971
rect 8024 12928 8076 12937
rect 10232 12928 10284 12980
rect 10692 12928 10744 12980
rect 2964 12860 3016 12912
rect 3056 12792 3108 12844
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 4252 12792 4304 12844
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 8300 12860 8352 12912
rect 10140 12860 10192 12912
rect 4896 12792 4948 12844
rect 8668 12835 8720 12844
rect 1492 12724 1544 12776
rect 4068 12724 4120 12776
rect 7288 12767 7340 12776
rect 7288 12733 7297 12767
rect 7297 12733 7331 12767
rect 7331 12733 7340 12767
rect 7288 12724 7340 12733
rect 7748 12724 7800 12776
rect 1952 12656 2004 12708
rect 7196 12699 7248 12708
rect 7196 12665 7205 12699
rect 7205 12665 7239 12699
rect 7239 12665 7248 12699
rect 7196 12656 7248 12665
rect 8668 12801 8677 12835
rect 8677 12801 8711 12835
rect 8711 12801 8720 12835
rect 8668 12792 8720 12801
rect 11244 12792 11296 12844
rect 14372 12928 14424 12980
rect 16120 12928 16172 12980
rect 18328 12928 18380 12980
rect 18696 12928 18748 12980
rect 18880 12971 18932 12980
rect 18880 12937 18889 12971
rect 18889 12937 18923 12971
rect 18923 12937 18932 12971
rect 18880 12928 18932 12937
rect 19892 12971 19944 12980
rect 19892 12937 19901 12971
rect 19901 12937 19935 12971
rect 19935 12937 19944 12971
rect 19892 12928 19944 12937
rect 21272 12971 21324 12980
rect 21272 12937 21281 12971
rect 21281 12937 21315 12971
rect 21315 12937 21324 12971
rect 21272 12928 21324 12937
rect 22652 12971 22704 12980
rect 22652 12937 22661 12971
rect 22661 12937 22695 12971
rect 22695 12937 22704 12971
rect 22652 12928 22704 12937
rect 22836 12928 22888 12980
rect 19156 12860 19208 12912
rect 19248 12860 19300 12912
rect 21180 12860 21232 12912
rect 22560 12860 22612 12912
rect 15844 12792 15896 12844
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 8576 12767 8628 12776
rect 8576 12733 8585 12767
rect 8585 12733 8619 12767
rect 8619 12733 8628 12767
rect 8576 12724 8628 12733
rect 9588 12724 9640 12776
rect 13268 12767 13320 12776
rect 10968 12656 11020 12708
rect 11336 12656 11388 12708
rect 2504 12588 2556 12640
rect 3148 12631 3200 12640
rect 3148 12597 3157 12631
rect 3157 12597 3191 12631
rect 3191 12597 3200 12631
rect 3148 12588 3200 12597
rect 7840 12588 7892 12640
rect 9956 12588 10008 12640
rect 11060 12588 11112 12640
rect 13268 12733 13302 12767
rect 13302 12733 13320 12767
rect 13268 12724 13320 12733
rect 21272 12724 21324 12776
rect 21916 12767 21968 12776
rect 21916 12733 21925 12767
rect 21925 12733 21959 12767
rect 21959 12733 21968 12767
rect 21916 12724 21968 12733
rect 22836 12724 22888 12776
rect 23112 12724 23164 12776
rect 23664 12767 23716 12776
rect 23664 12733 23673 12767
rect 23673 12733 23707 12767
rect 23707 12733 23716 12767
rect 23664 12724 23716 12733
rect 25044 12724 25096 12776
rect 16120 12656 16172 12708
rect 18512 12656 18564 12708
rect 11520 12588 11572 12640
rect 12440 12588 12492 12640
rect 13544 12588 13596 12640
rect 15660 12631 15712 12640
rect 15660 12597 15669 12631
rect 15669 12597 15703 12631
rect 15703 12597 15712 12631
rect 15660 12588 15712 12597
rect 18696 12631 18748 12640
rect 18696 12597 18705 12631
rect 18705 12597 18739 12631
rect 18739 12597 18748 12631
rect 18696 12588 18748 12597
rect 19064 12588 19116 12640
rect 25136 12588 25188 12640
rect 25320 12631 25372 12640
rect 25320 12597 25329 12631
rect 25329 12597 25363 12631
rect 25363 12597 25372 12631
rect 25320 12588 25372 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1492 12384 1544 12436
rect 1952 12384 2004 12436
rect 4068 12427 4120 12436
rect 4068 12393 4077 12427
rect 4077 12393 4111 12427
rect 4111 12393 4120 12427
rect 4068 12384 4120 12393
rect 4344 12384 4396 12436
rect 5172 12427 5224 12436
rect 5172 12393 5181 12427
rect 5181 12393 5215 12427
rect 5215 12393 5224 12427
rect 5172 12384 5224 12393
rect 6828 12384 6880 12436
rect 7288 12384 7340 12436
rect 8208 12384 8260 12436
rect 8484 12384 8536 12436
rect 8576 12384 8628 12436
rect 10048 12384 10100 12436
rect 12256 12384 12308 12436
rect 12992 12427 13044 12436
rect 12992 12393 13001 12427
rect 13001 12393 13035 12427
rect 13035 12393 13044 12427
rect 12992 12384 13044 12393
rect 14740 12384 14792 12436
rect 2044 12316 2096 12368
rect 10692 12316 10744 12368
rect 11152 12316 11204 12368
rect 15752 12384 15804 12436
rect 18052 12384 18104 12436
rect 18880 12384 18932 12436
rect 19524 12427 19576 12436
rect 19524 12393 19533 12427
rect 19533 12393 19567 12427
rect 19567 12393 19576 12427
rect 19524 12384 19576 12393
rect 21732 12384 21784 12436
rect 23204 12384 23256 12436
rect 23296 12384 23348 12436
rect 23480 12384 23532 12436
rect 24216 12384 24268 12436
rect 24676 12384 24728 12436
rect 2136 12248 2188 12300
rect 2872 12291 2924 12300
rect 2872 12257 2881 12291
rect 2881 12257 2915 12291
rect 2915 12257 2924 12291
rect 2872 12248 2924 12257
rect 4620 12248 4672 12300
rect 11060 12248 11112 12300
rect 11428 12248 11480 12300
rect 13360 12291 13412 12300
rect 13360 12257 13369 12291
rect 13369 12257 13403 12291
rect 13403 12257 13412 12291
rect 13360 12248 13412 12257
rect 13728 12248 13780 12300
rect 14280 12248 14332 12300
rect 15292 12248 15344 12300
rect 15568 12248 15620 12300
rect 19340 12316 19392 12368
rect 23112 12316 23164 12368
rect 3608 12180 3660 12232
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 13544 12223 13596 12232
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 15752 12223 15804 12232
rect 13544 12180 13596 12189
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 17500 12248 17552 12300
rect 19156 12291 19208 12300
rect 19156 12257 19165 12291
rect 19165 12257 19199 12291
rect 19199 12257 19208 12291
rect 19156 12248 19208 12257
rect 21640 12291 21692 12300
rect 21640 12257 21649 12291
rect 21649 12257 21683 12291
rect 21683 12257 21692 12291
rect 21640 12248 21692 12257
rect 23020 12248 23072 12300
rect 24124 12316 24176 12368
rect 24860 12248 24912 12300
rect 16304 12223 16356 12232
rect 16304 12189 16313 12223
rect 16313 12189 16347 12223
rect 16347 12189 16356 12223
rect 16304 12180 16356 12189
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 17408 12223 17460 12232
rect 17408 12189 17417 12223
rect 17417 12189 17451 12223
rect 17451 12189 17460 12223
rect 17408 12180 17460 12189
rect 18512 12180 18564 12232
rect 19248 12180 19300 12232
rect 19800 12223 19852 12232
rect 19800 12189 19809 12223
rect 19809 12189 19843 12223
rect 19843 12189 19852 12223
rect 19800 12180 19852 12189
rect 23940 12180 23992 12232
rect 24124 12180 24176 12232
rect 24400 12180 24452 12232
rect 24676 12180 24728 12232
rect 3148 12112 3200 12164
rect 4896 12112 4948 12164
rect 11336 12112 11388 12164
rect 12072 12112 12124 12164
rect 13268 12112 13320 12164
rect 24032 12112 24084 12164
rect 13452 12044 13504 12096
rect 14096 12087 14148 12096
rect 14096 12053 14105 12087
rect 14105 12053 14139 12087
rect 14139 12053 14148 12087
rect 14096 12044 14148 12053
rect 14372 12044 14424 12096
rect 16856 12087 16908 12096
rect 16856 12053 16865 12087
rect 16865 12053 16899 12087
rect 16899 12053 16908 12087
rect 16856 12044 16908 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1400 11840 1452 11892
rect 2044 11883 2096 11892
rect 2044 11849 2053 11883
rect 2053 11849 2087 11883
rect 2087 11849 2096 11883
rect 2044 11840 2096 11849
rect 2136 11840 2188 11892
rect 3148 11840 3200 11892
rect 4344 11840 4396 11892
rect 4712 11840 4764 11892
rect 11152 11883 11204 11892
rect 11152 11849 11161 11883
rect 11161 11849 11195 11883
rect 11195 11849 11204 11883
rect 11152 11840 11204 11849
rect 11980 11840 12032 11892
rect 12624 11840 12676 11892
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 16120 11883 16172 11892
rect 16120 11849 16129 11883
rect 16129 11849 16163 11883
rect 16163 11849 16172 11883
rect 16120 11840 16172 11849
rect 17316 11840 17368 11892
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 18236 11883 18288 11892
rect 18236 11849 18245 11883
rect 18245 11849 18279 11883
rect 18279 11849 18288 11883
rect 18236 11840 18288 11849
rect 21640 11840 21692 11892
rect 22284 11840 22336 11892
rect 23020 11883 23072 11892
rect 23020 11849 23029 11883
rect 23029 11849 23063 11883
rect 23063 11849 23072 11883
rect 23020 11840 23072 11849
rect 24860 11840 24912 11892
rect 25044 11883 25096 11892
rect 25044 11849 25053 11883
rect 25053 11849 25087 11883
rect 25087 11849 25096 11883
rect 25044 11840 25096 11849
rect 4620 11772 4672 11824
rect 11060 11772 11112 11824
rect 13360 11772 13412 11824
rect 16304 11772 16356 11824
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 3608 11704 3660 11713
rect 11244 11704 11296 11756
rect 12348 11704 12400 11756
rect 13544 11704 13596 11756
rect 14740 11704 14792 11756
rect 16488 11704 16540 11756
rect 21456 11747 21508 11756
rect 21456 11713 21465 11747
rect 21465 11713 21499 11747
rect 21499 11713 21508 11747
rect 21456 11704 21508 11713
rect 22284 11747 22336 11756
rect 22284 11713 22293 11747
rect 22293 11713 22327 11747
rect 22327 11713 22336 11747
rect 22284 11704 22336 11713
rect 1676 11636 1728 11688
rect 2412 11636 2464 11688
rect 3148 11636 3200 11688
rect 3516 11636 3568 11688
rect 13728 11679 13780 11688
rect 13728 11645 13737 11679
rect 13737 11645 13771 11679
rect 13771 11645 13780 11679
rect 13728 11636 13780 11645
rect 23848 11704 23900 11756
rect 24032 11704 24084 11756
rect 24952 11704 25004 11756
rect 14740 11568 14792 11620
rect 15752 11568 15804 11620
rect 3240 11500 3292 11552
rect 3976 11500 4028 11552
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 13452 11500 13504 11552
rect 14372 11543 14424 11552
rect 14372 11509 14381 11543
rect 14381 11509 14415 11543
rect 14415 11509 14424 11543
rect 14372 11500 14424 11509
rect 16396 11500 16448 11552
rect 23848 11543 23900 11552
rect 23848 11509 23857 11543
rect 23857 11509 23891 11543
rect 23891 11509 23900 11543
rect 23848 11500 23900 11509
rect 24124 11568 24176 11620
rect 24492 11543 24544 11552
rect 24492 11509 24501 11543
rect 24501 11509 24535 11543
rect 24535 11509 24544 11543
rect 24492 11500 24544 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2596 11296 2648 11348
rect 3148 11339 3200 11348
rect 3148 11305 3157 11339
rect 3157 11305 3191 11339
rect 3191 11305 3200 11339
rect 3148 11296 3200 11305
rect 3608 11296 3660 11348
rect 11428 11339 11480 11348
rect 11428 11305 11437 11339
rect 11437 11305 11471 11339
rect 11471 11305 11480 11339
rect 11428 11296 11480 11305
rect 12348 11339 12400 11348
rect 12348 11305 12357 11339
rect 12357 11305 12391 11339
rect 12391 11305 12400 11339
rect 12348 11296 12400 11305
rect 12532 11296 12584 11348
rect 15660 11296 15712 11348
rect 16488 11296 16540 11348
rect 16948 11296 17000 11348
rect 22744 11296 22796 11348
rect 13084 11228 13136 11280
rect 13452 11228 13504 11280
rect 15568 11228 15620 11280
rect 16120 11228 16172 11280
rect 16856 11228 16908 11280
rect 24676 11296 24728 11348
rect 26332 11228 26384 11280
rect 14740 11160 14792 11212
rect 15384 11160 15436 11212
rect 16028 11160 16080 11212
rect 22376 11203 22428 11212
rect 22376 11169 22385 11203
rect 22385 11169 22419 11203
rect 22419 11169 22428 11203
rect 22376 11160 22428 11169
rect 23480 11203 23532 11212
rect 23480 11169 23489 11203
rect 23489 11169 23523 11203
rect 23523 11169 23532 11203
rect 23480 11160 23532 11169
rect 24584 11203 24636 11212
rect 24584 11169 24593 11203
rect 24593 11169 24627 11203
rect 24627 11169 24636 11203
rect 24584 11160 24636 11169
rect 24860 11160 24912 11212
rect 13176 11092 13228 11144
rect 13728 11092 13780 11144
rect 15752 11092 15804 11144
rect 16304 11092 16356 11144
rect 24124 11135 24176 11144
rect 24124 11101 24133 11135
rect 24133 11101 24167 11135
rect 24167 11101 24176 11135
rect 24124 11092 24176 11101
rect 24492 11092 24544 11144
rect 14096 11024 14148 11076
rect 14648 11024 14700 11076
rect 16856 11067 16908 11076
rect 16856 11033 16865 11067
rect 16865 11033 16899 11067
rect 16899 11033 16908 11067
rect 16856 11024 16908 11033
rect 17408 11024 17460 11076
rect 23756 11024 23808 11076
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2504 10795 2556 10804
rect 2504 10761 2513 10795
rect 2513 10761 2547 10795
rect 2547 10761 2556 10795
rect 2504 10752 2556 10761
rect 13728 10795 13780 10804
rect 13728 10761 13737 10795
rect 13737 10761 13771 10795
rect 13771 10761 13780 10795
rect 13728 10752 13780 10761
rect 15384 10795 15436 10804
rect 15384 10761 15393 10795
rect 15393 10761 15427 10795
rect 15427 10761 15436 10795
rect 15384 10752 15436 10761
rect 15752 10795 15804 10804
rect 15752 10761 15761 10795
rect 15761 10761 15795 10795
rect 15795 10761 15804 10795
rect 15752 10752 15804 10761
rect 16120 10795 16172 10804
rect 16120 10761 16129 10795
rect 16129 10761 16163 10795
rect 16163 10761 16172 10795
rect 16120 10752 16172 10761
rect 22376 10795 22428 10804
rect 22376 10761 22385 10795
rect 22385 10761 22419 10795
rect 22419 10761 22428 10795
rect 22376 10752 22428 10761
rect 23480 10752 23532 10804
rect 23940 10752 23992 10804
rect 24860 10752 24912 10804
rect 25780 10752 25832 10804
rect 24400 10659 24452 10668
rect 24400 10625 24409 10659
rect 24409 10625 24443 10659
rect 24443 10625 24452 10659
rect 24400 10616 24452 10625
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 13084 10455 13136 10464
rect 13084 10421 13093 10455
rect 13093 10421 13127 10455
rect 13127 10421 13136 10455
rect 13084 10412 13136 10421
rect 13452 10455 13504 10464
rect 13452 10421 13461 10455
rect 13461 10421 13495 10455
rect 13495 10421 13504 10455
rect 13452 10412 13504 10421
rect 14648 10455 14700 10464
rect 14648 10421 14657 10455
rect 14657 10421 14691 10455
rect 14691 10421 14700 10455
rect 14648 10412 14700 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 24768 10251 24820 10260
rect 24768 10217 24777 10251
rect 24777 10217 24811 10251
rect 24811 10217 24820 10251
rect 24768 10208 24820 10217
rect 24676 10072 24728 10124
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 24216 9596 24268 9648
rect 25136 9503 25188 9512
rect 25136 9469 25145 9503
rect 25145 9469 25179 9503
rect 25179 9469 25188 9503
rect 25136 9460 25188 9469
rect 19340 9392 19392 9444
rect 25964 9392 26016 9444
rect 24032 9324 24084 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 9588 8576 9640 8628
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 9588 5856 9640 5908
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1400 5312 1452 5364
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 572 2796 624 2848
rect 3332 2796 3384 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 14096 2635 14148 2644
rect 14096 2601 14105 2635
rect 14105 2601 14139 2635
rect 14139 2601 14148 2635
rect 14096 2592 14148 2601
rect 12716 2499 12768 2508
rect 12716 2465 12725 2499
rect 12725 2465 12759 2499
rect 12759 2465 12768 2499
rect 12716 2456 12768 2465
rect 25136 2252 25188 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 3054 27520 3110 28000
rect 3514 27704 3570 27713
rect 3514 27639 3570 27648
rect 308 25226 336 27520
rect 860 27418 888 27520
rect 768 27390 888 27418
rect 296 25220 348 25226
rect 296 25162 348 25168
rect 768 16017 796 27390
rect 1412 24188 1440 27520
rect 1964 25770 1992 27520
rect 1952 25764 2004 25770
rect 1952 25706 2004 25712
rect 2320 25356 2372 25362
rect 2320 25298 2372 25304
rect 1584 25152 1636 25158
rect 1584 25094 1636 25100
rect 1596 24721 1624 25094
rect 2332 24750 2360 25298
rect 2516 24993 2544 27520
rect 2778 25936 2834 25945
rect 2778 25871 2834 25880
rect 2792 25498 2820 25871
rect 2780 25492 2832 25498
rect 2780 25434 2832 25440
rect 2596 25356 2648 25362
rect 2596 25298 2648 25304
rect 2502 24984 2558 24993
rect 2502 24919 2558 24928
rect 2608 24834 2636 25298
rect 2686 25256 2742 25265
rect 2686 25191 2742 25200
rect 2700 24954 2728 25191
rect 2688 24948 2740 24954
rect 2688 24890 2740 24896
rect 2608 24806 2728 24834
rect 2320 24744 2372 24750
rect 1582 24712 1638 24721
rect 2320 24686 2372 24692
rect 1582 24647 1638 24656
rect 1584 24608 1636 24614
rect 1584 24550 1636 24556
rect 1412 24160 1532 24188
rect 1400 24064 1452 24070
rect 1400 24006 1452 24012
rect 1412 21049 1440 24006
rect 1504 22001 1532 24160
rect 1596 22273 1624 24550
rect 1768 24268 1820 24274
rect 1768 24210 1820 24216
rect 1780 24070 1808 24210
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1676 23520 1728 23526
rect 1676 23462 1728 23468
rect 1582 22264 1638 22273
rect 1582 22199 1638 22208
rect 1490 21992 1546 22001
rect 1490 21927 1546 21936
rect 1492 21888 1544 21894
rect 1492 21830 1544 21836
rect 1504 21486 1532 21830
rect 1492 21480 1544 21486
rect 1492 21422 1544 21428
rect 1504 21146 1532 21422
rect 1492 21140 1544 21146
rect 1492 21082 1544 21088
rect 1398 21040 1454 21049
rect 1398 20975 1454 20984
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 18970 1440 20878
rect 1688 20369 1716 23462
rect 1780 21554 1808 24006
rect 2136 23860 2188 23866
rect 2136 23802 2188 23808
rect 1952 23520 2004 23526
rect 1952 23462 2004 23468
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1674 20360 1730 20369
rect 1674 20295 1730 20304
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 19825 1624 20198
rect 1582 19816 1638 19825
rect 1582 19751 1638 19760
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1872 19378 1900 19654
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1676 19168 1728 19174
rect 1676 19110 1728 19116
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1412 18426 1440 18906
rect 1400 18420 1452 18426
rect 1400 18362 1452 18368
rect 1688 17542 1716 19110
rect 1872 18630 1900 19314
rect 1964 19281 1992 23462
rect 2148 22574 2176 23802
rect 2226 23624 2282 23633
rect 2226 23559 2282 23568
rect 2240 23254 2268 23559
rect 2228 23248 2280 23254
rect 2228 23190 2280 23196
rect 2240 22778 2268 23190
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 2136 22568 2188 22574
rect 2136 22510 2188 22516
rect 2044 20256 2096 20262
rect 2042 20224 2044 20233
rect 2096 20224 2098 20233
rect 2042 20159 2098 20168
rect 2228 19304 2280 19310
rect 1950 19272 2006 19281
rect 2228 19246 2280 19252
rect 1950 19207 2006 19216
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 1860 18624 1912 18630
rect 1860 18566 1912 18572
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1780 17746 1808 18158
rect 1872 17746 1900 18566
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1688 17105 1716 17478
rect 1674 17096 1730 17105
rect 1964 17082 1992 18566
rect 2056 18086 2084 18702
rect 2240 18630 2268 19246
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 1674 17031 1730 17040
rect 1780 17054 1992 17082
rect 1582 16688 1638 16697
rect 1780 16658 1808 17054
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1858 16688 1914 16697
rect 1582 16623 1638 16632
rect 1768 16652 1820 16658
rect 1398 16144 1454 16153
rect 1398 16079 1454 16088
rect 754 16008 810 16017
rect 754 15943 810 15952
rect 1412 11898 1440 16079
rect 1492 15972 1544 15978
rect 1492 15914 1544 15920
rect 1504 12782 1532 15914
rect 1596 12986 1624 16623
rect 1858 16623 1914 16632
rect 1768 16594 1820 16600
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1780 16046 1808 16390
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1688 15201 1716 15302
rect 1674 15192 1730 15201
rect 1674 15127 1730 15136
rect 1688 15026 1716 15127
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1676 14884 1728 14890
rect 1676 14826 1728 14832
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1504 12442 1532 12718
rect 1492 12436 1544 12442
rect 1492 12378 1544 12384
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 1688 11694 1716 14826
rect 1780 13530 1808 15982
rect 1872 13938 1900 16623
rect 1964 14346 1992 16934
rect 2056 16538 2084 18022
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 2240 16794 2268 16934
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2228 16584 2280 16590
rect 2056 16510 2176 16538
rect 2228 16526 2280 16532
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1964 13870 1992 14282
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1964 12714 1992 13126
rect 1952 12708 2004 12714
rect 1952 12650 2004 12656
rect 1964 12442 1992 12650
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 2056 12374 2084 14350
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 2056 11898 2084 12310
rect 2148 12306 2176 16510
rect 2240 15706 2268 16526
rect 2332 16289 2360 24686
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2424 23361 2452 24550
rect 2594 24440 2650 24449
rect 2594 24375 2650 24384
rect 2504 23656 2556 23662
rect 2504 23598 2556 23604
rect 2410 23352 2466 23361
rect 2410 23287 2466 23296
rect 2516 22273 2544 23598
rect 2608 23322 2636 24375
rect 2700 24154 2728 24806
rect 2780 24200 2832 24206
rect 2700 24148 2780 24154
rect 3068 24177 3096 27520
rect 3528 27334 3556 27639
rect 3606 27520 3662 28000
rect 4158 27520 4214 28000
rect 4710 27520 4766 28000
rect 5262 27520 5318 28000
rect 5814 27520 5870 28000
rect 6366 27520 6422 28000
rect 6918 27520 6974 28000
rect 7562 27520 7618 28000
rect 8114 27520 8170 28000
rect 8666 27520 8722 28000
rect 9218 27520 9274 28000
rect 9770 27520 9826 28000
rect 10322 27520 10378 28000
rect 10874 27520 10930 28000
rect 11426 27520 11482 28000
rect 11978 27520 12034 28000
rect 12530 27520 12586 28000
rect 13082 27520 13138 28000
rect 13634 27520 13690 28000
rect 14278 27520 14334 28000
rect 14830 27520 14886 28000
rect 15382 27520 15438 28000
rect 15934 27520 15990 28000
rect 16486 27520 16542 28000
rect 17038 27520 17094 28000
rect 17590 27520 17646 28000
rect 18142 27520 18198 28000
rect 18694 27520 18750 28000
rect 19246 27520 19302 28000
rect 19798 27520 19854 28000
rect 20350 27520 20406 28000
rect 20902 27520 20958 28000
rect 21546 27520 21602 28000
rect 22098 27520 22154 28000
rect 22650 27520 22706 28000
rect 23202 27520 23258 28000
rect 23754 27520 23810 28000
rect 24306 27520 24362 28000
rect 24858 27520 24914 28000
rect 25410 27520 25466 28000
rect 25594 27704 25650 27713
rect 25594 27639 25650 27648
rect 3516 27328 3568 27334
rect 3516 27270 3568 27276
rect 3148 24744 3200 24750
rect 3148 24686 3200 24692
rect 2700 24142 2832 24148
rect 3054 24168 3110 24177
rect 2700 24126 2820 24142
rect 2700 23866 2728 24126
rect 3054 24103 3110 24112
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2688 23860 2740 23866
rect 2688 23802 2740 23808
rect 2688 23520 2740 23526
rect 2688 23462 2740 23468
rect 2596 23316 2648 23322
rect 2596 23258 2648 23264
rect 2608 22642 2636 23258
rect 2596 22636 2648 22642
rect 2596 22578 2648 22584
rect 2502 22264 2558 22273
rect 2502 22199 2558 22208
rect 2412 21888 2464 21894
rect 2412 21830 2464 21836
rect 2424 21729 2452 21830
rect 2410 21720 2466 21729
rect 2516 21690 2544 22199
rect 2596 22024 2648 22030
rect 2596 21966 2648 21972
rect 2410 21655 2466 21664
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 2608 21457 2636 21966
rect 2700 21593 2728 23462
rect 2792 22817 2820 24006
rect 2778 22808 2834 22817
rect 2778 22743 2834 22752
rect 2778 22264 2834 22273
rect 2778 22199 2780 22208
rect 2832 22199 2834 22208
rect 2780 22170 2832 22176
rect 2686 21584 2742 21593
rect 2686 21519 2742 21528
rect 2594 21448 2650 21457
rect 2594 21383 2650 21392
rect 2608 21010 2636 21383
rect 2872 21344 2924 21350
rect 2872 21286 2924 21292
rect 2884 21078 2912 21286
rect 2872 21072 2924 21078
rect 2872 21014 2924 21020
rect 2596 21004 2648 21010
rect 2596 20946 2648 20952
rect 2884 20942 2912 21014
rect 2872 20936 2924 20942
rect 3160 20913 3188 24686
rect 3238 24304 3294 24313
rect 3238 24239 3240 24248
rect 3292 24239 3294 24248
rect 3240 24210 3292 24216
rect 3252 23866 3280 24210
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3516 23520 3568 23526
rect 3516 23462 3568 23468
rect 3528 23254 3556 23462
rect 3516 23248 3568 23254
rect 3516 23190 3568 23196
rect 3330 22672 3386 22681
rect 3330 22607 3386 22616
rect 3238 21992 3294 22001
rect 3238 21927 3294 21936
rect 3146 20904 3202 20913
rect 2872 20878 2924 20884
rect 2504 20868 2556 20874
rect 2504 20810 2556 20816
rect 3068 20862 3146 20890
rect 2516 20602 2544 20810
rect 2504 20596 2556 20602
rect 2504 20538 2556 20544
rect 2412 20392 2464 20398
rect 2412 20334 2464 20340
rect 2424 18766 2452 20334
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2884 20058 2912 20198
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2792 19514 2820 19858
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2884 19718 2912 19790
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2884 19446 2912 19654
rect 2872 19440 2924 19446
rect 2872 19382 2924 19388
rect 2872 19236 2924 19242
rect 2872 19178 2924 19184
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 2502 18184 2558 18193
rect 2412 18148 2464 18154
rect 2502 18119 2558 18128
rect 2412 18090 2464 18096
rect 2424 16590 2452 18090
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2318 16280 2374 16289
rect 2424 16250 2452 16526
rect 2318 16215 2374 16224
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2412 15972 2464 15978
rect 2412 15914 2464 15920
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2424 15638 2452 15914
rect 2412 15632 2464 15638
rect 2412 15574 2464 15580
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 2228 15428 2280 15434
rect 2228 15370 2280 15376
rect 2240 14618 2268 15370
rect 2332 15162 2360 15506
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 2424 15094 2452 15574
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2148 11898 2176 12242
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2424 11694 2452 15030
rect 2516 14618 2544 18119
rect 2780 18080 2832 18086
rect 2700 18028 2780 18034
rect 2700 18022 2832 18028
rect 2700 18006 2820 18022
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2608 17270 2636 17682
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 2608 15502 2636 17206
rect 2700 17202 2728 18006
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2884 16726 2912 19178
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2976 18329 3004 19110
rect 2962 18320 3018 18329
rect 2962 18255 3018 18264
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2700 16096 2728 16186
rect 2780 16108 2832 16114
rect 2700 16068 2780 16096
rect 2780 16050 2832 16056
rect 2884 16046 2912 16662
rect 2976 16182 3004 17002
rect 3068 16658 3096 20862
rect 3146 20839 3202 20848
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3160 19990 3188 20402
rect 3148 19984 3200 19990
rect 3252 19961 3280 21927
rect 3148 19926 3200 19932
rect 3238 19952 3294 19961
rect 3160 19446 3188 19926
rect 3238 19887 3294 19896
rect 3148 19440 3200 19446
rect 3148 19382 3200 19388
rect 3148 18148 3200 18154
rect 3148 18090 3200 18096
rect 3160 17882 3188 18090
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3252 17134 3280 17478
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 3344 16946 3372 22607
rect 3516 22024 3568 22030
rect 3516 21966 3568 21972
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3436 19825 3464 21830
rect 3528 21418 3556 21966
rect 3516 21412 3568 21418
rect 3516 21354 3568 21360
rect 3528 21162 3556 21354
rect 3620 21321 3648 27520
rect 3790 27160 3846 27169
rect 3790 27095 3846 27104
rect 3804 24954 3832 27095
rect 4066 26480 4122 26489
rect 4066 26415 4122 26424
rect 4080 25650 4108 26415
rect 4172 25809 4200 27520
rect 4620 25968 4672 25974
rect 4620 25910 4672 25916
rect 4158 25800 4214 25809
rect 4158 25735 4214 25744
rect 4080 25622 4200 25650
rect 3792 24948 3844 24954
rect 3792 24890 3844 24896
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 3606 21312 3662 21321
rect 3606 21247 3662 21256
rect 3528 21134 3648 21162
rect 3620 21078 3648 21134
rect 3608 21072 3660 21078
rect 3608 21014 3660 21020
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3528 20058 3556 20742
rect 3620 20505 3648 21014
rect 3606 20496 3662 20505
rect 3606 20431 3608 20440
rect 3660 20431 3662 20440
rect 3608 20402 3660 20408
rect 3620 20371 3648 20402
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3620 19938 3648 20198
rect 3528 19910 3648 19938
rect 3422 19816 3478 19825
rect 3422 19751 3478 19760
rect 3436 19242 3464 19751
rect 3528 19378 3556 19910
rect 3712 19718 3740 24550
rect 4172 24410 4200 25622
rect 4344 25356 4396 25362
rect 4344 25298 4396 25304
rect 4356 24750 4384 25298
rect 4344 24744 4396 24750
rect 4344 24686 4396 24692
rect 4252 24608 4304 24614
rect 4252 24550 4304 24556
rect 4160 24404 4212 24410
rect 4160 24346 4212 24352
rect 3790 24032 3846 24041
rect 3790 23967 3846 23976
rect 3804 23866 3832 23967
rect 3792 23860 3844 23866
rect 3792 23802 3844 23808
rect 4066 23488 4122 23497
rect 4066 23423 4122 23432
rect 4080 23322 4108 23423
rect 4068 23316 4120 23322
rect 4068 23258 4120 23264
rect 3976 23248 4028 23254
rect 3976 23190 4028 23196
rect 3884 23044 3936 23050
rect 3884 22986 3936 22992
rect 3896 22001 3924 22986
rect 3988 22574 4016 23190
rect 3976 22568 4028 22574
rect 3976 22510 4028 22516
rect 3988 22030 4016 22510
rect 4160 22500 4212 22506
rect 4160 22442 4212 22448
rect 4068 22432 4120 22438
rect 4068 22374 4120 22380
rect 4080 22166 4108 22374
rect 4068 22160 4120 22166
rect 4068 22102 4120 22108
rect 3976 22024 4028 22030
rect 3882 21992 3938 22001
rect 3976 21966 4028 21972
rect 3882 21927 3938 21936
rect 3792 21888 3844 21894
rect 3792 21830 3844 21836
rect 3700 19712 3752 19718
rect 3700 19654 3752 19660
rect 3698 19408 3754 19417
rect 3516 19372 3568 19378
rect 3698 19343 3754 19352
rect 3516 19314 3568 19320
rect 3424 19236 3476 19242
rect 3424 19178 3476 19184
rect 3528 18970 3556 19314
rect 3606 19136 3662 19145
rect 3606 19071 3662 19080
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3436 17649 3464 18566
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3422 17640 3478 17649
rect 3422 17575 3478 17584
rect 3252 16918 3372 16946
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 2964 16176 3016 16182
rect 2964 16118 3016 16124
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2792 15026 2820 15506
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 3068 14958 3096 15302
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 2964 14884 3016 14890
rect 2964 14826 3016 14832
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2792 14657 2820 14758
rect 2778 14648 2834 14657
rect 2504 14612 2556 14618
rect 2778 14583 2834 14592
rect 2504 14554 2556 14560
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 13546 2820 14418
rect 2976 13870 3004 14826
rect 3068 14074 3096 14894
rect 3252 14385 3280 16918
rect 3330 16824 3386 16833
rect 3330 16759 3386 16768
rect 3344 16726 3372 16759
rect 3332 16720 3384 16726
rect 3332 16662 3384 16668
rect 3344 15910 3372 16662
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3528 15552 3556 18158
rect 3620 17338 3648 19071
rect 3712 18222 3740 19343
rect 3804 19310 3832 21830
rect 3896 19666 3924 21927
rect 3988 21486 4016 21966
rect 4080 21622 4108 22102
rect 4172 21690 4200 22442
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 4068 21616 4120 21622
rect 4068 21558 4120 21564
rect 3976 21480 4028 21486
rect 3976 21422 4028 21428
rect 3988 20466 4016 21422
rect 4080 20942 4108 21558
rect 4160 21072 4212 21078
rect 4160 21014 4212 21020
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 4080 20602 4108 20878
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 4068 20052 4120 20058
rect 4172 20040 4200 21014
rect 4264 20369 4292 24550
rect 4356 24206 4384 24686
rect 4632 24274 4660 25910
rect 4724 24614 4752 27520
rect 4896 27328 4948 27334
rect 4896 27270 4948 27276
rect 4908 24954 4936 27270
rect 4896 24948 4948 24954
rect 4896 24890 4948 24896
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 5276 24426 5304 27520
rect 5828 25514 5856 27520
rect 5828 25486 6132 25514
rect 6000 25356 6052 25362
rect 6000 25298 6052 25304
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6012 24682 6040 25298
rect 6000 24676 6052 24682
rect 6000 24618 6052 24624
rect 5448 24608 5500 24614
rect 6104 24585 6132 25486
rect 6276 25152 6328 25158
rect 6276 25094 6328 25100
rect 5448 24550 5500 24556
rect 6090 24576 6146 24585
rect 4724 24398 5304 24426
rect 4620 24268 4672 24274
rect 4620 24210 4672 24216
rect 4344 24200 4396 24206
rect 4344 24142 4396 24148
rect 4632 23866 4660 24210
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 4528 23656 4580 23662
rect 4528 23598 4580 23604
rect 4540 20754 4568 23598
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 4632 20942 4660 21626
rect 4620 20936 4672 20942
rect 4620 20878 4672 20884
rect 4356 20726 4568 20754
rect 4250 20360 4306 20369
rect 4250 20295 4306 20304
rect 4120 20012 4200 20040
rect 4068 19994 4120 20000
rect 3896 19638 4200 19666
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 3792 19304 3844 19310
rect 3792 19246 3844 19252
rect 3804 18970 3832 19246
rect 3882 19136 3938 19145
rect 3882 19071 3938 19080
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 3700 18216 3752 18222
rect 3700 18158 3752 18164
rect 3792 18080 3844 18086
rect 3792 18022 3844 18028
rect 3698 17912 3754 17921
rect 3804 17882 3832 18022
rect 3698 17847 3754 17856
rect 3792 17876 3844 17882
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3712 16794 3740 17847
rect 3792 17818 3844 17824
rect 3896 17762 3924 19071
rect 3804 17734 3924 17762
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3608 16652 3660 16658
rect 3608 16594 3660 16600
rect 3436 15524 3556 15552
rect 3330 14648 3386 14657
rect 3330 14583 3386 14592
rect 3238 14376 3294 14385
rect 3238 14311 3294 14320
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2700 13518 2820 13546
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2516 12646 2544 13330
rect 2608 13002 2636 13466
rect 2700 13462 2728 13518
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2792 13297 2820 13518
rect 2964 13320 3016 13326
rect 2778 13288 2834 13297
rect 2964 13262 3016 13268
rect 2778 13223 2834 13232
rect 2608 12986 2820 13002
rect 2608 12980 2832 12986
rect 2608 12974 2780 12980
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 1688 11354 1716 11630
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 2516 10810 2544 12582
rect 2608 11354 2636 12974
rect 2780 12922 2832 12928
rect 2976 12918 3004 13262
rect 2964 12912 3016 12918
rect 2964 12854 3016 12860
rect 3068 12850 3096 14010
rect 3252 13734 3280 14214
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 1398 10704 1454 10713
rect 1398 10639 1454 10648
rect 1412 10606 1440 10639
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1582 10568 1638 10577
rect 1582 10503 1638 10512
rect 1596 10470 1624 10503
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1400 8424 1452 8430
rect 1398 8392 1400 8401
rect 1452 8392 1454 8401
rect 1398 8327 1454 8336
rect 1398 5808 1454 5817
rect 1398 5743 1400 5752
rect 1452 5743 1454 5752
rect 1400 5714 1452 5720
rect 1412 5370 1440 5714
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 2778 3496 2834 3505
rect 2778 3431 2834 3440
rect 572 2848 624 2854
rect 572 2790 624 2796
rect 584 2689 612 2790
rect 570 2680 626 2689
rect 570 2615 626 2624
rect 2792 480 2820 3431
rect 2884 3369 2912 12242
rect 3160 12170 3188 12582
rect 3148 12164 3200 12170
rect 3148 12106 3200 12112
rect 3160 11898 3188 12106
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3160 11354 3188 11630
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 2870 3360 2926 3369
rect 2870 3295 2926 3304
rect 3252 921 3280 11494
rect 3344 2854 3372 14583
rect 3436 13705 3464 15524
rect 3514 15464 3570 15473
rect 3514 15399 3570 15408
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 3422 13152 3478 13161
rect 3422 13087 3478 13096
rect 3436 12209 3464 13087
rect 3528 12753 3556 15399
rect 3620 14618 3648 16594
rect 3804 14929 3832 17734
rect 3884 15496 3936 15502
rect 3882 15464 3884 15473
rect 3936 15464 3938 15473
rect 3882 15399 3938 15408
rect 3790 14920 3846 14929
rect 3790 14855 3846 14864
rect 3882 14784 3938 14793
rect 3882 14719 3938 14728
rect 3896 14618 3924 14719
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3884 14340 3936 14346
rect 3884 14282 3936 14288
rect 3608 13796 3660 13802
rect 3608 13738 3660 13744
rect 3620 13190 3648 13738
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3514 12744 3570 12753
rect 3514 12679 3570 12688
rect 3620 12238 3648 13126
rect 3804 12850 3832 13466
rect 3896 13462 3924 14282
rect 3988 13462 4016 19450
rect 4172 18290 4200 19638
rect 4250 18592 4306 18601
rect 4250 18527 4306 18536
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4066 18048 4122 18057
rect 4066 17983 4122 17992
rect 4080 17746 4108 17983
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 4172 17202 4200 18226
rect 4264 17882 4292 18527
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4356 17762 4384 20726
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 4436 19984 4488 19990
rect 4436 19926 4488 19932
rect 4448 19514 4476 19926
rect 4540 19922 4568 20402
rect 4632 20058 4660 20878
rect 4620 20052 4672 20058
rect 4620 19994 4672 20000
rect 4528 19916 4580 19922
rect 4528 19858 4580 19864
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4540 19378 4568 19858
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 4356 17734 4568 17762
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4448 17270 4476 17614
rect 4436 17264 4488 17270
rect 4436 17206 4488 17212
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4068 16992 4120 16998
rect 4356 16969 4384 17138
rect 4068 16934 4120 16940
rect 4342 16960 4398 16969
rect 4080 16674 4108 16934
rect 4342 16895 4398 16904
rect 4080 16646 4292 16674
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 4066 16144 4122 16153
rect 4066 16079 4122 16088
rect 3884 13456 3936 13462
rect 3884 13398 3936 13404
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 3882 13288 3938 13297
rect 4080 13258 4108 16079
rect 4172 15910 4200 16526
rect 4160 15904 4212 15910
rect 4158 15872 4160 15881
rect 4212 15872 4214 15881
rect 4158 15807 4214 15816
rect 4264 15609 4292 16646
rect 4356 16250 4384 16895
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4356 15706 4384 16186
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4250 15600 4306 15609
rect 4160 15564 4212 15570
rect 4306 15558 4384 15586
rect 4250 15535 4306 15544
rect 4160 15506 4212 15512
rect 4172 14822 4200 15506
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4172 13326 4200 14758
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 3882 13223 3938 13232
rect 4068 13252 4120 13258
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3804 12730 3832 12786
rect 3712 12702 3832 12730
rect 3608 12232 3660 12238
rect 3422 12200 3478 12209
rect 3608 12174 3660 12180
rect 3422 12135 3478 12144
rect 3620 11762 3648 12174
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 3528 2145 3556 11630
rect 3620 11354 3648 11698
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3712 4978 3740 12702
rect 3896 11234 3924 13223
rect 4068 13194 4120 13200
rect 4264 12850 4292 13398
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4080 12442 4108 12718
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4264 12186 4292 12786
rect 4356 12442 4384 15558
rect 4448 14657 4476 17206
rect 4540 15065 4568 17734
rect 4618 16280 4674 16289
rect 4618 16215 4674 16224
rect 4526 15056 4582 15065
rect 4526 14991 4582 15000
rect 4434 14648 4490 14657
rect 4434 14583 4490 14592
rect 4448 13734 4476 14583
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 3988 12158 4292 12186
rect 3988 11558 4016 12158
rect 4066 11928 4122 11937
rect 4356 11898 4384 12378
rect 4632 12306 4660 16215
rect 4724 15745 4752 24398
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4816 22522 4844 24142
rect 4896 24064 4948 24070
rect 4896 24006 4948 24012
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 4908 23662 4936 24006
rect 5080 23860 5132 23866
rect 5080 23802 5132 23808
rect 4896 23656 4948 23662
rect 4896 23598 4948 23604
rect 4908 22778 4936 23598
rect 4988 23112 5040 23118
rect 4988 23054 5040 23060
rect 5092 23066 5120 23802
rect 5276 23730 5304 24006
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5170 23624 5226 23633
rect 5170 23559 5226 23568
rect 5184 23526 5212 23559
rect 5172 23520 5224 23526
rect 5460 23508 5488 24550
rect 6090 24511 6146 24520
rect 6288 24274 6316 25094
rect 6380 24800 6408 27520
rect 6380 24772 6500 24800
rect 6368 24676 6420 24682
rect 6368 24618 6420 24624
rect 5540 24268 5592 24274
rect 5540 24210 5592 24216
rect 6276 24268 6328 24274
rect 6276 24210 6328 24216
rect 5172 23462 5224 23468
rect 5368 23480 5488 23508
rect 4896 22772 4948 22778
rect 4896 22714 4948 22720
rect 5000 22710 5028 23054
rect 5092 23038 5212 23066
rect 5080 22976 5132 22982
rect 5080 22918 5132 22924
rect 4988 22704 5040 22710
rect 4988 22646 5040 22652
rect 5092 22642 5120 22918
rect 5080 22636 5132 22642
rect 5080 22578 5132 22584
rect 4816 22494 5120 22522
rect 4894 22400 4950 22409
rect 4894 22335 4950 22344
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 4816 18902 4844 19178
rect 4804 18896 4856 18902
rect 4804 18838 4856 18844
rect 4816 17882 4844 18838
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4804 16516 4856 16522
rect 4804 16458 4856 16464
rect 4816 16046 4844 16458
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4710 15736 4766 15745
rect 4710 15671 4766 15680
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4724 14074 4752 14418
rect 4816 14414 4844 15302
rect 4908 14550 4936 22335
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 5000 16454 5028 17002
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 5000 15366 5028 16390
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 4896 14544 4948 14550
rect 4896 14486 4948 14492
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4816 13308 4844 14350
rect 4908 14074 4936 14486
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4908 13530 4936 14010
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4896 13320 4948 13326
rect 4816 13280 4896 13308
rect 4896 13262 4948 13268
rect 4710 12880 4766 12889
rect 4908 12850 4936 13262
rect 4710 12815 4712 12824
rect 4764 12815 4766 12824
rect 4896 12844 4948 12850
rect 4712 12786 4764 12792
rect 4896 12786 4948 12792
rect 4710 12336 4766 12345
rect 4620 12300 4672 12306
rect 4710 12271 4766 12280
rect 4620 12242 4672 12248
rect 4066 11863 4122 11872
rect 4344 11892 4396 11898
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 4080 11257 4108 11863
rect 4344 11834 4396 11840
rect 4632 11830 4660 12242
rect 4724 12238 4752 12271
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4724 11898 4752 12174
rect 4908 12170 4936 12786
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4632 11529 4660 11766
rect 4618 11520 4674 11529
rect 4618 11455 4674 11464
rect 4066 11248 4122 11257
rect 3896 11206 4016 11234
rect 3882 11112 3938 11121
rect 3882 11047 3938 11056
rect 3896 5137 3924 11047
rect 3882 5128 3938 5137
rect 3882 5063 3938 5072
rect 3712 4950 3924 4978
rect 3514 2136 3570 2145
rect 3514 2071 3570 2080
rect 3896 1465 3924 4950
rect 3988 4434 4016 11206
rect 4066 11183 4122 11192
rect 4066 9616 4122 9625
rect 4066 9551 4122 9560
rect 4080 8809 4108 9551
rect 4066 8800 4122 8809
rect 4066 8735 4122 8744
rect 4066 7848 4122 7857
rect 4066 7783 4122 7792
rect 4080 7041 4108 7783
rect 4066 7032 4122 7041
rect 4066 6967 4122 6976
rect 4066 5264 4122 5273
rect 4066 5199 4122 5208
rect 4080 4593 4108 5199
rect 5092 5137 5120 22494
rect 5184 22250 5212 23038
rect 5368 22438 5396 23480
rect 5448 23316 5500 23322
rect 5552 23304 5580 24210
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5500 23276 5580 23304
rect 5448 23258 5500 23264
rect 6184 23180 6236 23186
rect 6184 23122 6236 23128
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5816 22636 5868 22642
rect 5816 22578 5868 22584
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 5446 22264 5502 22273
rect 5184 22222 5396 22250
rect 5262 21720 5318 21729
rect 5262 21655 5318 21664
rect 5276 21486 5304 21655
rect 5264 21480 5316 21486
rect 5264 21422 5316 21428
rect 5276 21010 5304 21422
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5184 16794 5212 18702
rect 5276 17882 5304 18770
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5368 16794 5396 22222
rect 5828 22234 5856 22578
rect 6196 22574 6224 23122
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 5446 22199 5502 22208
rect 5816 22228 5868 22234
rect 5460 21554 5488 22199
rect 5816 22170 5868 22176
rect 6196 22166 6224 22510
rect 6184 22160 6236 22166
rect 6184 22102 6236 22108
rect 6090 21992 6146 22001
rect 6090 21927 6092 21936
rect 6144 21927 6146 21936
rect 6092 21898 6144 21904
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6196 21690 6224 22102
rect 6288 21894 6316 24210
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 5448 21548 5500 21554
rect 5448 21490 5500 21496
rect 5460 21146 5488 21490
rect 6288 21146 6316 21830
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 6380 21026 6408 24618
rect 6472 23905 6500 24772
rect 6932 24698 6960 27520
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 7208 24818 7236 25094
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 6932 24670 7144 24698
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 6932 24449 6960 24550
rect 6918 24440 6974 24449
rect 6918 24375 6974 24384
rect 6552 24336 6604 24342
rect 6552 24278 6604 24284
rect 6458 23896 6514 23905
rect 6458 23831 6514 23840
rect 6564 23662 6592 24278
rect 6920 24132 6972 24138
rect 6920 24074 6972 24080
rect 6552 23656 6604 23662
rect 6552 23598 6604 23604
rect 6564 23526 6592 23598
rect 6932 23526 6960 24074
rect 7012 24064 7064 24070
rect 7012 24006 7064 24012
rect 7024 23730 7052 24006
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 6552 23520 6604 23526
rect 6920 23520 6972 23526
rect 6552 23462 6604 23468
rect 6840 23480 6920 23508
rect 6564 22982 6592 23462
rect 6552 22976 6604 22982
rect 6552 22918 6604 22924
rect 6564 22642 6592 22918
rect 6552 22636 6604 22642
rect 6552 22578 6604 22584
rect 6736 22024 6788 22030
rect 6656 21984 6736 22012
rect 6656 21350 6684 21984
rect 6736 21966 6788 21972
rect 6840 21962 6868 23480
rect 7116 23474 7144 24670
rect 7208 24410 7236 24754
rect 7196 24404 7248 24410
rect 7196 24346 7248 24352
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 6920 23462 6972 23468
rect 7024 23446 7144 23474
rect 7024 22778 7052 23446
rect 7102 23352 7158 23361
rect 7300 23322 7328 23666
rect 7102 23287 7158 23296
rect 7288 23316 7340 23322
rect 7012 22772 7064 22778
rect 7012 22714 7064 22720
rect 7116 22234 7144 23287
rect 7288 23258 7340 23264
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7196 22976 7248 22982
rect 7196 22918 7248 22924
rect 7208 22438 7236 22918
rect 7286 22536 7342 22545
rect 7286 22471 7288 22480
rect 7340 22471 7342 22480
rect 7288 22442 7340 22448
rect 7196 22432 7248 22438
rect 7194 22400 7196 22409
rect 7248 22400 7250 22409
rect 7194 22335 7250 22344
rect 7104 22228 7156 22234
rect 7104 22170 7156 22176
rect 6828 21956 6880 21962
rect 6828 21898 6880 21904
rect 7116 21350 7144 22170
rect 7392 21894 7420 23054
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7484 22030 7512 22578
rect 7472 22024 7524 22030
rect 7472 21966 7524 21972
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 7392 21486 7420 21830
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 6092 21004 6144 21010
rect 6092 20946 6144 20952
rect 6196 20998 6408 21026
rect 6552 21004 6604 21010
rect 6104 20806 6132 20946
rect 6092 20800 6144 20806
rect 6092 20742 6144 20748
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5998 20632 6054 20641
rect 5998 20567 6000 20576
rect 6052 20567 6054 20576
rect 6000 20538 6052 20544
rect 5540 20324 5592 20330
rect 5540 20266 5592 20272
rect 5552 19174 5580 20266
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5998 19272 6054 19281
rect 5998 19207 6054 19216
rect 6012 19174 6040 19207
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6104 18850 6132 20742
rect 6012 18822 6132 18850
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5908 18352 5960 18358
rect 5908 18294 5960 18300
rect 5920 17678 5948 18294
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 5920 17524 5948 17614
rect 6012 17592 6040 18822
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 6104 18222 6132 18702
rect 6092 18216 6144 18222
rect 6090 18184 6092 18193
rect 6144 18184 6146 18193
rect 6090 18119 6146 18128
rect 6012 17564 6132 17592
rect 5920 17496 6040 17524
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 5184 16046 5212 16390
rect 5368 16250 5396 16730
rect 6012 16590 6040 17496
rect 6104 17202 6132 17564
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 6090 17096 6146 17105
rect 6090 17031 6146 17040
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 16250 6040 16526
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5170 15192 5226 15201
rect 5170 15127 5172 15136
rect 5224 15127 5226 15136
rect 5172 15098 5224 15104
rect 5276 14793 5304 15846
rect 5262 14784 5318 14793
rect 5262 14719 5318 14728
rect 5354 14648 5410 14657
rect 5354 14583 5410 14592
rect 5368 14550 5396 14583
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5170 14376 5226 14385
rect 5170 14311 5226 14320
rect 5184 14074 5212 14311
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5368 13870 5396 14486
rect 5460 14482 5488 16118
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 5538 15464 5594 15473
rect 5538 15399 5540 15408
rect 5592 15399 5594 15408
rect 5540 15370 5592 15376
rect 5552 14958 5580 15370
rect 6012 15366 6040 16050
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5632 14816 5684 14822
rect 5630 14784 5632 14793
rect 5684 14784 5686 14793
rect 5630 14719 5686 14728
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 6012 14278 6040 15302
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5184 13530 5212 13670
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5170 12880 5226 12889
rect 5170 12815 5226 12824
rect 5184 12442 5212 12815
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5552 12238 5580 13874
rect 5644 13530 5672 13874
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 6012 13394 6040 14214
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6012 12986 6040 13330
rect 6104 12986 6132 17031
rect 6196 16794 6224 20998
rect 6552 20946 6604 20952
rect 6564 20602 6592 20946
rect 6656 20777 6684 21286
rect 7116 21049 7144 21286
rect 7102 21040 7158 21049
rect 7102 20975 7158 20984
rect 6920 20936 6972 20942
rect 6972 20884 7052 20890
rect 6920 20878 7052 20884
rect 6736 20868 6788 20874
rect 6932 20862 7052 20878
rect 6736 20810 6788 20816
rect 6642 20768 6698 20777
rect 6642 20703 6698 20712
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6642 20224 6698 20233
rect 6642 20159 6698 20168
rect 6276 19848 6328 19854
rect 6276 19790 6328 19796
rect 6288 18902 6316 19790
rect 6276 18896 6328 18902
rect 6276 18838 6328 18844
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6288 16998 6316 17682
rect 6380 17542 6408 18770
rect 6552 18692 6604 18698
rect 6552 18634 6604 18640
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6196 16182 6224 16594
rect 6288 16561 6316 16934
rect 6274 16552 6330 16561
rect 6274 16487 6330 16496
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6184 16176 6236 16182
rect 6184 16118 6236 16124
rect 6288 15910 6316 16390
rect 6380 16153 6408 17478
rect 6472 16833 6500 18566
rect 6564 18426 6592 18634
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6564 17338 6592 18362
rect 6656 17377 6684 20159
rect 6748 20058 6776 20810
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6932 20058 6960 20742
rect 7024 20602 7052 20862
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 7392 20398 7420 21422
rect 7576 20942 7604 27520
rect 8128 24834 8156 27520
rect 7852 24806 8156 24834
rect 8392 24812 8444 24818
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 7656 24064 7708 24070
rect 7656 24006 7708 24012
rect 7668 23186 7696 24006
rect 7760 23361 7788 24550
rect 7746 23352 7802 23361
rect 7746 23287 7802 23296
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 7668 22234 7696 23122
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 7668 21146 7696 21422
rect 7746 21176 7802 21185
rect 7656 21140 7708 21146
rect 7746 21111 7802 21120
rect 7656 21082 7708 21088
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7576 20602 7604 20878
rect 7564 20596 7616 20602
rect 7564 20538 7616 20544
rect 7562 20496 7618 20505
rect 7562 20431 7618 20440
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6748 19378 6776 19994
rect 7194 19952 7250 19961
rect 7194 19887 7250 19896
rect 7288 19916 7340 19922
rect 6918 19816 6974 19825
rect 6918 19751 6920 19760
rect 6972 19751 6974 19760
rect 6920 19722 6972 19728
rect 7208 19718 7236 19887
rect 7288 19858 7340 19864
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7300 19514 7328 19858
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6748 18358 6776 19314
rect 6840 18970 6868 19450
rect 7576 19417 7604 20431
rect 7562 19408 7618 19417
rect 7472 19372 7524 19378
rect 7562 19343 7618 19352
rect 7472 19314 7524 19320
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6736 18352 6788 18358
rect 6736 18294 6788 18300
rect 6826 18320 6882 18329
rect 6642 17368 6698 17377
rect 6552 17332 6604 17338
rect 6748 17338 6776 18294
rect 6826 18255 6882 18264
rect 6840 18222 6868 18255
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6840 18034 6868 18158
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 7116 18057 7144 18090
rect 7102 18048 7158 18057
rect 6840 18006 6960 18034
rect 6932 17746 6960 18006
rect 7102 17983 7158 17992
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 7208 17542 7236 19110
rect 7300 18737 7328 19110
rect 7484 18970 7512 19314
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7286 18728 7342 18737
rect 7286 18663 7342 18672
rect 7656 18692 7708 18698
rect 7656 18634 7708 18640
rect 7668 18086 7696 18634
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7668 17746 7696 18022
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7668 17338 7696 17682
rect 6642 17303 6698 17312
rect 6736 17332 6788 17338
rect 6552 17274 6604 17280
rect 6736 17274 6788 17280
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 6918 17232 6974 17241
rect 6552 17196 6604 17202
rect 7760 17202 7788 21111
rect 7852 20210 7880 24806
rect 8392 24754 8444 24760
rect 7932 24744 7984 24750
rect 7932 24686 7984 24692
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 7944 20346 7972 24686
rect 8312 24313 8340 24686
rect 8298 24304 8354 24313
rect 8298 24239 8354 24248
rect 8116 24064 8168 24070
rect 8116 24006 8168 24012
rect 8128 22001 8156 24006
rect 8298 23896 8354 23905
rect 8298 23831 8300 23840
rect 8352 23831 8354 23840
rect 8300 23802 8352 23808
rect 8300 23724 8352 23730
rect 8300 23666 8352 23672
rect 8208 22636 8260 22642
rect 8312 22624 8340 23666
rect 8404 22982 8432 24754
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8496 24410 8524 24550
rect 8484 24404 8536 24410
rect 8484 24346 8536 24352
rect 8574 23216 8630 23225
rect 8574 23151 8630 23160
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 8260 22596 8340 22624
rect 8208 22578 8260 22584
rect 8404 22522 8432 22918
rect 8220 22494 8432 22522
rect 8114 21992 8170 22001
rect 8114 21927 8170 21936
rect 8022 21312 8078 21321
rect 8022 21247 8078 21256
rect 8036 21146 8064 21247
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 8128 21078 8156 21927
rect 8220 21486 8248 22494
rect 8392 22432 8444 22438
rect 8392 22374 8444 22380
rect 8404 22273 8432 22374
rect 8390 22264 8446 22273
rect 8390 22199 8446 22208
rect 8208 21480 8260 21486
rect 8208 21422 8260 21428
rect 8390 21448 8446 21457
rect 8390 21383 8446 21392
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 8116 21072 8168 21078
rect 8116 21014 8168 21020
rect 7944 20318 8064 20346
rect 8128 20330 8156 21014
rect 8312 21010 8340 21082
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8036 20262 8064 20318
rect 8116 20324 8168 20330
rect 8116 20266 8168 20272
rect 8024 20256 8076 20262
rect 7852 20182 7972 20210
rect 8024 20198 8076 20204
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7852 18970 7880 19994
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 7944 18465 7972 20182
rect 8208 20052 8260 20058
rect 8312 20040 8340 20946
rect 8404 20913 8432 21383
rect 8588 21146 8616 23151
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8680 21026 8708 27520
rect 9232 27470 9260 27520
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 8760 25696 8812 25702
rect 8760 25638 8812 25644
rect 8772 25498 8800 25638
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 9312 25152 9364 25158
rect 9312 25094 9364 25100
rect 9324 24954 9352 25094
rect 9312 24948 9364 24954
rect 9312 24890 9364 24896
rect 9128 24744 9180 24750
rect 9128 24686 9180 24692
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8956 24177 8984 24550
rect 9036 24336 9088 24342
rect 9036 24278 9088 24284
rect 8942 24168 8998 24177
rect 8942 24103 8998 24112
rect 8944 24064 8996 24070
rect 8944 24006 8996 24012
rect 8852 23860 8904 23866
rect 8852 23802 8904 23808
rect 8864 23769 8892 23802
rect 8850 23760 8906 23769
rect 8956 23730 8984 24006
rect 8850 23695 8906 23704
rect 8944 23724 8996 23730
rect 8864 23594 8892 23695
rect 8944 23666 8996 23672
rect 8852 23588 8904 23594
rect 8852 23530 8904 23536
rect 9048 23322 9076 24278
rect 9036 23316 9088 23322
rect 9036 23258 9088 23264
rect 9140 22953 9168 24686
rect 9126 22944 9182 22953
rect 9126 22879 9182 22888
rect 8944 22772 8996 22778
rect 8944 22714 8996 22720
rect 8758 21992 8814 22001
rect 8758 21927 8814 21936
rect 8772 21690 8800 21927
rect 8760 21684 8812 21690
rect 8760 21626 8812 21632
rect 8496 20998 8708 21026
rect 8390 20904 8446 20913
rect 8390 20839 8446 20848
rect 8260 20012 8340 20040
rect 8208 19994 8260 20000
rect 8496 18952 8524 20998
rect 8668 20936 8720 20942
rect 8668 20878 8720 20884
rect 8680 20058 8708 20878
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 8588 19417 8616 19790
rect 8574 19408 8630 19417
rect 8574 19343 8630 19352
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8680 19174 8708 19246
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8312 18924 8524 18952
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 7930 18456 7986 18465
rect 7852 18414 7930 18442
rect 6918 17167 6974 17176
rect 7748 17196 7800 17202
rect 6552 17138 6604 17144
rect 6458 16824 6514 16833
rect 6458 16759 6514 16768
rect 6460 16720 6512 16726
rect 6460 16662 6512 16668
rect 6366 16144 6422 16153
rect 6366 16079 6422 16088
rect 6472 15994 6500 16662
rect 6564 16658 6592 17138
rect 6932 16794 6960 17167
rect 7748 17138 7800 17144
rect 7654 16960 7710 16969
rect 7654 16895 7710 16904
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 7668 16726 7696 16895
rect 7656 16720 7708 16726
rect 6734 16688 6790 16697
rect 6552 16652 6604 16658
rect 7656 16662 7708 16668
rect 6734 16623 6736 16632
rect 6552 16594 6604 16600
rect 6788 16623 6790 16632
rect 6736 16594 6788 16600
rect 6380 15966 6500 15994
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6182 15328 6238 15337
rect 6182 15263 6238 15272
rect 6196 13297 6224 15263
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6288 15065 6316 15098
rect 6274 15056 6330 15065
rect 6274 14991 6330 15000
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6288 14550 6316 14894
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 6288 14074 6316 14486
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6380 13433 6408 15966
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6472 14385 6500 15506
rect 6564 15337 6592 16594
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 6918 16144 6974 16153
rect 6918 16079 6974 16088
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6550 15328 6606 15337
rect 6550 15263 6606 15272
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6458 14376 6514 14385
rect 6458 14311 6514 14320
rect 6564 14074 6592 14962
rect 6656 14657 6684 15846
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6642 14648 6698 14657
rect 6748 14618 6776 15438
rect 6642 14583 6698 14592
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6840 13870 6868 14418
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 13462 6868 13806
rect 6828 13456 6880 13462
rect 6366 13424 6422 13433
rect 6828 13398 6880 13404
rect 6366 13359 6422 13368
rect 6182 13288 6238 13297
rect 6840 13258 6868 13398
rect 6182 13223 6238 13232
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6840 12442 6868 13194
rect 6932 12481 6960 16079
rect 7024 15162 7052 16390
rect 7116 16046 7144 16390
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7562 15872 7618 15881
rect 7562 15807 7618 15816
rect 7576 15366 7604 15807
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7378 15056 7434 15065
rect 7378 14991 7434 15000
rect 7392 14890 7420 14991
rect 7380 14884 7432 14890
rect 7380 14826 7432 14832
rect 7576 14822 7604 15302
rect 7668 15026 7696 15574
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7472 14408 7524 14414
rect 7470 14376 7472 14385
rect 7524 14376 7526 14385
rect 7470 14311 7526 14320
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7116 13530 7144 13806
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7194 13016 7250 13025
rect 7194 12951 7250 12960
rect 7208 12714 7236 12951
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7196 12708 7248 12714
rect 7196 12650 7248 12656
rect 6918 12472 6974 12481
rect 6828 12436 6880 12442
rect 7300 12442 7328 12718
rect 6918 12407 6974 12416
rect 7288 12436 7340 12442
rect 6828 12378 6880 12384
rect 7288 12378 7340 12384
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 7576 11801 7604 14758
rect 7852 13376 7880 18414
rect 7930 18391 7986 18400
rect 8036 18193 8064 18566
rect 8116 18216 8168 18222
rect 8022 18184 8078 18193
rect 8116 18158 8168 18164
rect 8022 18119 8078 18128
rect 8128 17814 8156 18158
rect 8116 17808 8168 17814
rect 8116 17750 8168 17756
rect 8128 17252 8156 17750
rect 8036 17224 8156 17252
rect 8036 17134 8064 17224
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8206 16688 8262 16697
rect 8128 16646 8206 16674
rect 8128 16250 8156 16646
rect 8206 16623 8208 16632
rect 8260 16623 8262 16632
rect 8208 16594 8260 16600
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8220 16425 8248 16458
rect 8206 16416 8262 16425
rect 8206 16351 8262 16360
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7944 15366 7972 15982
rect 8220 15706 8248 16351
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 8022 15192 8078 15201
rect 8022 15127 8078 15136
rect 8036 14618 8064 15127
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8024 13456 8076 13462
rect 8024 13398 8076 13404
rect 7760 13348 7880 13376
rect 7760 12782 7788 13348
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7852 12646 7880 13194
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7944 12889 7972 13126
rect 8036 12986 8064 13398
rect 8312 13326 8340 18924
rect 8588 18873 8616 19110
rect 8574 18864 8630 18873
rect 8392 18828 8444 18834
rect 8574 18799 8630 18808
rect 8392 18770 8444 18776
rect 8404 16794 8432 18770
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8496 18426 8524 18702
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8496 17882 8524 18362
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8574 16552 8630 16561
rect 8574 16487 8630 16496
rect 8390 15736 8446 15745
rect 8390 15671 8446 15680
rect 8484 15700 8536 15706
rect 8404 15570 8432 15671
rect 8484 15642 8536 15648
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8404 15094 8432 15506
rect 8496 15162 8524 15642
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8392 15088 8444 15094
rect 8392 15030 8444 15036
rect 8404 14482 8432 15030
rect 8496 14618 8524 15098
rect 8588 15026 8616 16487
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8404 13938 8432 14418
rect 8496 14074 8524 14554
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8496 13326 8524 13670
rect 8300 13320 8352 13326
rect 8220 13280 8300 13308
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7930 12880 7986 12889
rect 7930 12815 7986 12824
rect 8220 12866 8248 13280
rect 8300 13262 8352 13268
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8574 13288 8630 13297
rect 8300 12912 8352 12918
rect 8220 12860 8300 12866
rect 8220 12854 8352 12860
rect 8220 12838 8340 12854
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 8220 12442 8248 12838
rect 8496 12442 8524 13262
rect 8574 13223 8630 13232
rect 8588 12782 8616 13223
rect 8680 12850 8708 19110
rect 8758 17776 8814 17785
rect 8758 17711 8814 17720
rect 8772 17610 8800 17711
rect 8760 17604 8812 17610
rect 8760 17546 8812 17552
rect 8772 17134 8800 17546
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8760 16720 8812 16726
rect 8760 16662 8812 16668
rect 8772 14618 8800 16662
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8588 12442 8616 12718
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8496 12345 8524 12378
rect 8482 12336 8538 12345
rect 8482 12271 8538 12280
rect 7562 11792 7618 11801
rect 7562 11727 7618 11736
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 8298 5672 8354 5681
rect 8298 5607 8354 5616
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5078 5128 5134 5137
rect 5078 5063 5134 5072
rect 4066 4584 4122 4593
rect 4066 4519 4122 4528
rect 3988 4406 4108 4434
rect 3882 1456 3938 1465
rect 3882 1391 3938 1400
rect 3238 912 3294 921
rect 3238 847 3294 856
rect 2778 0 2834 480
rect 4080 377 4108 4406
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 8312 3913 8340 5607
rect 8298 3904 8354 3913
rect 8298 3839 8354 3848
rect 8864 3641 8892 20198
rect 8956 19802 8984 22714
rect 9036 22636 9088 22642
rect 9036 22578 9088 22584
rect 9048 21962 9076 22578
rect 9128 22092 9180 22098
rect 9128 22034 9180 22040
rect 9036 21956 9088 21962
rect 9036 21898 9088 21904
rect 9048 20641 9076 21898
rect 9140 21729 9168 22034
rect 9126 21720 9182 21729
rect 9126 21655 9128 21664
rect 9180 21655 9182 21664
rect 9128 21626 9180 21632
rect 9416 21554 9444 27406
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 9508 24206 9536 24754
rect 9784 24410 9812 27520
rect 10336 25786 10364 27520
rect 10152 25758 10364 25786
rect 10692 25832 10744 25838
rect 10692 25774 10744 25780
rect 9956 25356 10008 25362
rect 9956 25298 10008 25304
rect 9968 24614 9996 25298
rect 9956 24608 10008 24614
rect 9862 24576 9918 24585
rect 9956 24550 10008 24556
rect 9862 24511 9918 24520
rect 9772 24404 9824 24410
rect 9772 24346 9824 24352
rect 9496 24200 9548 24206
rect 9496 24142 9548 24148
rect 9784 23866 9812 24346
rect 9876 24342 9904 24511
rect 9864 24336 9916 24342
rect 9968 24313 9996 24550
rect 9864 24278 9916 24284
rect 9954 24304 10010 24313
rect 9876 24018 9904 24278
rect 9954 24239 10010 24248
rect 9876 23990 9996 24018
rect 9772 23860 9824 23866
rect 9824 23820 9904 23848
rect 9772 23802 9824 23808
rect 9772 23520 9824 23526
rect 9692 23480 9772 23508
rect 9588 23316 9640 23322
rect 9692 23304 9720 23480
rect 9772 23462 9824 23468
rect 9640 23276 9720 23304
rect 9770 23352 9826 23361
rect 9770 23287 9772 23296
rect 9588 23258 9640 23264
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9508 22778 9536 23054
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 9588 22092 9640 22098
rect 9588 22034 9640 22040
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9034 20632 9090 20641
rect 9034 20567 9090 20576
rect 8956 19774 9076 19802
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 8956 18222 8984 19654
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8956 16250 8984 16526
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 8956 15638 8984 16186
rect 9048 15910 9076 19774
rect 9140 19514 9168 21490
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9416 20398 9444 20742
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9416 20262 9444 20334
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9416 19718 9444 20198
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 9140 18698 9168 19314
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9128 18692 9180 18698
rect 9128 18634 9180 18640
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 8944 15632 8996 15638
rect 9140 15609 9168 17478
rect 8944 15574 8996 15580
rect 9126 15600 9182 15609
rect 9126 15535 9182 15544
rect 9126 13832 9182 13841
rect 9126 13767 9128 13776
rect 9180 13767 9182 13776
rect 9128 13738 9180 13744
rect 9140 13530 9168 13738
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9232 11937 9260 19110
rect 9324 15706 9352 19382
rect 9404 18896 9456 18902
rect 9404 18838 9456 18844
rect 9416 17882 9444 18838
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9416 15978 9444 16934
rect 9404 15972 9456 15978
rect 9404 15914 9456 15920
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9416 15502 9444 15914
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9416 15162 9444 15438
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9218 11928 9274 11937
rect 9218 11863 9274 11872
rect 9232 10033 9260 11863
rect 9508 10713 9536 21966
rect 9600 20788 9628 22034
rect 9692 21690 9720 23276
rect 9824 23287 9826 23296
rect 9772 23258 9824 23264
rect 9772 23044 9824 23050
rect 9772 22986 9824 22992
rect 9784 22710 9812 22986
rect 9772 22704 9824 22710
rect 9772 22646 9824 22652
rect 9784 22001 9812 22646
rect 9770 21992 9826 22001
rect 9770 21927 9826 21936
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9680 21344 9732 21350
rect 9678 21312 9680 21321
rect 9732 21312 9734 21321
rect 9678 21247 9734 21256
rect 9784 21185 9812 21830
rect 9770 21176 9826 21185
rect 9770 21111 9826 21120
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 9680 20800 9732 20806
rect 9600 20760 9680 20788
rect 9680 20742 9732 20748
rect 9692 20346 9720 20742
rect 9784 20466 9812 20946
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9692 20318 9812 20346
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9692 18970 9720 19314
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9588 18692 9640 18698
rect 9588 18634 9640 18640
rect 9600 18358 9628 18634
rect 9784 18601 9812 20318
rect 9876 19922 9904 23820
rect 9968 23730 9996 23990
rect 10152 23905 10180 25758
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10704 25498 10732 25774
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10888 24800 10916 27520
rect 10968 26036 11020 26042
rect 10968 25978 11020 25984
rect 10704 24772 10916 24800
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10704 24154 10732 24772
rect 10980 24698 11008 25978
rect 11244 25424 11296 25430
rect 11244 25366 11296 25372
rect 11256 24818 11284 25366
rect 11336 25152 11388 25158
rect 11336 25094 11388 25100
rect 11244 24812 11296 24818
rect 11244 24754 11296 24760
rect 10876 24676 10928 24682
rect 10980 24670 11192 24698
rect 10876 24618 10928 24624
rect 10784 24608 10836 24614
rect 10784 24550 10836 24556
rect 10612 24126 10732 24154
rect 10138 23896 10194 23905
rect 10138 23831 10194 23840
rect 10152 23746 10180 23831
rect 9956 23724 10008 23730
rect 9956 23666 10008 23672
rect 10060 23718 10180 23746
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9876 19242 9904 19858
rect 9968 19310 9996 23666
rect 10060 23662 10088 23718
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 10060 21894 10088 23122
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 10060 21350 10088 21490
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 10060 20806 10088 21286
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 10060 20330 10088 20742
rect 10048 20324 10100 20330
rect 10048 20266 10100 20272
rect 10060 19854 10088 20266
rect 10152 20058 10180 23598
rect 10612 23594 10640 24126
rect 10692 24064 10744 24070
rect 10692 24006 10744 24012
rect 10704 23730 10732 24006
rect 10692 23724 10744 23730
rect 10692 23666 10744 23672
rect 10600 23588 10652 23594
rect 10600 23530 10652 23536
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 10612 22574 10640 23054
rect 10600 22568 10652 22574
rect 10600 22510 10652 22516
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10336 20330 10364 20946
rect 10704 20584 10732 23666
rect 10796 23662 10824 24550
rect 10888 24449 10916 24618
rect 10968 24608 11020 24614
rect 10966 24576 10968 24585
rect 11020 24576 11022 24585
rect 10966 24511 11022 24520
rect 10874 24440 10930 24449
rect 10874 24375 10930 24384
rect 11060 24132 11112 24138
rect 11060 24074 11112 24080
rect 11072 24018 11100 24074
rect 10980 23990 11100 24018
rect 10876 23792 10928 23798
rect 10876 23734 10928 23740
rect 10784 23656 10836 23662
rect 10784 23598 10836 23604
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10796 23118 10824 23462
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10796 22506 10824 22918
rect 10784 22500 10836 22506
rect 10784 22442 10836 22448
rect 10784 22228 10836 22234
rect 10784 22170 10836 22176
rect 10796 21876 10824 22170
rect 10888 21978 10916 23734
rect 10980 22778 11008 23990
rect 10968 22772 11020 22778
rect 10968 22714 11020 22720
rect 11164 22658 11192 24670
rect 11348 24410 11376 25094
rect 11336 24404 11388 24410
rect 11336 24346 11388 24352
rect 11348 23662 11376 24346
rect 11440 24290 11468 27520
rect 11612 26240 11664 26246
rect 11612 26182 11664 26188
rect 11624 25498 11652 26182
rect 11612 25492 11664 25498
rect 11612 25434 11664 25440
rect 11992 24698 12020 27520
rect 12164 25288 12216 25294
rect 12164 25230 12216 25236
rect 11808 24670 12020 24698
rect 11440 24262 11560 24290
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 11440 23866 11468 24142
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 11336 23656 11388 23662
rect 11336 23598 11388 23604
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 10980 22630 11192 22658
rect 10980 22098 11008 22630
rect 10968 22092 11020 22098
rect 10968 22034 11020 22040
rect 10888 21950 11100 21978
rect 10968 21888 11020 21894
rect 10796 21848 10916 21876
rect 10784 20596 10836 20602
rect 10704 20556 10784 20584
rect 10324 20324 10376 20330
rect 10324 20266 10376 20272
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 10060 19514 10088 19790
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 10138 19272 10194 19281
rect 9864 19236 9916 19242
rect 10138 19207 10194 19216
rect 9864 19178 9916 19184
rect 10152 19174 10180 19207
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10704 18902 10732 20556
rect 10784 20538 10836 20544
rect 10782 20088 10838 20097
rect 10782 20023 10784 20032
rect 10836 20023 10838 20032
rect 10784 19994 10836 20000
rect 10692 18896 10744 18902
rect 10692 18838 10744 18844
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 9770 18592 9826 18601
rect 9770 18527 9826 18536
rect 9954 18456 10010 18465
rect 9954 18391 10010 18400
rect 9968 18358 9996 18391
rect 9588 18352 9640 18358
rect 9588 18294 9640 18300
rect 9956 18352 10008 18358
rect 9956 18294 10008 18300
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9876 17338 9904 17682
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9678 16416 9734 16425
rect 9678 16351 9734 16360
rect 9692 16250 9720 16351
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9876 15502 9904 16594
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9680 15360 9732 15366
rect 9784 15337 9812 15438
rect 9680 15302 9732 15308
rect 9770 15328 9826 15337
rect 9692 15178 9720 15302
rect 9770 15263 9826 15272
rect 9692 15150 9812 15178
rect 9784 14958 9812 15150
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9784 14618 9812 14894
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 12866 9720 14214
rect 9784 13870 9812 14554
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9784 13530 9812 13806
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9784 13258 9812 13466
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9968 13025 9996 18022
rect 10060 17882 10088 18090
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10704 17678 10732 18702
rect 10888 18154 10916 21848
rect 10968 21830 11020 21836
rect 10980 21350 11008 21830
rect 11072 21486 11100 21950
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 10968 21344 11020 21350
rect 11020 21292 11100 21298
rect 10968 21286 11100 21292
rect 10980 21270 11100 21286
rect 11072 20058 11100 21270
rect 11256 21146 11284 23258
rect 11348 23118 11376 23598
rect 11532 23225 11560 24262
rect 11518 23216 11574 23225
rect 11518 23151 11574 23160
rect 11612 23180 11664 23186
rect 11612 23122 11664 23128
rect 11336 23112 11388 23118
rect 11388 23072 11560 23100
rect 11336 23054 11388 23060
rect 11336 22568 11388 22574
rect 11336 22510 11388 22516
rect 11348 22166 11376 22510
rect 11532 22386 11560 23072
rect 11624 22642 11652 23122
rect 11612 22636 11664 22642
rect 11664 22596 11744 22624
rect 11612 22578 11664 22584
rect 11532 22358 11652 22386
rect 11336 22160 11388 22166
rect 11336 22102 11388 22108
rect 11348 21690 11376 22102
rect 11624 22098 11652 22358
rect 11612 22092 11664 22098
rect 11612 22034 11664 22040
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11244 21140 11296 21146
rect 11244 21082 11296 21088
rect 11624 21078 11652 22034
rect 11716 22001 11744 22596
rect 11808 22234 11836 24670
rect 12176 24614 12204 25230
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 11888 24608 11940 24614
rect 11888 24550 11940 24556
rect 12164 24608 12216 24614
rect 12164 24550 12216 24556
rect 11900 23202 11928 24550
rect 12162 24304 12218 24313
rect 12072 24268 12124 24274
rect 12162 24239 12218 24248
rect 12072 24210 12124 24216
rect 12084 23322 12112 24210
rect 12072 23316 12124 23322
rect 12072 23258 12124 23264
rect 11900 23174 12112 23202
rect 11796 22228 11848 22234
rect 11796 22170 11848 22176
rect 11702 21992 11758 22001
rect 11702 21927 11758 21936
rect 11612 21072 11664 21078
rect 11612 21014 11664 21020
rect 11624 20330 11652 21014
rect 11796 20596 11848 20602
rect 11796 20538 11848 20544
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11612 20324 11664 20330
rect 11612 20266 11664 20272
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 10980 19174 11008 19858
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 10966 19000 11022 19009
rect 10966 18935 11022 18944
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10782 17912 10838 17921
rect 10782 17847 10838 17856
rect 10876 17876 10928 17882
rect 10796 17814 10824 17847
rect 10876 17818 10928 17824
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10690 17232 10746 17241
rect 10888 17202 10916 17818
rect 10690 17167 10692 17176
rect 10744 17167 10746 17176
rect 10876 17196 10928 17202
rect 10692 17138 10744 17144
rect 10876 17138 10928 17144
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10140 16992 10192 16998
rect 10796 16969 10824 17002
rect 10140 16934 10192 16940
rect 10782 16960 10838 16969
rect 10152 16794 10180 16934
rect 10289 16892 10585 16912
rect 10782 16895 10838 16904
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10888 16794 10916 17138
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10980 16658 11008 18935
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 11072 18290 11100 18566
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 11072 17134 11100 17614
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11072 16658 11100 17070
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 11072 16538 11100 16594
rect 10888 16510 11100 16538
rect 10690 16144 10746 16153
rect 10690 16079 10746 16088
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 10152 15745 10180 15914
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10138 15736 10194 15745
rect 10289 15728 10585 15748
rect 10138 15671 10194 15680
rect 10704 15502 10732 16079
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10324 15496 10376 15502
rect 10322 15464 10324 15473
rect 10692 15496 10744 15502
rect 10376 15464 10378 15473
rect 10692 15438 10744 15444
rect 10322 15399 10378 15408
rect 10704 14890 10732 15438
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10046 14512 10102 14521
rect 10046 14447 10048 14456
rect 10100 14447 10102 14456
rect 10048 14418 10100 14424
rect 10152 14414 10180 14826
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14482 10732 14826
rect 10796 14618 10824 15846
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10152 14074 10180 14350
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10690 13560 10746 13569
rect 10690 13495 10692 13504
rect 10744 13495 10746 13504
rect 10692 13466 10744 13472
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 9954 13016 10010 13025
rect 9954 12951 10010 12960
rect 9600 12838 9720 12866
rect 9600 12782 9628 12838
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9956 12640 10008 12646
rect 10060 12628 10088 13194
rect 10152 12918 10180 13262
rect 10244 12986 10272 13262
rect 10704 12986 10732 13466
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10140 12912 10192 12918
rect 10888 12866 10916 16510
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11072 16114 11100 16390
rect 11164 16153 11192 17478
rect 11150 16144 11206 16153
rect 11060 16108 11112 16114
rect 11150 16079 11206 16088
rect 11060 16050 11112 16056
rect 11072 15706 11100 16050
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11164 15638 11192 15846
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 11072 15162 11100 15506
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10966 14784 11022 14793
rect 10966 14719 11022 14728
rect 10980 14618 11008 14719
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11256 13802 11284 19110
rect 11348 17728 11376 19246
rect 11440 18630 11468 19654
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11428 17740 11480 17746
rect 11348 17700 11428 17728
rect 11428 17682 11480 17688
rect 11440 17270 11468 17682
rect 11610 17504 11666 17513
rect 11610 17439 11666 17448
rect 11624 17338 11652 17439
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11440 16250 11468 16594
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11334 16144 11390 16153
rect 11334 16079 11390 16088
rect 11348 15978 11376 16079
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11440 15366 11468 16186
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11716 14929 11744 20402
rect 11808 19689 11836 20538
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 11992 19854 12020 20334
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11794 19680 11850 19689
rect 11794 19615 11850 19624
rect 11992 18970 12020 19790
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 12084 18426 12112 23174
rect 12176 21570 12204 24239
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 12268 23866 12296 24142
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12268 23594 12296 23802
rect 12256 23588 12308 23594
rect 12256 23530 12308 23536
rect 12360 22624 12388 24006
rect 12452 23254 12480 25094
rect 12440 23248 12492 23254
rect 12440 23190 12492 23196
rect 12544 23118 12572 27520
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 12636 25226 12664 25842
rect 12900 25356 12952 25362
rect 12900 25298 12952 25304
rect 12624 25220 12676 25226
rect 12624 25162 12676 25168
rect 12912 24721 12940 25298
rect 12992 24744 13044 24750
rect 12898 24712 12954 24721
rect 12992 24686 13044 24692
rect 12898 24647 12954 24656
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12820 23769 12848 24550
rect 12806 23760 12862 23769
rect 12806 23695 12862 23704
rect 12716 23588 12768 23594
rect 12716 23530 12768 23536
rect 12728 23322 12756 23530
rect 12716 23316 12768 23322
rect 12716 23258 12768 23264
rect 12624 23180 12676 23186
rect 12624 23122 12676 23128
rect 12532 23112 12584 23118
rect 12532 23054 12584 23060
rect 12440 22636 12492 22642
rect 12360 22596 12440 22624
rect 12360 21690 12388 22596
rect 12440 22578 12492 22584
rect 12532 22568 12584 22574
rect 12532 22510 12584 22516
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12452 21729 12480 22374
rect 12438 21720 12494 21729
rect 12348 21684 12400 21690
rect 12438 21655 12494 21664
rect 12348 21626 12400 21632
rect 12176 21542 12296 21570
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 12176 21078 12204 21422
rect 12164 21072 12216 21078
rect 12164 21014 12216 21020
rect 12164 20256 12216 20262
rect 12162 20224 12164 20233
rect 12216 20224 12218 20233
rect 12162 20159 12218 20168
rect 12268 20058 12296 21542
rect 12348 21548 12400 21554
rect 12544 21536 12572 22510
rect 12636 22030 12664 23122
rect 12728 22778 12756 23258
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12820 22574 12848 22918
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 12912 22386 12940 24647
rect 13004 24070 13032 24686
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 13004 23905 13032 24006
rect 12990 23896 13046 23905
rect 12990 23831 13046 23840
rect 12728 22358 12940 22386
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12622 21856 12678 21865
rect 12622 21791 12678 21800
rect 12400 21508 12572 21536
rect 12348 21490 12400 21496
rect 12636 21146 12664 21791
rect 12624 21140 12676 21146
rect 12624 21082 12676 21088
rect 12348 20800 12400 20806
rect 12348 20742 12400 20748
rect 12360 20398 12388 20742
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12256 20052 12308 20058
rect 12176 20012 12256 20040
rect 12176 19446 12204 20012
rect 12256 19994 12308 20000
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12268 19514 12296 19858
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12164 19440 12216 19446
rect 12164 19382 12216 19388
rect 12176 18737 12204 19382
rect 12162 18728 12218 18737
rect 12162 18663 12218 18672
rect 12268 18442 12296 19450
rect 12360 19145 12388 20334
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12452 20097 12480 20198
rect 12438 20088 12494 20097
rect 12636 20058 12664 21082
rect 12438 20023 12494 20032
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12346 19136 12402 19145
rect 12346 19071 12402 19080
rect 12544 18970 12572 19246
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12176 18414 12296 18442
rect 12072 17536 12124 17542
rect 12176 17524 12204 18414
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12268 17746 12296 18226
rect 12360 17882 12388 18566
rect 12544 18426 12572 18770
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 12544 17542 12572 18362
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12124 17496 12204 17524
rect 12532 17536 12584 17542
rect 12072 17478 12124 17484
rect 12532 17478 12584 17484
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11702 14920 11758 14929
rect 11702 14855 11758 14864
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 10140 12854 10192 12860
rect 10008 12600 10088 12628
rect 9956 12582 10008 12588
rect 10060 12442 10088 12600
rect 10704 12838 10916 12866
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10704 12374 10732 12838
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10692 12368 10744 12374
rect 10138 12336 10194 12345
rect 10692 12310 10744 12316
rect 10138 12271 10194 12280
rect 10152 11529 10180 12271
rect 10690 11928 10746 11937
rect 10980 11914 11008 12650
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11072 12306 11100 12582
rect 11164 12374 11192 13126
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10980 11886 11100 11914
rect 11164 11898 11192 12310
rect 11256 12238 11284 12786
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 10690 11863 10746 11872
rect 10138 11520 10194 11529
rect 10138 11455 10194 11464
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11393 10732 11863
rect 11072 11830 11100 11886
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 11256 11762 11284 12174
rect 11348 12170 11376 12650
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11532 12481 11560 12582
rect 11518 12472 11574 12481
rect 11518 12407 11574 12416
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11336 12164 11388 12170
rect 11336 12106 11388 12112
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 10690 11384 10746 11393
rect 11440 11354 11468 12242
rect 10690 11319 10746 11328
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 9494 10704 9550 10713
rect 9494 10639 9550 10648
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 9218 10024 9274 10033
rect 9218 9959 9274 9968
rect 11716 9489 11744 14855
rect 11808 14278 11836 16594
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11900 15570 11928 16050
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11992 14113 12020 14486
rect 11978 14104 12034 14113
rect 11978 14039 12034 14048
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11900 13705 11928 13806
rect 11992 13734 12020 14039
rect 11980 13728 12032 13734
rect 11886 13696 11942 13705
rect 11980 13670 12032 13676
rect 11886 13631 11942 13640
rect 11992 13530 12020 13670
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 11992 12238 12020 13466
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11992 11898 12020 12174
rect 12084 12170 12112 17478
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12176 16182 12204 16934
rect 12544 16454 12572 16934
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 16182 12572 16390
rect 12164 16176 12216 16182
rect 12164 16118 12216 16124
rect 12532 16176 12584 16182
rect 12532 16118 12584 16124
rect 12636 15978 12664 18022
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 15638 12480 15846
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 12176 15162 12204 15302
rect 12360 15162 12388 15574
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12452 15026 12480 15438
rect 12622 15328 12678 15337
rect 12622 15263 12678 15272
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12636 14618 12664 15263
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 12176 13938 12204 14214
rect 12440 14000 12492 14006
rect 12438 13968 12440 13977
rect 12492 13968 12494 13977
rect 12164 13932 12216 13938
rect 12438 13903 12494 13912
rect 12164 13874 12216 13880
rect 12176 13841 12204 13874
rect 12440 13864 12492 13870
rect 12162 13832 12218 13841
rect 12440 13806 12492 13812
rect 12162 13767 12218 13776
rect 12256 13796 12308 13802
rect 12256 13738 12308 13744
rect 12268 13190 12296 13738
rect 12452 13716 12480 13806
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12532 13728 12584 13734
rect 12452 13688 12532 13716
rect 12532 13670 12584 13676
rect 12636 13530 12664 13738
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12728 13410 12756 22358
rect 13096 22273 13124 27520
rect 13452 26172 13504 26178
rect 13452 26114 13504 26120
rect 13266 25392 13322 25401
rect 13322 25336 13400 25344
rect 13266 25327 13268 25336
rect 13320 25316 13400 25336
rect 13268 25298 13320 25304
rect 13372 24886 13400 25316
rect 13360 24880 13412 24886
rect 13360 24822 13412 24828
rect 13268 24608 13320 24614
rect 13320 24568 13400 24596
rect 13268 24550 13320 24556
rect 13266 23352 13322 23361
rect 13266 23287 13322 23296
rect 13082 22264 13138 22273
rect 13280 22234 13308 23287
rect 13082 22199 13138 22208
rect 13268 22228 13320 22234
rect 13268 22170 13320 22176
rect 12900 22160 12952 22166
rect 12900 22102 12952 22108
rect 13084 22160 13136 22166
rect 13084 22102 13136 22108
rect 12820 20534 12848 20565
rect 12808 20528 12860 20534
rect 12806 20496 12808 20505
rect 12860 20496 12862 20505
rect 12806 20431 12862 20440
rect 12820 20398 12848 20431
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12806 20224 12862 20233
rect 12806 20159 12862 20168
rect 12820 18902 12848 20159
rect 12912 19174 12940 22102
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 13004 20466 13032 21830
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 13004 19854 13032 20402
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 13096 19310 13124 22102
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13188 21350 13216 21966
rect 13176 21344 13228 21350
rect 13176 21286 13228 21292
rect 13266 21312 13322 21321
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12820 17610 12848 18022
rect 12808 17604 12860 17610
rect 12808 17546 12860 17552
rect 13004 17134 13032 18838
rect 13096 18057 13124 19110
rect 13082 18048 13138 18057
rect 13082 17983 13138 17992
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 13004 16833 13032 17070
rect 13082 16960 13138 16969
rect 13082 16895 13138 16904
rect 12990 16824 13046 16833
rect 12990 16759 13046 16768
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 12912 15570 12940 16526
rect 13096 15978 13124 16895
rect 13084 15972 13136 15978
rect 13084 15914 13136 15920
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12912 15201 12940 15506
rect 12898 15192 12954 15201
rect 12898 15127 12954 15136
rect 13004 15042 13032 15846
rect 13096 15366 13124 15914
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 12912 15014 13032 15042
rect 12808 14816 12860 14822
rect 12806 14784 12808 14793
rect 12860 14784 12862 14793
rect 12806 14719 12862 14728
rect 12820 14618 12848 14719
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12544 13382 12756 13410
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12268 12442 12296 13126
rect 12452 12646 12480 13330
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12360 11354 12388 11698
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 11702 9480 11758 9489
rect 11702 9415 11758 9424
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 9586 9072 9642 9081
rect 9586 9007 9642 9016
rect 9600 8634 9628 9007
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 9586 6216 9642 6225
rect 9586 6151 9642 6160
rect 9600 5914 9628 6151
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 8850 3632 8906 3641
rect 8850 3567 8906 3576
rect 12452 3505 12480 12582
rect 12544 11354 12572 13382
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12636 11898 12664 13262
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12820 11257 12848 14350
rect 12806 11248 12862 11257
rect 12806 11183 12862 11192
rect 12438 3496 12494 3505
rect 12438 3431 12494 3440
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 8298 2952 8354 2961
rect 8298 2887 8354 2896
rect 12438 2952 12494 2961
rect 12438 2887 12494 2896
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 8312 480 8340 2887
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 12452 2650 12480 2887
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12714 2544 12770 2553
rect 12714 2479 12716 2488
rect 12768 2479 12770 2488
rect 12716 2450 12768 2456
rect 4066 368 4122 377
rect 4066 303 4122 312
rect 8298 0 8354 480
rect 12912 105 12940 15014
rect 12990 13696 13046 13705
rect 12990 13631 13046 13640
rect 13004 12442 13032 13631
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12990 12064 13046 12073
rect 12990 11999 13046 12008
rect 13004 9625 13032 11999
rect 13096 11642 13124 15302
rect 13188 12073 13216 21286
rect 13266 21247 13322 21256
rect 13280 18426 13308 21247
rect 13372 21185 13400 24568
rect 13464 22506 13492 26114
rect 13648 24562 13676 27520
rect 14188 25356 14240 25362
rect 14188 25298 14240 25304
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 13556 24534 13676 24562
rect 13556 24177 13584 24534
rect 13634 24440 13690 24449
rect 14108 24410 14136 25094
rect 13634 24375 13636 24384
rect 13688 24375 13690 24384
rect 14096 24404 14148 24410
rect 13636 24346 13688 24352
rect 14096 24346 14148 24352
rect 13542 24168 13598 24177
rect 13542 24103 13598 24112
rect 13648 23322 13676 24346
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 13728 24064 13780 24070
rect 14108 24052 14136 24210
rect 14200 24206 14228 25298
rect 14292 24834 14320 27520
rect 14844 24834 14872 27520
rect 15396 25242 15424 27520
rect 15304 25214 15424 25242
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14924 24880 14976 24886
rect 14292 24806 14504 24834
rect 14370 24712 14426 24721
rect 14370 24647 14372 24656
rect 14424 24647 14426 24656
rect 14372 24618 14424 24624
rect 14280 24608 14332 24614
rect 14280 24550 14332 24556
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14108 24024 14228 24052
rect 13728 24006 13780 24012
rect 13740 23322 13768 24006
rect 14200 23526 14228 24024
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 14188 23520 14240 23526
rect 14188 23462 14240 23468
rect 13636 23316 13688 23322
rect 13636 23258 13688 23264
rect 13728 23316 13780 23322
rect 13728 23258 13780 23264
rect 13740 23202 13768 23258
rect 13556 23174 13768 23202
rect 13452 22500 13504 22506
rect 13452 22442 13504 22448
rect 13556 22166 13584 23174
rect 13636 23112 13688 23118
rect 13636 23054 13688 23060
rect 13726 23080 13782 23089
rect 13544 22160 13596 22166
rect 13544 22102 13596 22108
rect 13450 21992 13506 22001
rect 13450 21927 13506 21936
rect 13358 21176 13414 21185
rect 13464 21146 13492 21927
rect 13542 21720 13598 21729
rect 13542 21655 13598 21664
rect 13358 21111 13414 21120
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13372 20754 13400 20946
rect 13464 20942 13492 21082
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13372 20726 13492 20754
rect 13358 20632 13414 20641
rect 13358 20567 13414 20576
rect 13372 19990 13400 20567
rect 13464 20262 13492 20726
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 13372 19310 13400 19926
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13268 18420 13320 18426
rect 13268 18362 13320 18368
rect 13464 18154 13492 20198
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13358 17640 13414 17649
rect 13280 16658 13308 17614
rect 13358 17575 13360 17584
rect 13412 17575 13414 17584
rect 13360 17546 13412 17552
rect 13464 17377 13492 17682
rect 13450 17368 13506 17377
rect 13450 17303 13452 17312
rect 13504 17303 13506 17312
rect 13452 17274 13504 17280
rect 13464 17243 13492 17274
rect 13556 16697 13584 21655
rect 13542 16688 13598 16697
rect 13268 16652 13320 16658
rect 13542 16623 13544 16632
rect 13268 16594 13320 16600
rect 13596 16623 13598 16632
rect 13544 16594 13596 16600
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13372 13569 13400 15846
rect 13464 15706 13492 16390
rect 13556 16250 13584 16594
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13464 15502 13492 15642
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13556 15162 13584 16050
rect 13648 15910 13676 23054
rect 13726 23015 13782 23024
rect 13740 21554 13768 23015
rect 13832 22642 13860 23462
rect 14096 23112 14148 23118
rect 14200 23089 14228 23462
rect 14096 23054 14148 23060
rect 14186 23080 14242 23089
rect 14108 22778 14136 23054
rect 14186 23015 14242 23024
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 14200 22681 14228 23015
rect 14186 22672 14242 22681
rect 13820 22636 13872 22642
rect 14186 22607 14242 22616
rect 13820 22578 13872 22584
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 13820 22500 13872 22506
rect 13820 22442 13872 22448
rect 13832 22234 13860 22442
rect 13820 22228 13872 22234
rect 13820 22170 13872 22176
rect 13912 22024 13964 22030
rect 13910 21992 13912 22001
rect 14004 22024 14056 22030
rect 13964 21992 13966 22001
rect 14004 21966 14056 21972
rect 13910 21927 13966 21936
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13820 21072 13872 21078
rect 13740 21032 13820 21060
rect 13740 20058 13768 21032
rect 13820 21014 13872 21020
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 13832 20602 13860 20878
rect 13924 20806 13952 21830
rect 14016 21350 14044 21966
rect 14108 21350 14136 22510
rect 14292 21962 14320 24550
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14384 22098 14412 22918
rect 14372 22092 14424 22098
rect 14372 22034 14424 22040
rect 14280 21956 14332 21962
rect 14280 21898 14332 21904
rect 14292 21418 14320 21898
rect 14280 21412 14332 21418
rect 14280 21354 14332 21360
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 14096 21344 14148 21350
rect 14476 21321 14504 24806
rect 14568 24806 14872 24834
rect 14922 24848 14924 24857
rect 14976 24848 14978 24857
rect 14568 21865 14596 24806
rect 14922 24783 14978 24792
rect 15106 24848 15162 24857
rect 15106 24783 15162 24792
rect 15120 24614 15148 24783
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 15304 24426 15332 25214
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 15212 24398 15332 24426
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14554 21856 14610 21865
rect 14554 21791 14610 21800
rect 14660 21570 14688 24142
rect 14740 24132 14792 24138
rect 14740 24074 14792 24080
rect 14752 23526 14780 24074
rect 14844 23730 14872 24346
rect 15212 24313 15240 24398
rect 15198 24304 15254 24313
rect 15198 24239 15254 24248
rect 15292 24268 15344 24274
rect 15292 24210 15344 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15304 23848 15332 24210
rect 15396 24052 15424 25094
rect 15580 24614 15608 25230
rect 15660 25152 15712 25158
rect 15660 25094 15712 25100
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 15474 24440 15530 24449
rect 15474 24375 15476 24384
rect 15528 24375 15530 24384
rect 15476 24346 15528 24352
rect 15476 24064 15528 24070
rect 15396 24024 15476 24052
rect 15476 24006 15528 24012
rect 15120 23820 15332 23848
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 14740 23520 14792 23526
rect 14740 23462 14792 23468
rect 14752 22438 14780 23462
rect 15120 23322 15148 23820
rect 15488 23594 15516 24006
rect 15476 23588 15528 23594
rect 15476 23530 15528 23536
rect 15488 23322 15516 23530
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 15476 23316 15528 23322
rect 15476 23258 15528 23264
rect 15292 23112 15344 23118
rect 15580 23066 15608 24550
rect 15672 24274 15700 25094
rect 15948 24834 15976 27520
rect 16500 25378 16528 27520
rect 16854 25800 16910 25809
rect 16854 25735 16910 25744
rect 16316 25350 16528 25378
rect 16580 25356 16632 25362
rect 15948 24806 16252 24834
rect 15750 24712 15806 24721
rect 15750 24647 15806 24656
rect 15660 24268 15712 24274
rect 15660 24210 15712 24216
rect 15658 24168 15714 24177
rect 15658 24103 15714 24112
rect 15292 23054 15344 23060
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14740 22432 14792 22438
rect 14740 22374 14792 22380
rect 14752 22001 14780 22374
rect 15304 22273 15332 23054
rect 15488 23038 15608 23066
rect 15384 22500 15436 22506
rect 15384 22442 15436 22448
rect 15290 22264 15346 22273
rect 15290 22199 15346 22208
rect 14738 21992 14794 22001
rect 14738 21927 14794 21936
rect 14832 21956 14884 21962
rect 14832 21898 14884 21904
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14568 21542 14688 21570
rect 14096 21286 14148 21292
rect 14462 21312 14518 21321
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13832 19514 13860 20266
rect 13924 20233 13952 20742
rect 13910 20224 13966 20233
rect 13910 20159 13966 20168
rect 14016 20074 14044 21286
rect 14108 20398 14136 21286
rect 14462 21247 14518 21256
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 13924 20046 14044 20074
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 13832 18970 13860 19178
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13740 17649 13768 18770
rect 13832 18426 13860 18906
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 13726 17640 13782 17649
rect 13726 17575 13782 17584
rect 13832 17241 13860 17750
rect 13818 17232 13874 17241
rect 13818 17167 13874 17176
rect 13924 17082 13952 20046
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 14016 18630 14044 19790
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 14016 18290 14044 18566
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13832 17054 13952 17082
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13740 16232 13768 16730
rect 13832 16561 13860 17054
rect 14016 16998 14044 18226
rect 14108 18057 14136 19858
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14200 18086 14228 18226
rect 14188 18080 14240 18086
rect 14094 18048 14150 18057
rect 14188 18022 14240 18028
rect 14094 17983 14150 17992
rect 14200 17785 14228 18022
rect 14186 17776 14242 17785
rect 14186 17711 14242 17720
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 13912 16584 13964 16590
rect 13818 16552 13874 16561
rect 13912 16526 13964 16532
rect 13818 16487 13874 16496
rect 13820 16244 13872 16250
rect 13740 16204 13820 16232
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13648 15162 13676 15438
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13556 14482 13584 15098
rect 13740 14958 13768 16204
rect 13820 16186 13872 16192
rect 13924 16114 13952 16526
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 14016 15994 14044 16934
rect 13924 15966 14044 15994
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13740 14414 13768 14486
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13820 13728 13872 13734
rect 13818 13696 13820 13705
rect 13872 13696 13874 13705
rect 13818 13631 13874 13640
rect 13358 13560 13414 13569
rect 13358 13495 13414 13504
rect 13818 13288 13874 13297
rect 13818 13223 13820 13232
rect 13872 13223 13874 13232
rect 13820 13194 13872 13200
rect 13266 12880 13322 12889
rect 13266 12815 13322 12824
rect 13280 12782 13308 12815
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13174 12064 13230 12073
rect 13174 11999 13230 12008
rect 13096 11614 13216 11642
rect 13084 11552 13136 11558
rect 13082 11520 13084 11529
rect 13136 11520 13138 11529
rect 13082 11455 13138 11464
rect 13096 11286 13124 11455
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 13096 11121 13124 11222
rect 13188 11150 13216 11614
rect 13176 11144 13228 11150
rect 13082 11112 13138 11121
rect 13176 11086 13228 11092
rect 13082 11047 13138 11056
rect 13188 10962 13216 11086
rect 13096 10934 13216 10962
rect 13096 10470 13124 10934
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12990 9616 13046 9625
rect 12990 9551 13046 9560
rect 13096 3505 13124 10406
rect 13280 5545 13308 12106
rect 13372 11830 13400 12242
rect 13556 12238 13584 12582
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13464 11558 13492 12038
rect 13556 11762 13584 12174
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13740 11694 13768 12242
rect 13728 11688 13780 11694
rect 13726 11656 13728 11665
rect 13780 11656 13782 11665
rect 13726 11591 13782 11600
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 11286 13492 11494
rect 13452 11280 13504 11286
rect 13452 11222 13504 11228
rect 13464 10470 13492 11222
rect 13728 11144 13780 11150
rect 13924 11132 13952 15966
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14016 14113 14044 14214
rect 14002 14104 14058 14113
rect 14002 14039 14058 14048
rect 14016 13938 14044 14039
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 14108 12617 14136 17274
rect 14292 13569 14320 20878
rect 14476 20777 14504 21247
rect 14462 20768 14518 20777
rect 14462 20703 14518 20712
rect 14370 20224 14426 20233
rect 14370 20159 14426 20168
rect 14384 19553 14412 20159
rect 14462 20088 14518 20097
rect 14462 20023 14518 20032
rect 14476 19825 14504 20023
rect 14462 19816 14518 19825
rect 14462 19751 14518 19760
rect 14370 19544 14426 19553
rect 14370 19479 14426 19488
rect 14462 18864 14518 18873
rect 14462 18799 14464 18808
rect 14516 18799 14518 18808
rect 14464 18770 14516 18776
rect 14370 18592 14426 18601
rect 14370 18527 14426 18536
rect 14384 18426 14412 18527
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14476 18222 14504 18770
rect 14464 18216 14516 18222
rect 14370 18184 14426 18193
rect 14464 18158 14516 18164
rect 14370 18119 14426 18128
rect 14384 18086 14412 18119
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14462 18048 14518 18057
rect 14384 17882 14412 18022
rect 14462 17983 14518 17992
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14476 17762 14504 17983
rect 14568 17921 14596 21542
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14660 20398 14688 21422
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14660 20058 14688 20334
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14660 19281 14688 19654
rect 14646 19272 14702 19281
rect 14646 19207 14702 19216
rect 14752 19009 14780 21830
rect 14844 21690 14872 21898
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 15292 21412 15344 21418
rect 15292 21354 15344 21360
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14844 20602 14872 20742
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14738 19000 14794 19009
rect 14648 18964 14700 18970
rect 15304 18986 15332 21354
rect 15396 20534 15424 22442
rect 15488 21418 15516 23038
rect 15672 22710 15700 24103
rect 15660 22704 15712 22710
rect 15660 22646 15712 22652
rect 15660 22024 15712 22030
rect 15566 21992 15622 22001
rect 15660 21966 15712 21972
rect 15566 21927 15622 21936
rect 15476 21412 15528 21418
rect 15476 21354 15528 21360
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15384 20528 15436 20534
rect 15384 20470 15436 20476
rect 15384 20324 15436 20330
rect 15384 20266 15436 20272
rect 15396 19922 15424 20266
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15396 19156 15424 19858
rect 15488 19718 15516 20878
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15476 19168 15528 19174
rect 15396 19128 15476 19156
rect 15476 19110 15528 19116
rect 15304 18958 15516 18986
rect 14738 18935 14794 18944
rect 14648 18906 14700 18912
rect 14660 18873 14688 18906
rect 14646 18864 14702 18873
rect 14646 18799 14702 18808
rect 15384 18828 15436 18834
rect 14554 17912 14610 17921
rect 14554 17847 14610 17856
rect 14476 17734 14596 17762
rect 14462 16552 14518 16561
rect 14462 16487 14518 16496
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 14384 15706 14412 16050
rect 14476 16046 14504 16487
rect 14568 16266 14596 17734
rect 14660 17134 14688 18799
rect 15384 18770 15436 18776
rect 15396 18737 15424 18770
rect 15382 18728 15438 18737
rect 15382 18663 15438 18672
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14738 17912 14794 17921
rect 14738 17847 14794 17856
rect 14752 17814 14780 17847
rect 14740 17808 14792 17814
rect 14740 17750 14792 17756
rect 14752 17338 14780 17750
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14844 17202 14872 17478
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15106 17232 15162 17241
rect 14832 17196 14884 17202
rect 15106 17167 15108 17176
rect 14832 17138 14884 17144
rect 15160 17167 15162 17176
rect 15108 17138 15160 17144
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 15014 17096 15070 17105
rect 14660 16794 14688 17070
rect 15014 17031 15016 17040
rect 15068 17031 15070 17040
rect 15016 17002 15068 17008
rect 15028 16794 15056 17002
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15382 16280 15438 16289
rect 14568 16238 14872 16266
rect 14554 16144 14610 16153
rect 14554 16079 14610 16088
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14476 15570 14504 15982
rect 14568 15978 14596 16079
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14554 15600 14610 15609
rect 14464 15564 14516 15570
rect 14554 15535 14610 15544
rect 14464 15506 14516 15512
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14384 13870 14412 14894
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14278 13560 14334 13569
rect 14278 13495 14334 13504
rect 14280 13456 14332 13462
rect 14280 13398 14332 13404
rect 14094 12608 14150 12617
rect 14094 12543 14150 12552
rect 14292 12306 14320 13398
rect 14384 12986 14412 13806
rect 14568 13462 14596 15535
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14660 13870 14688 14214
rect 14752 14074 14780 14826
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14384 12102 14412 12922
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 13780 11104 13952 11132
rect 13728 11086 13780 11092
rect 13740 10810 13768 11086
rect 14108 11082 14136 12038
rect 14568 11898 14596 13126
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14660 11642 14688 13806
rect 14752 12442 14780 14010
rect 14844 12481 14872 16238
rect 15488 16266 15516 18958
rect 15580 18426 15608 21927
rect 15672 20330 15700 21966
rect 15660 20324 15712 20330
rect 15660 20266 15712 20272
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15672 18766 15700 19110
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15580 17746 15608 18362
rect 15764 17882 15792 24647
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 16028 24608 16080 24614
rect 16028 24550 16080 24556
rect 15948 24206 15976 24550
rect 15936 24200 15988 24206
rect 15936 24142 15988 24148
rect 15844 24132 15896 24138
rect 15844 24074 15896 24080
rect 15856 23866 15884 24074
rect 15948 23866 15976 24142
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 15856 23526 15884 23802
rect 15844 23520 15896 23526
rect 15844 23462 15896 23468
rect 15856 22778 15884 23462
rect 15936 23180 15988 23186
rect 15936 23122 15988 23128
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15856 21622 15884 22374
rect 15948 22030 15976 23122
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15948 21690 15976 21830
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 15844 21616 15896 21622
rect 15844 21558 15896 21564
rect 16040 21536 16068 24550
rect 16120 23248 16172 23254
rect 16120 23190 16172 23196
rect 15948 21508 16068 21536
rect 15844 21344 15896 21350
rect 15842 21312 15844 21321
rect 15896 21312 15898 21321
rect 15842 21247 15898 21256
rect 15842 20904 15898 20913
rect 15842 20839 15844 20848
rect 15896 20839 15898 20848
rect 15844 20810 15896 20816
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 15856 19310 15884 19858
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15856 17202 15884 19246
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15438 16238 15516 16266
rect 15382 16215 15438 16224
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 14958 15332 15438
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15304 14657 15332 14894
rect 15290 14648 15346 14657
rect 15290 14583 15346 14592
rect 15396 14550 15424 16215
rect 15764 16114 15792 16594
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15948 15994 15976 21508
rect 16132 21468 16160 23190
rect 16040 21440 16160 21468
rect 16040 18902 16068 21440
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 16132 21146 16160 21286
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 16132 20262 16160 20878
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16028 18896 16080 18902
rect 16028 18838 16080 18844
rect 16132 17785 16160 20198
rect 16224 17921 16252 24806
rect 16316 21962 16344 25350
rect 16580 25298 16632 25304
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 16408 24698 16436 25230
rect 16488 24744 16540 24750
rect 16408 24692 16488 24698
rect 16408 24686 16540 24692
rect 16408 24670 16528 24686
rect 16396 24608 16448 24614
rect 16396 24550 16448 24556
rect 16408 24449 16436 24550
rect 16394 24440 16450 24449
rect 16394 24375 16450 24384
rect 16396 24336 16448 24342
rect 16396 24278 16448 24284
rect 16408 23186 16436 24278
rect 16500 23322 16528 24670
rect 16592 24410 16620 25298
rect 16672 25152 16724 25158
rect 16672 25094 16724 25100
rect 16580 24404 16632 24410
rect 16580 24346 16632 24352
rect 16684 24342 16712 25094
rect 16868 24993 16896 25735
rect 17052 25294 17080 27520
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 17224 25220 17276 25226
rect 17224 25162 17276 25168
rect 16854 24984 16910 24993
rect 17236 24954 17264 25162
rect 16854 24919 16910 24928
rect 17224 24948 17276 24954
rect 16672 24336 16724 24342
rect 16672 24278 16724 24284
rect 16580 23520 16632 23526
rect 16580 23462 16632 23468
rect 16488 23316 16540 23322
rect 16488 23258 16540 23264
rect 16396 23180 16448 23186
rect 16396 23122 16448 23128
rect 16500 23066 16528 23258
rect 16592 23254 16620 23462
rect 16580 23248 16632 23254
rect 16580 23190 16632 23196
rect 16500 23038 16620 23066
rect 16396 22704 16448 22710
rect 16396 22646 16448 22652
rect 16304 21956 16356 21962
rect 16304 21898 16356 21904
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16316 21350 16344 21626
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16316 19990 16344 21286
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16408 19258 16436 22646
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 16500 20380 16528 22374
rect 16592 21894 16620 23038
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16684 22438 16712 22918
rect 16672 22432 16724 22438
rect 16670 22400 16672 22409
rect 16724 22400 16726 22409
rect 16670 22335 16726 22344
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16580 20392 16632 20398
rect 16500 20352 16580 20380
rect 16580 20334 16632 20340
rect 16684 20058 16712 21422
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16868 19904 16896 24919
rect 17224 24890 17276 24896
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 17052 22098 17080 24550
rect 17314 24032 17370 24041
rect 17314 23967 17370 23976
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16960 21078 16988 21286
rect 16948 21072 17000 21078
rect 16948 21014 17000 21020
rect 16960 20330 16988 21014
rect 17052 21010 17080 22034
rect 17040 21004 17092 21010
rect 17040 20946 17092 20952
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 16592 19876 16896 19904
rect 16316 19145 16344 19246
rect 16408 19230 16528 19258
rect 16396 19168 16448 19174
rect 16302 19136 16358 19145
rect 16396 19110 16448 19116
rect 16302 19071 16358 19080
rect 16408 19009 16436 19110
rect 16394 19000 16450 19009
rect 16394 18935 16450 18944
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16408 18193 16436 18702
rect 16394 18184 16450 18193
rect 16394 18119 16450 18128
rect 16210 17912 16266 17921
rect 16210 17847 16266 17856
rect 16118 17776 16174 17785
rect 16118 17711 16174 17720
rect 16302 17776 16358 17785
rect 16302 17711 16304 17720
rect 16132 17377 16160 17711
rect 16356 17711 16358 17720
rect 16304 17682 16356 17688
rect 16118 17368 16174 17377
rect 16118 17303 16174 17312
rect 16210 17096 16266 17105
rect 16316 17066 16344 17682
rect 16408 17678 16436 18119
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16210 17031 16266 17040
rect 16304 17060 16356 17066
rect 16224 16998 16252 17031
rect 16304 17002 16356 17008
rect 16212 16992 16264 16998
rect 16408 16946 16436 17614
rect 16212 16934 16264 16940
rect 16316 16918 16436 16946
rect 16316 16726 16344 16918
rect 16394 16824 16450 16833
rect 16394 16759 16450 16768
rect 16304 16720 16356 16726
rect 16304 16662 16356 16668
rect 15948 15966 16252 15994
rect 15568 15904 15620 15910
rect 15936 15904 15988 15910
rect 15568 15846 15620 15852
rect 15750 15872 15806 15881
rect 15580 15473 15608 15846
rect 15936 15846 15988 15852
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 15750 15807 15806 15816
rect 15764 15473 15792 15807
rect 15844 15564 15896 15570
rect 15844 15506 15896 15512
rect 15566 15464 15622 15473
rect 15566 15399 15622 15408
rect 15750 15464 15806 15473
rect 15750 15399 15806 15408
rect 15856 14822 15884 15506
rect 15948 15366 15976 15846
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14830 12472 14886 12481
rect 14740 12436 14792 12442
rect 14830 12407 14886 12416
rect 14740 12378 14792 12384
rect 14752 11762 14780 12378
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14292 11614 14688 11642
rect 14738 11656 14794 11665
rect 14292 11121 14320 11614
rect 14738 11591 14740 11600
rect 14792 11591 14794 11600
rect 14740 11562 14792 11568
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14278 11112 14334 11121
rect 14096 11076 14148 11082
rect 14278 11047 14334 11056
rect 14096 11018 14148 11024
rect 14292 10962 14320 11047
rect 14108 10934 14320 10962
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13464 10169 13492 10406
rect 13450 10160 13506 10169
rect 13450 10095 13506 10104
rect 13266 5536 13322 5545
rect 13266 5471 13322 5480
rect 13726 5128 13782 5137
rect 13726 5063 13782 5072
rect 13740 4049 13768 5063
rect 13726 4040 13782 4049
rect 13726 3975 13782 3984
rect 13910 3632 13966 3641
rect 13910 3567 13966 3576
rect 13082 3496 13138 3505
rect 13082 3431 13138 3440
rect 13924 480 13952 3567
rect 14108 2650 14136 10934
rect 14384 5681 14412 11494
rect 14752 11218 14780 11562
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14660 10470 14688 11018
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14554 9616 14610 9625
rect 14554 9551 14610 9560
rect 14370 5672 14426 5681
rect 14370 5607 14426 5616
rect 14186 5536 14242 5545
rect 14186 5471 14242 5480
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14200 1465 14228 5471
rect 14568 5273 14596 9551
rect 14554 5264 14610 5273
rect 14554 5199 14610 5208
rect 14660 2553 14688 10406
rect 14752 9081 14780 11154
rect 14738 9072 14794 9081
rect 14738 9007 14794 9016
rect 14844 3641 14872 12407
rect 15304 12306 15332 14350
rect 15856 14278 15884 14758
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15752 13456 15804 13462
rect 15752 13398 15804 13404
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15580 11286 15608 12242
rect 15672 11354 15700 12582
rect 15764 12442 15792 13398
rect 15856 13326 15884 14214
rect 15948 13530 15976 15302
rect 16132 14822 16160 15846
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15856 12850 15884 13262
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15764 11665 15792 12174
rect 15750 11656 15806 11665
rect 15750 11591 15752 11600
rect 15804 11591 15806 11600
rect 15752 11562 15804 11568
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 16040 11218 16068 14010
rect 16132 12986 16160 14758
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 16132 11898 16160 12650
rect 16224 12345 16252 15966
rect 16408 15638 16436 16759
rect 16396 15632 16448 15638
rect 16396 15574 16448 15580
rect 16408 14618 16436 15574
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16500 14550 16528 19230
rect 16592 14618 16620 19876
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16776 19310 16804 19722
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16868 18970 16896 19110
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 16960 18834 16988 19314
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16960 18426 16988 18770
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16960 18290 16988 18362
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16868 16794 16896 18022
rect 16946 17912 17002 17921
rect 16946 17847 17002 17856
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16764 16720 16816 16726
rect 16816 16668 16896 16674
rect 16764 16662 16896 16668
rect 16776 16646 16896 16662
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16684 15910 16712 16050
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16684 15706 16712 15846
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16488 14544 16540 14550
rect 16488 14486 16540 14492
rect 16302 14376 16358 14385
rect 16302 14311 16304 14320
rect 16356 14311 16358 14320
rect 16304 14282 16356 14288
rect 16500 14074 16528 14486
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16488 13524 16540 13530
rect 16592 13512 16620 14554
rect 16684 14521 16712 14758
rect 16670 14512 16726 14521
rect 16670 14447 16726 14456
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16776 13530 16804 14350
rect 16868 13818 16896 16646
rect 16960 13938 16988 17847
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17040 16516 17092 16522
rect 17040 16458 17092 16464
rect 17052 16250 17080 16458
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 17130 16144 17186 16153
rect 17130 16079 17186 16088
rect 17038 15192 17094 15201
rect 17038 15127 17040 15136
rect 17092 15127 17094 15136
rect 17040 15098 17092 15104
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16868 13790 16988 13818
rect 16854 13696 16910 13705
rect 16854 13631 16910 13640
rect 16868 13530 16896 13631
rect 16540 13484 16620 13512
rect 16764 13524 16816 13530
rect 16488 13466 16540 13472
rect 16764 13466 16816 13472
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16210 12336 16266 12345
rect 16210 12271 16266 12280
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16316 11830 16344 12174
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16120 11280 16172 11286
rect 16120 11222 16172 11228
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15396 10810 15424 11154
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15764 10810 15792 11086
rect 16132 10810 16160 11222
rect 16316 11150 16344 11766
rect 16500 11762 16528 13466
rect 16762 13016 16818 13025
rect 16762 12951 16818 12960
rect 16776 12850 16804 12951
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 16408 4593 16436 11494
rect 16500 11354 16528 11698
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16868 11286 16896 12038
rect 16960 11354 16988 13790
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16854 11112 16910 11121
rect 16854 11047 16856 11056
rect 16908 11047 16910 11056
rect 16856 11018 16908 11024
rect 17144 10985 17172 16079
rect 17236 16017 17264 16526
rect 17222 16008 17278 16017
rect 17222 15943 17224 15952
rect 17276 15943 17278 15952
rect 17224 15914 17276 15920
rect 17328 15570 17356 23967
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17512 23322 17540 23462
rect 17500 23316 17552 23322
rect 17500 23258 17552 23264
rect 17406 22536 17462 22545
rect 17406 22471 17408 22480
rect 17460 22471 17462 22480
rect 17408 22442 17460 22448
rect 17604 22148 17632 27520
rect 18156 26246 18184 27520
rect 18144 26240 18196 26246
rect 18144 26182 18196 26188
rect 18708 25838 18736 27520
rect 18696 25832 18748 25838
rect 18696 25774 18748 25780
rect 19260 25702 19288 27520
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 19248 25696 19300 25702
rect 19248 25638 19300 25644
rect 18788 25356 18840 25362
rect 18788 25298 18840 25304
rect 18052 25288 18104 25294
rect 18052 25230 18104 25236
rect 18064 24954 18092 25230
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18052 24948 18104 24954
rect 18104 24908 18276 24936
rect 18052 24890 18104 24896
rect 18052 24268 18104 24274
rect 18052 24210 18104 24216
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 17880 23633 17908 24142
rect 17866 23624 17922 23633
rect 17866 23559 17922 23568
rect 18064 22778 18092 24210
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 18064 22273 18092 22374
rect 18050 22264 18106 22273
rect 18050 22199 18052 22208
rect 18104 22199 18106 22208
rect 18052 22170 18104 22176
rect 17512 22120 17632 22148
rect 17512 19446 17540 22120
rect 18248 22080 18276 24908
rect 18616 24818 18644 25094
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18800 24614 18828 25298
rect 19156 25288 19208 25294
rect 19156 25230 19208 25236
rect 18604 24608 18656 24614
rect 18604 24550 18656 24556
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18524 23322 18552 24142
rect 18616 24070 18644 24550
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18328 23316 18380 23322
rect 18328 23258 18380 23264
rect 18512 23316 18564 23322
rect 18512 23258 18564 23264
rect 18340 22642 18368 23258
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18340 22234 18368 22578
rect 18524 22234 18552 23258
rect 18328 22228 18380 22234
rect 18328 22170 18380 22176
rect 18512 22228 18564 22234
rect 18512 22170 18564 22176
rect 18156 22052 18276 22080
rect 17776 22024 17828 22030
rect 17776 21966 17828 21972
rect 17788 21622 17816 21966
rect 17776 21616 17828 21622
rect 17774 21584 17776 21593
rect 17828 21584 17830 21593
rect 17830 21542 17908 21570
rect 17774 21519 17830 21528
rect 17592 21412 17644 21418
rect 17592 21354 17644 21360
rect 17604 21185 17632 21354
rect 17590 21176 17646 21185
rect 17590 21111 17646 21120
rect 17604 21078 17632 21111
rect 17592 21072 17644 21078
rect 17592 21014 17644 21020
rect 17774 20360 17830 20369
rect 17774 20295 17830 20304
rect 17788 20058 17816 20295
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 17880 19922 17908 21542
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17972 20466 18000 20742
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17500 19440 17552 19446
rect 17500 19382 17552 19388
rect 17604 18601 17632 19450
rect 17788 18850 17816 19654
rect 17880 19514 17908 19858
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17972 19174 18000 19382
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17696 18834 18000 18850
rect 17696 18828 18012 18834
rect 17696 18822 17960 18828
rect 17590 18592 17646 18601
rect 17590 18527 17646 18536
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17512 18086 17540 18226
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17512 17882 17540 18022
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17696 17746 17724 18822
rect 17960 18770 18012 18776
rect 17776 18216 17828 18222
rect 17776 18158 17828 18164
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17696 17270 17724 17682
rect 17788 17338 17816 18158
rect 17868 18148 17920 18154
rect 17868 18090 17920 18096
rect 17880 17864 17908 18090
rect 17960 17876 18012 17882
rect 17880 17836 17960 17864
rect 17960 17818 18012 17824
rect 18064 17814 18092 20198
rect 18156 19242 18184 22052
rect 18512 21616 18564 21622
rect 18512 21558 18564 21564
rect 18524 21457 18552 21558
rect 18510 21448 18566 21457
rect 18510 21383 18566 21392
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18432 21146 18460 21286
rect 18420 21140 18472 21146
rect 18420 21082 18472 21088
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18248 19281 18276 19994
rect 18432 19990 18460 20198
rect 18420 19984 18472 19990
rect 18420 19926 18472 19932
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18340 19310 18368 19654
rect 18328 19304 18380 19310
rect 18234 19272 18290 19281
rect 18144 19236 18196 19242
rect 18328 19246 18380 19252
rect 18234 19207 18290 19216
rect 18144 19178 18196 19184
rect 18248 18902 18276 19207
rect 18236 18896 18288 18902
rect 18236 18838 18288 18844
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18156 18290 18184 18566
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18052 17808 18104 17814
rect 18052 17750 18104 17756
rect 18064 17338 18092 17750
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 17684 17264 17736 17270
rect 17684 17206 17736 17212
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17420 15706 17448 16390
rect 17682 16008 17738 16017
rect 17682 15943 17738 15952
rect 17696 15706 17724 15943
rect 17788 15910 17816 16526
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17222 15464 17278 15473
rect 17222 15399 17278 15408
rect 17236 15026 17264 15399
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17236 12220 17264 14962
rect 17328 14618 17356 15506
rect 17788 15337 17816 15846
rect 17774 15328 17830 15337
rect 17774 15263 17830 15272
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17788 14657 17816 14894
rect 17774 14648 17830 14657
rect 17316 14612 17368 14618
rect 17774 14583 17830 14592
rect 17316 14554 17368 14560
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17604 14414 17632 14486
rect 17788 14414 17816 14583
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 17604 14074 17632 14350
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 17420 13870 17448 13942
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17420 13530 17448 13806
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17498 13288 17554 13297
rect 17788 13258 17816 14350
rect 17880 14074 17908 15098
rect 18064 14958 18092 15982
rect 18156 15978 18184 18226
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 18248 17649 18276 18022
rect 18340 17921 18368 19246
rect 18432 19145 18460 19926
rect 18418 19136 18474 19145
rect 18418 19071 18474 19080
rect 18326 17912 18382 17921
rect 18326 17847 18382 17856
rect 18234 17640 18290 17649
rect 18234 17575 18290 17584
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 18156 15706 18184 15914
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17880 13870 17908 14010
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 17866 13560 17922 13569
rect 18248 13530 18276 13670
rect 17866 13495 17922 13504
rect 18236 13524 18288 13530
rect 17498 13223 17554 13232
rect 17776 13252 17828 13258
rect 17512 12306 17540 13223
rect 17776 13194 17828 13200
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17316 12232 17368 12238
rect 17236 12192 17316 12220
rect 17316 12174 17368 12180
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17328 11898 17356 12174
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17420 11082 17448 12174
rect 17512 11898 17540 12242
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17880 11801 17908 13495
rect 18236 13466 18288 13472
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 18064 13161 18092 13330
rect 18236 13252 18288 13258
rect 18236 13194 18288 13200
rect 18050 13152 18106 13161
rect 18050 13087 18106 13096
rect 18064 12442 18092 13087
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18248 11898 18276 13194
rect 18340 12986 18368 13466
rect 18432 13394 18460 19071
rect 18524 17490 18552 21383
rect 18616 20777 18644 24006
rect 18708 23866 18736 24142
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 18708 23254 18736 23802
rect 18696 23248 18748 23254
rect 18696 23190 18748 23196
rect 18708 22778 18736 23190
rect 18696 22772 18748 22778
rect 18696 22714 18748 22720
rect 18602 20768 18658 20777
rect 18602 20703 18658 20712
rect 18694 19000 18750 19009
rect 18694 18935 18750 18944
rect 18708 18902 18736 18935
rect 18696 18896 18748 18902
rect 18696 18838 18748 18844
rect 18708 18222 18736 18838
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18800 17762 18828 24550
rect 19168 24070 19196 25230
rect 19352 24818 19380 25910
rect 19812 25786 19840 27520
rect 19444 25758 19840 25786
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19444 24721 19472 25758
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19524 25152 19576 25158
rect 19524 25094 19576 25100
rect 19430 24712 19486 24721
rect 19430 24647 19486 24656
rect 19536 24410 19564 25094
rect 20166 24984 20222 24993
rect 20166 24919 20222 24928
rect 20076 24880 20128 24886
rect 20076 24822 20128 24828
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 19524 24404 19576 24410
rect 19524 24346 19576 24352
rect 19260 24313 19288 24346
rect 19246 24304 19302 24313
rect 19246 24239 19302 24248
rect 19340 24268 19392 24274
rect 19340 24210 19392 24216
rect 19248 24132 19300 24138
rect 19248 24074 19300 24080
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18708 17734 18828 17762
rect 18524 17462 18644 17490
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18524 15706 18552 16526
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18616 15586 18644 17462
rect 18524 15558 18644 15586
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18524 13161 18552 15558
rect 18708 15065 18736 17734
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18800 17338 18828 17614
rect 18892 17338 18920 22578
rect 18972 22092 19024 22098
rect 18972 22034 19024 22040
rect 18984 21622 19012 22034
rect 18972 21616 19024 21622
rect 18972 21558 19024 21564
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 19076 20233 19104 21286
rect 19168 21078 19196 24006
rect 19260 23662 19288 24074
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19260 23186 19288 23598
rect 19352 23526 19380 24210
rect 19536 24138 19564 24346
rect 19524 24132 19576 24138
rect 19524 24074 19576 24080
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19248 23180 19300 23186
rect 19248 23122 19300 23128
rect 19248 22636 19300 22642
rect 19352 22624 19380 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19996 22778 20024 24550
rect 20088 24410 20116 24822
rect 20180 24682 20208 24919
rect 20364 24698 20392 27520
rect 20812 25764 20864 25770
rect 20812 25706 20864 25712
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20168 24676 20220 24682
rect 20168 24618 20220 24624
rect 20272 24670 20392 24698
rect 20180 24410 20208 24618
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 20168 24404 20220 24410
rect 20168 24346 20220 24352
rect 20272 23769 20300 24670
rect 20352 24132 20404 24138
rect 20352 24074 20404 24080
rect 20258 23760 20314 23769
rect 20364 23730 20392 24074
rect 20258 23695 20314 23704
rect 20352 23724 20404 23730
rect 20352 23666 20404 23672
rect 20456 23610 20484 24754
rect 20272 23582 20484 23610
rect 20548 23594 20576 24754
rect 20720 24608 20772 24614
rect 20640 24568 20720 24596
rect 20536 23588 20588 23594
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 19300 22596 19380 22624
rect 19248 22578 19300 22584
rect 19996 22574 20024 22714
rect 19984 22568 20036 22574
rect 19522 22536 19578 22545
rect 19984 22510 20036 22516
rect 19522 22471 19578 22480
rect 19338 22400 19394 22409
rect 19338 22335 19394 22344
rect 19352 21690 19380 22335
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19156 21072 19208 21078
rect 19156 21014 19208 21020
rect 19168 20330 19196 21014
rect 19352 20788 19380 21082
rect 19444 20806 19472 21422
rect 19260 20760 19380 20788
rect 19432 20800 19484 20806
rect 19260 20602 19288 20760
rect 19432 20742 19484 20748
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 19062 20224 19118 20233
rect 19062 20159 19118 20168
rect 19338 20088 19394 20097
rect 19338 20023 19394 20032
rect 19352 19854 19380 20023
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18984 18290 19012 19246
rect 19064 19236 19116 19242
rect 19064 19178 19116 19184
rect 19076 18970 19104 19178
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 19156 18828 19208 18834
rect 19156 18770 19208 18776
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 19168 17814 19196 18770
rect 19260 18329 19288 19654
rect 19352 19514 19380 19790
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19352 18902 19380 19450
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19352 18465 19380 18838
rect 19338 18456 19394 18465
rect 19338 18391 19394 18400
rect 19246 18320 19302 18329
rect 19246 18255 19302 18264
rect 19248 18216 19300 18222
rect 19352 18204 19380 18391
rect 19300 18176 19380 18204
rect 19248 18158 19300 18164
rect 19156 17808 19208 17814
rect 19156 17750 19208 17756
rect 19062 17640 19118 17649
rect 19062 17575 19118 17584
rect 19076 17542 19104 17575
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18800 16153 18828 17274
rect 18892 16697 18920 17274
rect 19076 17134 19104 17478
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 18878 16688 18934 16697
rect 18878 16623 18934 16632
rect 18786 16144 18842 16153
rect 18786 16079 18842 16088
rect 18786 15872 18842 15881
rect 18786 15807 18842 15816
rect 18694 15056 18750 15065
rect 18694 14991 18750 15000
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18510 13152 18566 13161
rect 18510 13087 18566 13096
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18524 12238 18552 12650
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 17866 11792 17922 11801
rect 17866 11727 17922 11736
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17130 10976 17186 10985
rect 17130 10911 17186 10920
rect 17144 6905 17172 10911
rect 18616 9489 18644 13738
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18708 13530 18736 13670
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18708 12986 18736 13262
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18696 12640 18748 12646
rect 18694 12608 18696 12617
rect 18748 12608 18750 12617
rect 18694 12543 18750 12552
rect 17958 9480 18014 9489
rect 17958 9415 18014 9424
rect 18602 9480 18658 9489
rect 18602 9415 18658 9424
rect 17972 7721 18000 9415
rect 17958 7712 18014 7721
rect 17958 7647 18014 7656
rect 17130 6896 17186 6905
rect 17130 6831 17186 6840
rect 17314 6896 17370 6905
rect 17314 6831 17370 6840
rect 17328 6361 17356 6831
rect 18800 6361 18828 15807
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18892 15162 18920 15506
rect 18984 15366 19012 17070
rect 19168 16810 19196 17750
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 19260 16810 19288 17070
rect 19076 16794 19196 16810
rect 19251 16794 19288 16810
rect 19064 16788 19196 16794
rect 19116 16782 19196 16788
rect 19248 16788 19300 16794
rect 19064 16730 19116 16736
rect 19248 16730 19300 16736
rect 19154 16688 19210 16697
rect 19260 16674 19288 16730
rect 19154 16623 19210 16632
rect 19251 16646 19288 16674
rect 19062 16552 19118 16561
rect 19168 16522 19196 16623
rect 19251 16572 19279 16646
rect 19251 16544 19288 16572
rect 19062 16487 19118 16496
rect 19156 16516 19208 16522
rect 19076 16153 19104 16487
rect 19260 16504 19288 16544
rect 19340 16516 19392 16522
rect 19260 16476 19340 16504
rect 19156 16458 19208 16464
rect 19340 16458 19392 16464
rect 19062 16144 19118 16153
rect 19062 16079 19118 16088
rect 19246 15736 19302 15745
rect 19302 15706 19380 15722
rect 19302 15700 19392 15706
rect 19302 15694 19340 15700
rect 19246 15671 19302 15680
rect 19340 15642 19392 15648
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 19248 15360 19300 15366
rect 19300 15308 19380 15314
rect 19248 15302 19380 15308
rect 19260 15286 19380 15302
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18970 15056 19026 15065
rect 18970 14991 19026 15000
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18892 12442 18920 12922
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18984 11121 19012 14991
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19260 14618 19288 14826
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19260 14056 19288 14554
rect 19352 14278 19380 15286
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19168 14028 19288 14056
rect 19168 13326 19196 14028
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 19168 12918 19196 13262
rect 19260 12918 19288 13874
rect 19340 13796 19392 13802
rect 19340 13738 19392 13744
rect 19352 13190 19380 13738
rect 19444 13705 19472 20742
rect 19536 20058 19564 22471
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19524 19916 19576 19922
rect 19996 19904 20024 21830
rect 20088 21146 20116 22170
rect 20076 21140 20128 21146
rect 20076 21082 20128 21088
rect 20088 20466 20116 21082
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 20074 20088 20130 20097
rect 20074 20023 20130 20032
rect 19524 19858 19576 19864
rect 19904 19876 20024 19904
rect 19536 18970 19564 19858
rect 19904 19310 19932 19876
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19536 18426 19564 18906
rect 19996 18834 20024 19722
rect 20088 19242 20116 20023
rect 20180 19990 20208 20946
rect 20168 19984 20220 19990
rect 20168 19926 20220 19932
rect 20076 19236 20128 19242
rect 20076 19178 20128 19184
rect 20088 18970 20116 19178
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19536 17066 19564 18226
rect 19996 18154 20024 18770
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19996 17882 20024 18090
rect 19984 17876 20036 17882
rect 20272 17864 20300 23582
rect 20536 23530 20588 23536
rect 20352 23520 20404 23526
rect 20352 23462 20404 23468
rect 20364 19394 20392 23462
rect 20548 23322 20576 23530
rect 20536 23316 20588 23322
rect 20536 23258 20588 23264
rect 20548 22166 20576 23258
rect 20640 22778 20668 24568
rect 20720 24550 20772 24556
rect 20824 24206 20852 25706
rect 20916 25362 20944 27520
rect 20904 25356 20956 25362
rect 20904 25298 20956 25304
rect 21180 25356 21232 25362
rect 21180 25298 21232 25304
rect 21192 24614 21220 25298
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21180 24608 21232 24614
rect 21180 24550 21232 24556
rect 21088 24268 21140 24274
rect 21088 24210 21140 24216
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 20720 24064 20772 24070
rect 20720 24006 20772 24012
rect 20628 22772 20680 22778
rect 20628 22714 20680 22720
rect 20536 22160 20588 22166
rect 20536 22102 20588 22108
rect 20536 21956 20588 21962
rect 20536 21898 20588 21904
rect 20548 21554 20576 21898
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20456 19718 20484 20198
rect 20548 19854 20576 21490
rect 20732 21418 20760 24006
rect 20824 23526 20852 24142
rect 20812 23520 20864 23526
rect 20812 23462 20864 23468
rect 20994 23352 21050 23361
rect 20994 23287 21050 23296
rect 20904 22500 20956 22506
rect 20904 22442 20956 22448
rect 20916 22234 20944 22442
rect 20904 22228 20956 22234
rect 20904 22170 20956 22176
rect 20720 21412 20772 21418
rect 20720 21354 20772 21360
rect 20732 21146 20760 21354
rect 20720 21140 20772 21146
rect 20720 21082 20772 21088
rect 20812 21072 20864 21078
rect 20812 21014 20864 21020
rect 20628 20392 20680 20398
rect 20824 20346 20852 21014
rect 20680 20340 20852 20346
rect 20628 20334 20852 20340
rect 20640 20318 20852 20334
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20628 19508 20680 19514
rect 20824 19496 20852 20318
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20680 19468 20852 19496
rect 20628 19450 20680 19456
rect 20364 19366 20852 19394
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20364 18426 20392 18566
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 20272 17836 20484 17864
rect 19984 17818 20036 17824
rect 19524 17060 19576 17066
rect 19524 17002 19576 17008
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19996 16794 20024 17818
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19720 16250 19748 16526
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19996 16182 20024 16730
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19996 15706 20024 16118
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 20272 15502 20300 15846
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20272 15162 20300 15438
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19616 14544 19668 14550
rect 19616 14486 19668 14492
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19430 13696 19486 13705
rect 19430 13631 19486 13640
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 19260 12730 19288 12854
rect 19168 12702 19288 12730
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 18970 11112 19026 11121
rect 18970 11047 19026 11056
rect 19076 7313 19104 12582
rect 19168 12306 19196 12702
rect 19352 12374 19380 13126
rect 19536 12442 19564 14214
rect 19628 13938 19656 14486
rect 19996 14414 20024 14826
rect 20180 14414 20208 14894
rect 20272 14550 20300 15098
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20260 14544 20312 14550
rect 20260 14486 20312 14492
rect 19984 14408 20036 14414
rect 19982 14376 19984 14385
rect 20168 14408 20220 14414
rect 20036 14376 20038 14385
rect 20168 14350 20220 14356
rect 20258 14376 20314 14385
rect 19982 14311 20038 14320
rect 20258 14311 20314 14320
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 20272 13870 20300 14311
rect 20364 14074 20392 14758
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20456 13705 20484 17836
rect 20548 15570 20576 19246
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20732 18170 20760 19110
rect 20640 18142 20760 18170
rect 20640 17524 20668 18142
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20732 17814 20760 18022
rect 20720 17808 20772 17814
rect 20720 17750 20772 17756
rect 20732 17649 20760 17750
rect 20718 17640 20774 17649
rect 20718 17575 20774 17584
rect 20640 17496 20760 17524
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20640 16454 20668 16594
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20548 14958 20576 15506
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20442 13696 20498 13705
rect 19622 13628 19918 13648
rect 20442 13631 20498 13640
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 20548 13394 20576 14418
rect 20640 13530 20668 16390
rect 20732 15745 20760 17496
rect 20718 15736 20774 15745
rect 20824 15706 20852 19366
rect 20916 18970 20944 19790
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20902 18728 20958 18737
rect 20902 18663 20958 18672
rect 20916 17882 20944 18663
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20718 15671 20774 15680
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20720 15632 20772 15638
rect 20720 15574 20772 15580
rect 20732 15450 20760 15574
rect 20916 15450 20944 15846
rect 20732 15422 20944 15450
rect 20732 15366 20760 15422
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 19892 13252 19944 13258
rect 19892 13194 19944 13200
rect 19904 12986 19932 13194
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 20626 12608 20682 12617
rect 19622 12540 19918 12560
rect 20626 12543 20682 12552
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 19248 12232 19300 12238
rect 19800 12232 19852 12238
rect 19248 12174 19300 12180
rect 19798 12200 19800 12209
rect 19852 12200 19854 12209
rect 19260 7993 19288 12174
rect 19798 12135 19854 12144
rect 20640 12073 20668 12543
rect 20626 12064 20682 12073
rect 20626 11999 20682 12008
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19352 8945 19380 9386
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19338 8936 19394 8945
rect 19338 8871 19394 8880
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19246 7984 19302 7993
rect 19246 7919 19302 7928
rect 20732 7449 20760 15302
rect 20824 15026 20852 15302
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20812 14884 20864 14890
rect 20812 14826 20864 14832
rect 20824 13297 20852 14826
rect 20916 14618 20944 14962
rect 21008 14618 21036 23287
rect 21100 22982 21128 24210
rect 21270 23624 21326 23633
rect 21270 23559 21326 23568
rect 21088 22976 21140 22982
rect 21088 22918 21140 22924
rect 21100 22817 21128 22918
rect 21086 22808 21142 22817
rect 21086 22743 21142 22752
rect 21100 22574 21128 22743
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 21178 22400 21234 22409
rect 21178 22335 21234 22344
rect 21192 21690 21220 22335
rect 21284 22234 21312 23559
rect 21272 22228 21324 22234
rect 21272 22170 21324 22176
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 21284 21146 21312 22170
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21376 21350 21404 21966
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21362 20768 21418 20777
rect 21362 20703 21418 20712
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 21178 20224 21234 20233
rect 21100 20058 21128 20198
rect 21178 20159 21234 20168
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 21100 19378 21128 19994
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21086 19272 21142 19281
rect 21086 19207 21142 19216
rect 21100 18970 21128 19207
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 21086 18592 21142 18601
rect 21086 18527 21142 18536
rect 21100 18358 21128 18527
rect 21088 18352 21140 18358
rect 21088 18294 21140 18300
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 21100 16114 21128 16526
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 20810 13288 20866 13297
rect 20810 13223 20866 13232
rect 20916 10033 20944 14282
rect 21008 14074 21036 14418
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 21100 12481 21128 15914
rect 21192 12918 21220 20159
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 21284 19514 21312 19858
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21284 16794 21312 19450
rect 21376 19174 21404 20703
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 21376 18601 21404 18702
rect 21362 18592 21418 18601
rect 21362 18527 21418 18536
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21376 17882 21404 18362
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 21468 17762 21496 25230
rect 21560 22098 21588 27520
rect 21640 24132 21692 24138
rect 21640 24074 21692 24080
rect 21652 23186 21680 24074
rect 22112 23746 22140 27520
rect 22192 25424 22244 25430
rect 22192 25366 22244 25372
rect 22020 23718 22140 23746
rect 21916 23656 21968 23662
rect 21916 23598 21968 23604
rect 21732 23520 21784 23526
rect 21732 23462 21784 23468
rect 21744 23254 21772 23462
rect 21732 23248 21784 23254
rect 21732 23190 21784 23196
rect 21640 23180 21692 23186
rect 21640 23122 21692 23128
rect 21652 22166 21680 23122
rect 21744 22778 21772 23190
rect 21822 23080 21878 23089
rect 21822 23015 21878 23024
rect 21732 22772 21784 22778
rect 21732 22714 21784 22720
rect 21836 22710 21864 23015
rect 21824 22704 21876 22710
rect 21824 22646 21876 22652
rect 21732 22568 21784 22574
rect 21732 22510 21784 22516
rect 21640 22160 21692 22166
rect 21640 22102 21692 22108
rect 21548 22092 21600 22098
rect 21548 22034 21600 22040
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 21560 21350 21588 21830
rect 21744 21672 21772 22510
rect 21824 22092 21876 22098
rect 21824 22034 21876 22040
rect 21652 21644 21772 21672
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21560 20369 21588 21286
rect 21546 20360 21602 20369
rect 21546 20295 21602 20304
rect 21548 18896 21600 18902
rect 21548 18838 21600 18844
rect 21560 18358 21588 18838
rect 21548 18352 21600 18358
rect 21548 18294 21600 18300
rect 21376 17734 21496 17762
rect 21548 17740 21600 17746
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 21284 16250 21312 16730
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21284 12986 21312 16186
rect 21376 14482 21404 17734
rect 21548 17682 21600 17688
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21468 17066 21496 17614
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 21560 16697 21588 17682
rect 21546 16688 21602 16697
rect 21546 16623 21602 16632
rect 21456 15632 21508 15638
rect 21456 15574 21508 15580
rect 21468 14890 21496 15574
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21560 14618 21588 16623
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21652 14346 21680 21644
rect 21732 21548 21784 21554
rect 21732 21490 21784 21496
rect 21744 21146 21772 21490
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21836 20890 21864 22034
rect 21928 21962 21956 23598
rect 22020 23361 22048 23718
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 22006 23352 22062 23361
rect 22006 23287 22062 23296
rect 22006 23080 22062 23089
rect 22006 23015 22062 23024
rect 22020 22778 22048 23015
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 22006 22672 22062 22681
rect 22006 22607 22062 22616
rect 21916 21956 21968 21962
rect 21916 21898 21968 21904
rect 22020 21146 22048 22607
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 21744 20862 21864 20890
rect 21744 19496 21772 20862
rect 21824 20800 21876 20806
rect 21822 20768 21824 20777
rect 21876 20768 21878 20777
rect 21822 20703 21878 20712
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21836 20058 21864 20198
rect 21824 20052 21876 20058
rect 21824 19994 21876 20000
rect 22020 19990 22048 21082
rect 22008 19984 22060 19990
rect 22006 19952 22008 19961
rect 22060 19952 22062 19961
rect 22006 19887 22062 19896
rect 21916 19712 21968 19718
rect 21916 19654 21968 19660
rect 21744 19468 21864 19496
rect 21730 19408 21786 19417
rect 21730 19343 21786 19352
rect 21744 19310 21772 19343
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21744 18970 21772 19246
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21744 17134 21772 18702
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21744 16658 21772 17070
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21730 16280 21786 16289
rect 21730 16215 21786 16224
rect 21640 14340 21692 14346
rect 21640 14282 21692 14288
rect 21454 14240 21510 14249
rect 21454 14175 21510 14184
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21180 12912 21232 12918
rect 21180 12854 21232 12860
rect 21284 12782 21312 12922
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 21086 12472 21142 12481
rect 21086 12407 21142 12416
rect 20902 10024 20958 10033
rect 20902 9959 20958 9968
rect 20994 9072 21050 9081
rect 20994 9007 21050 9016
rect 20718 7440 20774 7449
rect 20718 7375 20774 7384
rect 19062 7304 19118 7313
rect 19062 7239 19118 7248
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 17314 6352 17370 6361
rect 17314 6287 17370 6296
rect 18786 6352 18842 6361
rect 18786 6287 18842 6296
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 21008 5137 21036 9007
rect 21284 7857 21312 12718
rect 21468 11762 21496 14175
rect 21638 13560 21694 13569
rect 21638 13495 21640 13504
rect 21692 13495 21694 13504
rect 21640 13466 21692 13472
rect 21744 12442 21772 16215
rect 21836 16017 21864 19468
rect 21928 19378 21956 19654
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 21928 17814 21956 18226
rect 21916 17808 21968 17814
rect 21916 17750 21968 17756
rect 22008 17604 22060 17610
rect 22008 17546 22060 17552
rect 21916 17060 21968 17066
rect 21916 17002 21968 17008
rect 21928 16794 21956 17002
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 22020 16674 22048 17546
rect 21928 16646 22048 16674
rect 21822 16008 21878 16017
rect 21822 15943 21878 15952
rect 21928 14958 21956 16646
rect 22008 16584 22060 16590
rect 22008 16526 22060 16532
rect 22020 15162 22048 16526
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21836 14346 21864 14758
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 21836 14074 21864 14282
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21928 14006 21956 14894
rect 22006 14784 22062 14793
rect 22006 14719 22062 14728
rect 22020 14618 22048 14719
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 21916 14000 21968 14006
rect 21916 13942 21968 13948
rect 22020 13870 22048 14554
rect 22112 14074 22140 23530
rect 22204 22574 22232 25366
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 22480 24954 22508 25298
rect 22468 24948 22520 24954
rect 22468 24890 22520 24896
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22296 23526 22324 24142
rect 22376 24132 22428 24138
rect 22376 24074 22428 24080
rect 22388 23866 22416 24074
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 22192 22568 22244 22574
rect 22192 22510 22244 22516
rect 22204 22234 22232 22510
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22204 21690 22232 21966
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 22204 20262 22232 20878
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22296 18902 22324 23462
rect 22388 20262 22416 23802
rect 22664 23662 22692 27520
rect 22744 26172 22796 26178
rect 22744 26114 22796 26120
rect 22756 25430 22784 26114
rect 22744 25424 22796 25430
rect 22744 25366 22796 25372
rect 23112 24676 23164 24682
rect 23112 24618 23164 24624
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22848 23594 22876 24210
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 22468 23588 22520 23594
rect 22468 23530 22520 23536
rect 22836 23588 22888 23594
rect 22836 23530 22888 23536
rect 22480 21554 22508 23530
rect 22560 23520 22612 23526
rect 22560 23462 22612 23468
rect 22572 22778 22600 23462
rect 23032 23322 23060 24142
rect 23020 23316 23072 23322
rect 23020 23258 23072 23264
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 23032 22658 23060 23258
rect 22940 22642 23060 22658
rect 22928 22636 23060 22642
rect 22980 22630 23060 22636
rect 22928 22578 22980 22584
rect 22560 22568 22612 22574
rect 22558 22536 22560 22545
rect 22612 22536 22614 22545
rect 22558 22471 22614 22480
rect 22652 22432 22704 22438
rect 22652 22374 22704 22380
rect 22558 22128 22614 22137
rect 22558 22063 22614 22072
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 22466 21448 22522 21457
rect 22466 21383 22522 21392
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22388 19174 22416 19858
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 22192 18692 22244 18698
rect 22192 18634 22244 18640
rect 22204 18154 22232 18634
rect 22282 18320 22338 18329
rect 22282 18255 22338 18264
rect 22296 18222 22324 18255
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 22296 17882 22324 18158
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 22204 16250 22232 17614
rect 22388 17116 22416 19110
rect 22296 17088 22416 17116
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22204 15094 22232 15982
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 22192 14884 22244 14890
rect 22192 14826 22244 14832
rect 22204 14657 22232 14826
rect 22190 14648 22246 14657
rect 22190 14583 22246 14592
rect 22296 14362 22324 17088
rect 22480 16969 22508 21383
rect 22466 16960 22522 16969
rect 22466 16895 22522 16904
rect 22572 16776 22600 22063
rect 22664 20505 22692 22374
rect 22940 22166 22968 22578
rect 22928 22160 22980 22166
rect 22928 22102 22980 22108
rect 22744 22092 22796 22098
rect 22744 22034 22796 22040
rect 22756 21486 22784 22034
rect 22940 21690 22968 22102
rect 22928 21684 22980 21690
rect 22928 21626 22980 21632
rect 22836 21548 22888 21554
rect 22836 21490 22888 21496
rect 22744 21480 22796 21486
rect 22744 21422 22796 21428
rect 22756 21146 22784 21422
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 22650 20496 22706 20505
rect 22650 20431 22706 20440
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22664 20097 22692 20198
rect 22650 20088 22706 20097
rect 22650 20023 22706 20032
rect 22756 19922 22784 21082
rect 22744 19916 22796 19922
rect 22744 19858 22796 19864
rect 22650 19816 22706 19825
rect 22848 19802 22876 21490
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 23032 20262 23060 20878
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 23032 20058 23060 20198
rect 23020 20052 23072 20058
rect 23020 19994 23072 20000
rect 22928 19916 22980 19922
rect 22928 19858 22980 19864
rect 22706 19774 22876 19802
rect 22650 19751 22706 19760
rect 22664 17134 22692 19751
rect 22940 19514 22968 19858
rect 23018 19680 23074 19689
rect 23018 19615 23074 19624
rect 22928 19508 22980 19514
rect 22928 19450 22980 19456
rect 22940 19281 22968 19450
rect 22926 19272 22982 19281
rect 22926 19207 22982 19216
rect 23032 18834 23060 19615
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 22928 18624 22980 18630
rect 22928 18566 22980 18572
rect 22834 18456 22890 18465
rect 22834 18391 22890 18400
rect 22742 17912 22798 17921
rect 22742 17847 22798 17856
rect 22652 17128 22704 17134
rect 22652 17070 22704 17076
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22480 16748 22600 16776
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 22388 15570 22416 16594
rect 22480 16590 22508 16748
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22480 16153 22508 16390
rect 22466 16144 22522 16153
rect 22466 16079 22522 16088
rect 22560 16108 22612 16114
rect 22560 16050 22612 16056
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22376 15564 22428 15570
rect 22376 15506 22428 15512
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22388 14482 22416 15098
rect 22480 14618 22508 15846
rect 22572 15706 22600 16050
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22664 15638 22692 16934
rect 22756 16114 22784 17847
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 22652 15632 22704 15638
rect 22652 15574 22704 15580
rect 22664 15162 22692 15574
rect 22744 15360 22796 15366
rect 22744 15302 22796 15308
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22560 15088 22612 15094
rect 22560 15030 22612 15036
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 22296 14334 22508 14362
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 22008 13864 22060 13870
rect 21822 13832 21878 13841
rect 22008 13806 22060 13812
rect 21822 13767 21878 13776
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21836 12322 21864 13767
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21928 12782 21956 13330
rect 21916 12776 21968 12782
rect 21914 12744 21916 12753
rect 21968 12744 21970 12753
rect 21914 12679 21970 12688
rect 21652 12306 21864 12322
rect 21640 12300 21864 12306
rect 21692 12294 21864 12300
rect 21640 12242 21692 12248
rect 21652 11898 21680 12242
rect 22296 11898 22324 14214
rect 22374 13560 22430 13569
rect 22374 13495 22430 13504
rect 22388 13297 22416 13495
rect 22374 13288 22430 13297
rect 22374 13223 22430 13232
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22282 11792 22338 11801
rect 21456 11756 21508 11762
rect 22282 11727 22284 11736
rect 21456 11698 21508 11704
rect 22336 11727 22338 11736
rect 22284 11698 22336 11704
rect 22374 11656 22430 11665
rect 22374 11591 22430 11600
rect 22388 11218 22416 11591
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 22388 10810 22416 11154
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22480 10169 22508 14334
rect 22572 14278 22600 15030
rect 22664 14822 22692 15098
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22650 14648 22706 14657
rect 22650 14583 22706 14592
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22558 13560 22614 13569
rect 22558 13495 22614 13504
rect 22572 13394 22600 13495
rect 22664 13394 22692 14583
rect 22560 13388 22612 13394
rect 22560 13330 22612 13336
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22572 12918 22600 13330
rect 22650 13016 22706 13025
rect 22650 12951 22652 12960
rect 22704 12951 22706 12960
rect 22652 12922 22704 12928
rect 22560 12912 22612 12918
rect 22560 12854 22612 12860
rect 22756 11354 22784 15302
rect 22848 12986 22876 18391
rect 22940 18057 22968 18566
rect 23032 18086 23060 18770
rect 23020 18080 23072 18086
rect 22926 18048 22982 18057
rect 23020 18022 23072 18028
rect 22926 17983 22982 17992
rect 22928 17672 22980 17678
rect 22926 17640 22928 17649
rect 23020 17672 23072 17678
rect 22980 17640 22982 17649
rect 23020 17614 23072 17620
rect 22926 17575 22982 17584
rect 22926 17368 22982 17377
rect 22926 17303 22982 17312
rect 22940 17270 22968 17303
rect 22928 17264 22980 17270
rect 22928 17206 22980 17212
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22940 16153 22968 17070
rect 23032 16794 23060 17614
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 23020 16652 23072 16658
rect 23020 16594 23072 16600
rect 23032 16182 23060 16594
rect 23020 16176 23072 16182
rect 22926 16144 22982 16153
rect 23020 16118 23072 16124
rect 22926 16079 22982 16088
rect 23124 15994 23152 24618
rect 22940 15966 23152 15994
rect 22940 14793 22968 15966
rect 23112 15904 23164 15910
rect 23032 15852 23112 15858
rect 23032 15846 23164 15852
rect 23032 15830 23152 15846
rect 22926 14784 22982 14793
rect 22926 14719 22982 14728
rect 22928 14612 22980 14618
rect 22928 14554 22980 14560
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22848 12782 22876 12922
rect 22836 12776 22888 12782
rect 22836 12718 22888 12724
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 22466 10160 22522 10169
rect 22466 10095 22522 10104
rect 22940 9353 22968 14554
rect 23032 12306 23060 15830
rect 23110 15736 23166 15745
rect 23110 15671 23166 15680
rect 23124 14618 23152 15671
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23124 14074 23152 14350
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23216 13530 23244 27520
rect 23768 24857 23796 27520
rect 24124 25356 24176 25362
rect 24124 25298 24176 25304
rect 24136 24954 24164 25298
rect 24320 25242 24348 27520
rect 24674 26480 24730 26489
rect 24674 26415 24730 26424
rect 24584 26036 24636 26042
rect 24584 25978 24636 25984
rect 24596 25362 24624 25978
rect 24584 25356 24636 25362
rect 24584 25298 24636 25304
rect 24228 25214 24348 25242
rect 24124 24948 24176 24954
rect 24124 24890 24176 24896
rect 24228 24857 24256 25214
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 23754 24848 23810 24857
rect 23754 24783 23810 24792
rect 24214 24848 24270 24857
rect 24214 24783 24270 24792
rect 24032 24744 24084 24750
rect 24032 24686 24084 24692
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23400 23882 23428 24550
rect 23938 24304 23994 24313
rect 23938 24239 23940 24248
rect 23992 24239 23994 24248
rect 23940 24210 23992 24216
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23492 24041 23520 24142
rect 23572 24064 23624 24070
rect 23478 24032 23534 24041
rect 23572 24006 23624 24012
rect 23478 23967 23534 23976
rect 23400 23854 23520 23882
rect 23388 23520 23440 23526
rect 23388 23462 23440 23468
rect 23400 22930 23428 23462
rect 23492 23050 23520 23854
rect 23584 23322 23612 24006
rect 24044 23866 24072 24686
rect 24688 24614 24716 26415
rect 24766 25936 24822 25945
rect 24766 25871 24822 25880
rect 24780 25498 24808 25871
rect 24768 25492 24820 25498
rect 24768 25434 24820 25440
rect 24766 25256 24822 25265
rect 24766 25191 24822 25200
rect 24780 24886 24808 25191
rect 24768 24880 24820 24886
rect 24768 24822 24820 24828
rect 24872 24818 24900 27520
rect 25044 25220 25096 25226
rect 25044 25162 25096 25168
rect 24860 24812 24912 24818
rect 24860 24754 24912 24760
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24674 24032 24730 24041
rect 24032 23860 24084 23866
rect 24032 23802 24084 23808
rect 24136 23526 24164 24006
rect 24289 23964 24585 23984
rect 24674 23967 24730 23976
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24032 23520 24084 23526
rect 24032 23462 24084 23468
rect 24124 23520 24176 23526
rect 24124 23462 24176 23468
rect 23572 23316 23624 23322
rect 23572 23258 23624 23264
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23860 23089 23888 23122
rect 23940 23112 23992 23118
rect 23846 23080 23902 23089
rect 23480 23044 23532 23050
rect 23940 23054 23992 23060
rect 23846 23015 23902 23024
rect 23480 22986 23532 22992
rect 23400 22902 23520 22930
rect 23492 22080 23520 22902
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23400 22052 23520 22080
rect 23400 20398 23428 22052
rect 23676 21978 23704 22374
rect 23860 22234 23888 23015
rect 23952 22506 23980 23054
rect 23940 22500 23992 22506
rect 23940 22442 23992 22448
rect 23952 22234 23980 22442
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 23940 22228 23992 22234
rect 23940 22170 23992 22176
rect 23656 21950 23704 21978
rect 23656 21876 23684 21950
rect 23848 21888 23900 21894
rect 23656 21848 23796 21876
rect 23768 20398 23796 21848
rect 23848 21830 23900 21836
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23664 20392 23716 20398
rect 23664 20334 23716 20340
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 23584 19258 23612 20198
rect 23676 19786 23704 20334
rect 23768 20058 23796 20334
rect 23756 20052 23808 20058
rect 23756 19994 23808 20000
rect 23664 19780 23716 19786
rect 23664 19722 23716 19728
rect 23400 19230 23612 19258
rect 23296 18964 23348 18970
rect 23296 18906 23348 18912
rect 23308 18465 23336 18906
rect 23294 18456 23350 18465
rect 23294 18391 23296 18400
rect 23348 18391 23350 18400
rect 23296 18362 23348 18368
rect 23296 18080 23348 18086
rect 23296 18022 23348 18028
rect 23308 15745 23336 18022
rect 23400 16810 23428 19230
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23492 18766 23520 19110
rect 23480 18760 23532 18766
rect 23860 18714 23888 21830
rect 23952 21486 23980 22170
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 23952 20262 23980 21082
rect 23940 20256 23992 20262
rect 23940 20198 23992 20204
rect 23480 18702 23532 18708
rect 23492 18426 23520 18702
rect 23572 18692 23624 18698
rect 23572 18634 23624 18640
rect 23676 18686 23888 18714
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23584 17785 23612 18634
rect 23570 17776 23626 17785
rect 23570 17711 23626 17720
rect 23676 17524 23704 18686
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23754 18320 23810 18329
rect 23754 18255 23810 18264
rect 23768 17921 23796 18255
rect 23860 18154 23888 18566
rect 23848 18148 23900 18154
rect 23848 18090 23900 18096
rect 23754 17912 23810 17921
rect 23754 17847 23810 17856
rect 23756 17808 23808 17814
rect 23756 17750 23808 17756
rect 23584 17496 23704 17524
rect 23400 16782 23520 16810
rect 23386 16688 23442 16697
rect 23386 16623 23442 16632
rect 23294 15736 23350 15745
rect 23294 15671 23350 15680
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23308 14618 23336 15506
rect 23400 15201 23428 16623
rect 23386 15192 23442 15201
rect 23386 15127 23442 15136
rect 23492 15076 23520 16782
rect 23400 15048 23520 15076
rect 23400 14770 23428 15048
rect 23478 14920 23534 14929
rect 23478 14855 23480 14864
rect 23532 14855 23534 14864
rect 23480 14826 23532 14832
rect 23400 14742 23520 14770
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 23308 13530 23336 14554
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23400 13870 23428 14418
rect 23492 14074 23520 14742
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23388 13864 23440 13870
rect 23440 13824 23520 13852
rect 23388 13806 23440 13812
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 23204 13388 23256 13394
rect 23204 13330 23256 13336
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23124 12374 23152 12718
rect 23216 12442 23244 13330
rect 23386 12472 23442 12481
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 23296 12436 23348 12442
rect 23492 12442 23520 13824
rect 23386 12407 23442 12416
rect 23480 12436 23532 12442
rect 23296 12378 23348 12384
rect 23112 12368 23164 12374
rect 23112 12310 23164 12316
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23032 11937 23060 12242
rect 23018 11928 23074 11937
rect 23018 11863 23020 11872
rect 23072 11863 23074 11872
rect 23020 11834 23072 11840
rect 23032 11803 23060 11834
rect 23308 10690 23336 12378
rect 23400 11778 23428 12407
rect 23480 12378 23532 12384
rect 23584 11880 23612 17496
rect 23662 17368 23718 17377
rect 23662 17303 23664 17312
rect 23716 17303 23718 17312
rect 23664 17274 23716 17280
rect 23662 16824 23718 16833
rect 23662 16759 23718 16768
rect 23676 15366 23704 16759
rect 23768 16250 23796 17750
rect 23860 17678 23888 18090
rect 23848 17672 23900 17678
rect 24044 17626 24072 23462
rect 24136 20890 24164 23462
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24398 22672 24454 22681
rect 24308 22636 24360 22642
rect 24398 22607 24454 22616
rect 24308 22578 24360 22584
rect 24320 22098 24348 22578
rect 24308 22092 24360 22098
rect 24308 22034 24360 22040
rect 24412 22030 24440 22607
rect 24400 22024 24452 22030
rect 24400 21966 24452 21972
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21593 24716 23967
rect 24872 23322 24900 24210
rect 24952 23520 25004 23526
rect 24952 23462 25004 23468
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24964 22438 24992 23462
rect 24952 22432 25004 22438
rect 24952 22374 25004 22380
rect 24766 22264 24822 22273
rect 25056 22250 25084 25162
rect 25228 23792 25280 23798
rect 25228 23734 25280 23740
rect 25240 22624 25268 23734
rect 25318 23216 25374 23225
rect 25318 23151 25320 23160
rect 25372 23151 25374 23160
rect 25320 23122 25372 23128
rect 25332 22778 25360 23122
rect 25320 22772 25372 22778
rect 25320 22714 25372 22720
rect 25240 22596 25360 22624
rect 25228 22500 25280 22506
rect 25228 22442 25280 22448
rect 25136 22432 25188 22438
rect 25134 22400 25136 22409
rect 25188 22400 25190 22409
rect 25134 22335 25190 22344
rect 25056 22222 25176 22250
rect 24766 22199 24822 22208
rect 24674 21584 24730 21593
rect 24674 21519 24730 21528
rect 24780 21434 24808 22199
rect 24860 21956 24912 21962
rect 24860 21898 24912 21904
rect 24688 21406 24808 21434
rect 24872 21418 24900 21898
rect 24952 21888 25004 21894
rect 24952 21830 25004 21836
rect 24860 21412 24912 21418
rect 24136 20862 24256 20890
rect 24122 20768 24178 20777
rect 24122 20703 24178 20712
rect 24136 20466 24164 20703
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 24122 19816 24178 19825
rect 24122 19751 24178 19760
rect 23848 17614 23900 17620
rect 23952 17598 24072 17626
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23860 16998 23888 17478
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 23860 16096 23888 16458
rect 23768 16068 23888 16096
rect 23768 15502 23796 16068
rect 23846 16008 23902 16017
rect 23846 15943 23902 15952
rect 23756 15496 23808 15502
rect 23756 15438 23808 15444
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23754 15328 23810 15337
rect 23754 15263 23810 15272
rect 23664 14952 23716 14958
rect 23664 14894 23716 14900
rect 23676 14278 23704 14894
rect 23664 14272 23716 14278
rect 23662 14240 23664 14249
rect 23716 14240 23718 14249
rect 23662 14175 23718 14184
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23676 13530 23704 13806
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23676 12782 23704 13466
rect 23664 12776 23716 12782
rect 23768 12753 23796 15263
rect 23860 14362 23888 15943
rect 23952 15162 23980 17598
rect 24032 17536 24084 17542
rect 24032 17478 24084 17484
rect 24044 17241 24072 17478
rect 24030 17232 24086 17241
rect 24030 17167 24086 17176
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 24044 14521 24072 16934
rect 24136 16522 24164 19751
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 24228 16266 24256 20862
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24308 20460 24360 20466
rect 24308 20402 24360 20408
rect 24320 20262 24348 20402
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 17864 24716 21406
rect 24860 21354 24912 21360
rect 24872 21298 24900 21354
rect 24964 21350 24992 21830
rect 24780 21270 24900 21298
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 24780 20602 24808 21270
rect 24964 21010 24992 21286
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 24950 20904 25006 20913
rect 24950 20839 25006 20848
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 24766 20360 24822 20369
rect 24822 20318 24900 20346
rect 24766 20295 24822 20304
rect 24872 20058 24900 20318
rect 24860 20052 24912 20058
rect 24860 19994 24912 20000
rect 24768 19984 24820 19990
rect 24768 19926 24820 19932
rect 24780 19310 24808 19926
rect 24768 19304 24820 19310
rect 24768 19246 24820 19252
rect 24780 18834 24808 19246
rect 24964 18902 24992 20839
rect 25044 20800 25096 20806
rect 25044 20742 25096 20748
rect 25056 20262 25084 20742
rect 25148 20466 25176 22222
rect 25240 22001 25268 22442
rect 25226 21992 25282 22001
rect 25226 21927 25282 21936
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 25332 20398 25360 22596
rect 25320 20392 25372 20398
rect 25320 20334 25372 20340
rect 25136 20324 25188 20330
rect 25136 20266 25188 20272
rect 25044 20256 25096 20262
rect 25044 20198 25096 20204
rect 25056 19990 25084 20198
rect 25044 19984 25096 19990
rect 25044 19926 25096 19932
rect 25042 19272 25098 19281
rect 25042 19207 25098 19216
rect 25056 19174 25084 19207
rect 25044 19168 25096 19174
rect 25044 19110 25096 19116
rect 24952 18896 25004 18902
rect 24952 18838 25004 18844
rect 25042 18864 25098 18873
rect 24768 18828 24820 18834
rect 24768 18770 24820 18776
rect 24780 18714 24808 18770
rect 24780 18686 24900 18714
rect 24872 18222 24900 18686
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 24964 17882 24992 18838
rect 25042 18799 25098 18808
rect 25056 18766 25084 18799
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 25056 18290 25084 18702
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 25042 18048 25098 18057
rect 25042 17983 25098 17992
rect 24952 17876 25004 17882
rect 24688 17836 24900 17864
rect 24398 17776 24454 17785
rect 24398 17711 24400 17720
rect 24452 17711 24454 17720
rect 24768 17740 24820 17746
rect 24400 17682 24452 17688
rect 24872 17728 24900 17836
rect 24952 17818 25004 17824
rect 24872 17700 24992 17728
rect 24768 17682 24820 17688
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24306 17232 24362 17241
rect 24688 17202 24716 17614
rect 24780 17513 24808 17682
rect 24858 17640 24914 17649
rect 24858 17575 24914 17584
rect 24766 17504 24822 17513
rect 24766 17439 24822 17448
rect 24766 17368 24822 17377
rect 24766 17303 24822 17312
rect 24306 17167 24362 17176
rect 24676 17196 24728 17202
rect 24320 16833 24348 17167
rect 24676 17138 24728 17144
rect 24676 16992 24728 16998
rect 24674 16960 24676 16969
rect 24728 16960 24730 16969
rect 24674 16895 24730 16904
rect 24306 16824 24362 16833
rect 24306 16759 24362 16768
rect 24674 16824 24730 16833
rect 24674 16759 24730 16768
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24136 16238 24256 16266
rect 24136 15434 24164 16238
rect 24216 16108 24268 16114
rect 24216 16050 24268 16056
rect 24228 15706 24256 16050
rect 24216 15700 24268 15706
rect 24216 15642 24268 15648
rect 24124 15428 24176 15434
rect 24124 15370 24176 15376
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15094 24716 16759
rect 24780 16153 24808 17303
rect 24872 16794 24900 17575
rect 24964 16833 24992 17700
rect 24950 16824 25006 16833
rect 24860 16788 24912 16794
rect 24950 16759 25006 16768
rect 24860 16730 24912 16736
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 24964 16561 24992 16594
rect 24950 16552 25006 16561
rect 24950 16487 25006 16496
rect 24860 16448 24912 16454
rect 24858 16416 24860 16425
rect 24912 16416 24914 16425
rect 24858 16351 24914 16360
rect 24964 16250 24992 16487
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 24766 16144 24822 16153
rect 24766 16079 24822 16088
rect 24768 15904 24820 15910
rect 24820 15852 24992 15858
rect 24768 15846 24992 15852
rect 24780 15830 24992 15846
rect 24860 15496 24912 15502
rect 24766 15464 24822 15473
rect 24860 15438 24912 15444
rect 24766 15399 24822 15408
rect 24780 15162 24808 15399
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24676 15088 24728 15094
rect 24676 15030 24728 15036
rect 24872 14634 24900 15438
rect 24780 14606 24900 14634
rect 24030 14512 24086 14521
rect 24030 14447 24086 14456
rect 24216 14476 24268 14482
rect 24216 14418 24268 14424
rect 23860 14334 23980 14362
rect 23664 12718 23716 12724
rect 23754 12744 23810 12753
rect 23754 12679 23810 12688
rect 23952 12322 23980 14334
rect 24228 13977 24256 14418
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24214 13968 24270 13977
rect 24214 13903 24270 13912
rect 24214 13424 24270 13433
rect 24032 13388 24084 13394
rect 24214 13359 24270 13368
rect 24032 13330 24084 13336
rect 23860 12294 23980 12322
rect 23584 11852 23796 11880
rect 23400 11750 23612 11778
rect 23480 11212 23532 11218
rect 23480 11154 23532 11160
rect 23492 10985 23520 11154
rect 23478 10976 23534 10985
rect 23478 10911 23534 10920
rect 23492 10810 23520 10911
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23308 10662 23520 10690
rect 22926 9344 22982 9353
rect 22926 9279 22982 9288
rect 23492 8945 23520 10662
rect 23584 10577 23612 11750
rect 23662 11248 23718 11257
rect 23662 11183 23718 11192
rect 23570 10568 23626 10577
rect 23570 10503 23626 10512
rect 23478 8936 23534 8945
rect 23478 8871 23534 8880
rect 21270 7848 21326 7857
rect 21270 7783 21326 7792
rect 23676 5817 23704 11183
rect 23768 11082 23796 11852
rect 23860 11762 23888 12294
rect 23940 12232 23992 12238
rect 23940 12174 23992 12180
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23848 11552 23900 11558
rect 23848 11494 23900 11500
rect 23756 11076 23808 11082
rect 23756 11018 23808 11024
rect 23860 9625 23888 11494
rect 23952 10810 23980 12174
rect 24044 12170 24072 13330
rect 24228 13326 24256 13359
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24122 12880 24178 12889
rect 24122 12815 24178 12824
rect 24136 12374 24164 12815
rect 24398 12472 24454 12481
rect 24216 12436 24268 12442
rect 24688 12442 24716 14350
rect 24398 12407 24454 12416
rect 24676 12436 24728 12442
rect 24216 12378 24268 12384
rect 24124 12368 24176 12374
rect 24124 12310 24176 12316
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 24032 12164 24084 12170
rect 24032 12106 24084 12112
rect 24032 11756 24084 11762
rect 24032 11698 24084 11704
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 23938 10160 23994 10169
rect 23938 10095 23994 10104
rect 23846 9616 23902 9625
rect 23846 9551 23902 9560
rect 23662 5808 23718 5817
rect 23662 5743 23718 5752
rect 20994 5128 21050 5137
rect 20994 5063 21050 5072
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 16394 4584 16450 4593
rect 16394 4519 16450 4528
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 19522 4040 19578 4049
rect 19522 3975 19578 3984
rect 14830 3632 14886 3641
rect 14830 3567 14886 3576
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14646 2544 14702 2553
rect 14646 2479 14702 2488
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14186 1456 14242 1465
rect 14186 1391 14242 1400
rect 19536 480 19564 3975
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 23952 3754 23980 10095
rect 24044 9382 24072 11698
rect 24136 11626 24164 12174
rect 24124 11620 24176 11626
rect 24124 11562 24176 11568
rect 24124 11144 24176 11150
rect 24124 11086 24176 11092
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 24136 3913 24164 11086
rect 24228 9654 24256 12378
rect 24412 12238 24440 12407
rect 24676 12378 24728 12384
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 24504 11150 24532 11494
rect 24582 11384 24638 11393
rect 24688 11354 24716 12174
rect 24582 11319 24638 11328
rect 24676 11348 24728 11354
rect 24596 11218 24624 11319
rect 24676 11290 24728 11296
rect 24584 11212 24636 11218
rect 24584 11154 24636 11160
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24398 10704 24454 10713
rect 24398 10639 24400 10648
rect 24452 10639 24454 10648
rect 24400 10610 24452 10616
rect 24780 10266 24808 14606
rect 24858 13968 24914 13977
rect 24858 13903 24914 13912
rect 24872 13530 24900 13903
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24872 11898 24900 12242
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24964 11762 24992 15830
rect 25056 15722 25084 17983
rect 25148 16794 25176 20266
rect 25320 19848 25372 19854
rect 25320 19790 25372 19796
rect 25332 19242 25360 19790
rect 25320 19236 25372 19242
rect 25320 19178 25372 19184
rect 25228 19168 25280 19174
rect 25228 19110 25280 19116
rect 25240 17218 25268 19110
rect 25424 17270 25452 27520
rect 25502 27160 25558 27169
rect 25502 27095 25558 27104
rect 25516 24410 25544 27095
rect 25504 24404 25556 24410
rect 25504 24346 25556 24352
rect 25608 23866 25636 27639
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 25872 25900 25924 25906
rect 25872 25842 25924 25848
rect 25780 24268 25832 24274
rect 25780 24210 25832 24216
rect 25792 23866 25820 24210
rect 25596 23860 25648 23866
rect 25596 23802 25648 23808
rect 25780 23860 25832 23866
rect 25780 23802 25832 23808
rect 25502 23352 25558 23361
rect 25502 23287 25504 23296
rect 25556 23287 25558 23296
rect 25504 23258 25556 23264
rect 25792 22545 25820 23802
rect 25778 22536 25834 22545
rect 25778 22471 25834 22480
rect 25502 21584 25558 21593
rect 25502 21519 25558 21528
rect 25412 17264 25464 17270
rect 25240 17190 25360 17218
rect 25412 17206 25464 17212
rect 25228 17128 25280 17134
rect 25226 17096 25228 17105
rect 25280 17096 25282 17105
rect 25226 17031 25282 17040
rect 25136 16788 25188 16794
rect 25136 16730 25188 16736
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 25056 15706 25176 15722
rect 25044 15700 25176 15706
rect 25096 15694 25176 15700
rect 25044 15642 25096 15648
rect 25044 15564 25096 15570
rect 25044 15506 25096 15512
rect 25056 15473 25084 15506
rect 25042 15464 25098 15473
rect 25042 15399 25098 15408
rect 25148 14618 25176 15694
rect 25240 15609 25268 15982
rect 25226 15600 25282 15609
rect 25226 15535 25282 15544
rect 25332 15502 25360 17190
rect 25412 17060 25464 17066
rect 25412 17002 25464 17008
rect 25320 15496 25372 15502
rect 25320 15438 25372 15444
rect 25332 15162 25360 15438
rect 25320 15156 25372 15162
rect 25320 15098 25372 15104
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 25424 13841 25452 17002
rect 25516 16250 25544 21519
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25700 20806 25728 21286
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 25594 20088 25650 20097
rect 25594 20023 25650 20032
rect 25608 19854 25636 20023
rect 25688 19916 25740 19922
rect 25688 19858 25740 19864
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25608 18902 25636 19790
rect 25700 19174 25728 19858
rect 25780 19236 25832 19242
rect 25780 19178 25832 19184
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25596 18896 25648 18902
rect 25596 18838 25648 18844
rect 25594 18184 25650 18193
rect 25594 18119 25596 18128
rect 25648 18119 25650 18128
rect 25596 18090 25648 18096
rect 25608 17882 25636 18090
rect 25596 17876 25648 17882
rect 25596 17818 25648 17824
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25608 16726 25636 16934
rect 25596 16720 25648 16726
rect 25596 16662 25648 16668
rect 25608 16250 25636 16662
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25596 16244 25648 16250
rect 25596 16186 25648 16192
rect 25410 13832 25466 13841
rect 25410 13767 25466 13776
rect 25044 13728 25096 13734
rect 25044 13670 25096 13676
rect 25056 12782 25084 13670
rect 25320 13388 25372 13394
rect 25320 13330 25372 13336
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 25056 11898 25084 12718
rect 25332 12646 25360 13330
rect 25136 12640 25188 12646
rect 25320 12640 25372 12646
rect 25136 12582 25188 12588
rect 25318 12608 25320 12617
rect 25372 12608 25374 12617
rect 25148 12481 25176 12582
rect 25318 12543 25374 12552
rect 25134 12472 25190 12481
rect 25134 12407 25190 12416
rect 25700 12209 25728 19110
rect 25686 12200 25742 12209
rect 25686 12135 25742 12144
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24872 10810 24900 11154
rect 25792 10810 25820 19178
rect 25884 18698 25912 25842
rect 25872 18692 25924 18698
rect 25872 18634 25924 18640
rect 25884 18426 25912 18634
rect 25872 18420 25924 18426
rect 25872 18362 25924 18368
rect 25872 17536 25924 17542
rect 25872 17478 25924 17484
rect 25884 13569 25912 17478
rect 25870 13560 25926 13569
rect 25870 13495 25926 13504
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 24766 10160 24822 10169
rect 24676 10124 24728 10130
rect 24766 10095 24822 10104
rect 24676 10066 24728 10072
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24216 9648 24268 9654
rect 24216 9590 24268 9596
rect 24688 9489 24716 10066
rect 24674 9480 24730 9489
rect 24674 9415 24730 9424
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24122 3904 24178 3913
rect 24122 3839 24178 3848
rect 23952 3726 24164 3754
rect 23478 3632 23534 3641
rect 23478 3567 23534 3576
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 12898 96 12954 105
rect 12898 31 12954 40
rect 13910 0 13966 480
rect 19522 0 19578 480
rect 23492 377 23520 3567
rect 24136 2689 24164 3726
rect 24674 3496 24730 3505
rect 24674 3431 24730 3440
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24122 2680 24178 2689
rect 24122 2615 24178 2624
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 2145 24716 3431
rect 24780 3369 24808 10095
rect 25136 9512 25188 9518
rect 25134 9480 25136 9489
rect 25188 9480 25190 9489
rect 25976 9450 26004 27520
rect 26528 27470 26556 27520
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 26516 27464 26568 27470
rect 26516 27406 26568 27412
rect 26056 24812 26108 24818
rect 26056 24754 26108 24760
rect 26068 13530 26096 24754
rect 26238 24712 26294 24721
rect 26238 24647 26294 24656
rect 26148 22024 26200 22030
rect 26148 21966 26200 21972
rect 26160 17542 26188 21966
rect 26252 20330 26280 24647
rect 26240 20324 26292 20330
rect 26240 20266 26292 20272
rect 26330 19136 26386 19145
rect 26330 19071 26386 19080
rect 26238 17912 26294 17921
rect 26238 17847 26294 17856
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26148 17264 26200 17270
rect 26252 17241 26280 17847
rect 26148 17206 26200 17212
rect 26238 17232 26294 17241
rect 26056 13524 26108 13530
rect 26056 13466 26108 13472
rect 26160 10441 26188 17206
rect 26238 17167 26294 17176
rect 26240 16176 26292 16182
rect 26240 16118 26292 16124
rect 26252 13161 26280 16118
rect 26238 13152 26294 13161
rect 26238 13087 26294 13096
rect 26344 11286 26372 19071
rect 26332 11280 26384 11286
rect 26332 11222 26384 11228
rect 26146 10432 26202 10441
rect 26146 10367 26202 10376
rect 25134 9415 25190 9424
rect 25964 9444 26016 9450
rect 25964 9386 26016 9392
rect 26436 6905 26464 27406
rect 27080 25430 27108 27520
rect 27068 25424 27120 25430
rect 27068 25366 27120 25372
rect 27632 24449 27660 27520
rect 27618 24440 27674 24449
rect 27618 24375 27674 24384
rect 26422 6896 26478 6905
rect 26422 6831 26478 6840
rect 24766 3360 24822 3369
rect 24766 3295 24822 3304
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 24674 2136 24730 2145
rect 24674 2071 24730 2080
rect 25148 480 25176 2246
rect 23478 368 23534 377
rect 23478 303 23534 312
rect 25134 0 25190 480
<< via2 >>
rect 3514 27648 3570 27704
rect 2778 25880 2834 25936
rect 2502 24928 2558 24984
rect 2686 25200 2742 25256
rect 1582 24656 1638 24712
rect 1582 22208 1638 22264
rect 1490 21936 1546 21992
rect 1398 20984 1454 21040
rect 1674 20304 1730 20360
rect 1582 19760 1638 19816
rect 2226 23568 2282 23624
rect 2042 20204 2044 20224
rect 2044 20204 2096 20224
rect 2096 20204 2098 20224
rect 2042 20168 2098 20204
rect 1950 19216 2006 19272
rect 1674 17040 1730 17096
rect 1582 16632 1638 16688
rect 1398 16088 1454 16144
rect 754 15952 810 16008
rect 1858 16632 1914 16688
rect 1674 15136 1730 15192
rect 2594 24384 2650 24440
rect 2410 23296 2466 23352
rect 25594 27648 25650 27704
rect 3054 24112 3110 24168
rect 2502 22208 2558 22264
rect 2410 21664 2466 21720
rect 2778 22752 2834 22808
rect 2778 22228 2834 22264
rect 2778 22208 2780 22228
rect 2780 22208 2832 22228
rect 2832 22208 2834 22228
rect 2686 21528 2742 21584
rect 2594 21392 2650 21448
rect 3238 24268 3294 24304
rect 3238 24248 3240 24268
rect 3240 24248 3292 24268
rect 3292 24248 3294 24268
rect 3330 22616 3386 22672
rect 3238 21936 3294 21992
rect 2502 18128 2558 18184
rect 2318 16224 2374 16280
rect 2962 18264 3018 18320
rect 3146 20848 3202 20904
rect 3238 19896 3294 19952
rect 3790 27104 3846 27160
rect 4066 26424 4122 26480
rect 4158 25744 4214 25800
rect 3606 21256 3662 21312
rect 3606 20460 3662 20496
rect 3606 20440 3608 20460
rect 3608 20440 3660 20460
rect 3660 20440 3662 20460
rect 3422 19760 3478 19816
rect 3790 23976 3846 24032
rect 4066 23432 4122 23488
rect 3882 21936 3938 21992
rect 3698 19352 3754 19408
rect 3606 19080 3662 19136
rect 3422 17584 3478 17640
rect 2778 14592 2834 14648
rect 3330 16768 3386 16824
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 4250 20304 4306 20360
rect 3882 19080 3938 19136
rect 3698 17856 3754 17912
rect 3330 14592 3386 14648
rect 3238 14320 3294 14376
rect 2778 13232 2834 13288
rect 1398 10648 1454 10704
rect 1582 10512 1638 10568
rect 1398 8372 1400 8392
rect 1400 8372 1452 8392
rect 1452 8372 1454 8392
rect 1398 8336 1454 8372
rect 1398 5772 1454 5808
rect 1398 5752 1400 5772
rect 1400 5752 1452 5772
rect 1452 5752 1454 5772
rect 2778 3440 2834 3496
rect 570 2624 626 2680
rect 2870 3304 2926 3360
rect 3514 15408 3570 15464
rect 3422 13640 3478 13696
rect 3422 13096 3478 13152
rect 3882 15444 3884 15464
rect 3884 15444 3936 15464
rect 3936 15444 3938 15464
rect 3882 15408 3938 15444
rect 3790 14864 3846 14920
rect 3882 14728 3938 14784
rect 3514 12688 3570 12744
rect 4250 18536 4306 18592
rect 4066 17992 4122 18048
rect 4342 16904 4398 16960
rect 4066 16088 4122 16144
rect 3882 13232 3938 13288
rect 4158 15852 4160 15872
rect 4160 15852 4212 15872
rect 4212 15852 4214 15872
rect 4158 15816 4214 15852
rect 4250 15544 4306 15600
rect 3422 12144 3478 12200
rect 4618 16224 4674 16280
rect 4526 15000 4582 15056
rect 4434 14592 4490 14648
rect 4066 11872 4122 11928
rect 5170 23568 5226 23624
rect 6090 24520 6146 24576
rect 4894 22344 4950 22400
rect 4710 15680 4766 15736
rect 4710 12844 4766 12880
rect 4710 12824 4712 12844
rect 4712 12824 4764 12844
rect 4764 12824 4766 12844
rect 4710 12280 4766 12336
rect 4618 11464 4674 11520
rect 3882 11056 3938 11112
rect 3882 5072 3938 5128
rect 3514 2080 3570 2136
rect 4066 11192 4122 11248
rect 4066 9560 4122 9616
rect 4066 8744 4122 8800
rect 4066 7792 4122 7848
rect 4066 6976 4122 7032
rect 4066 5208 4122 5264
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5262 21664 5318 21720
rect 5446 22208 5502 22264
rect 6090 21956 6146 21992
rect 6090 21936 6092 21956
rect 6092 21936 6144 21956
rect 6144 21936 6146 21956
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 6918 24384 6974 24440
rect 6458 23840 6514 23896
rect 7102 23296 7158 23352
rect 7286 22500 7342 22536
rect 7286 22480 7288 22500
rect 7288 22480 7340 22500
rect 7340 22480 7342 22500
rect 7194 22380 7196 22400
rect 7196 22380 7248 22400
rect 7248 22380 7250 22400
rect 7194 22344 7250 22380
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5998 20596 6054 20632
rect 5998 20576 6000 20596
rect 6000 20576 6052 20596
rect 6052 20576 6054 20596
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5998 19216 6054 19272
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 6090 18164 6092 18184
rect 6092 18164 6144 18184
rect 6144 18164 6146 18184
rect 6090 18128 6146 18164
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 6090 17040 6146 17096
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5170 15156 5226 15192
rect 5170 15136 5172 15156
rect 5172 15136 5224 15156
rect 5224 15136 5226 15156
rect 5262 14728 5318 14784
rect 5354 14592 5410 14648
rect 5170 14320 5226 14376
rect 5538 15428 5594 15464
rect 5538 15408 5540 15428
rect 5540 15408 5592 15428
rect 5592 15408 5594 15428
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5630 14764 5632 14784
rect 5632 14764 5684 14784
rect 5684 14764 5686 14784
rect 5630 14728 5686 14764
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5170 12824 5226 12880
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 7102 20984 7158 21040
rect 6642 20712 6698 20768
rect 6642 20168 6698 20224
rect 6274 16496 6330 16552
rect 7746 23296 7802 23352
rect 7746 21120 7802 21176
rect 7562 20440 7618 20496
rect 7194 19896 7250 19952
rect 6918 19780 6974 19816
rect 6918 19760 6920 19780
rect 6920 19760 6972 19780
rect 6972 19760 6974 19780
rect 7562 19352 7618 19408
rect 6642 17312 6698 17368
rect 6826 18264 6882 18320
rect 7102 17992 7158 18048
rect 7286 18672 7342 18728
rect 6918 17176 6974 17232
rect 8298 24248 8354 24304
rect 8298 23860 8354 23896
rect 8298 23840 8300 23860
rect 8300 23840 8352 23860
rect 8352 23840 8354 23860
rect 8574 23160 8630 23216
rect 8114 21936 8170 21992
rect 8022 21256 8078 21312
rect 8390 22208 8446 22264
rect 8390 21392 8446 21448
rect 8942 24112 8998 24168
rect 8850 23704 8906 23760
rect 9126 22888 9182 22944
rect 8758 21936 8814 21992
rect 8390 20848 8446 20904
rect 8574 19352 8630 19408
rect 6458 16768 6514 16824
rect 6366 16088 6422 16144
rect 7654 16904 7710 16960
rect 6734 16652 6790 16688
rect 6734 16632 6736 16652
rect 6736 16632 6788 16652
rect 6788 16632 6790 16652
rect 6182 15272 6238 15328
rect 6274 15000 6330 15056
rect 6918 16088 6974 16144
rect 6550 15272 6606 15328
rect 6458 14320 6514 14376
rect 6642 14592 6698 14648
rect 6366 13368 6422 13424
rect 6182 13232 6238 13288
rect 7562 15816 7618 15872
rect 7378 15000 7434 15056
rect 7470 14356 7472 14376
rect 7472 14356 7524 14376
rect 7524 14356 7526 14376
rect 7470 14320 7526 14356
rect 7194 12960 7250 13016
rect 6918 12416 6974 12472
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 7930 18400 7986 18456
rect 8022 18128 8078 18184
rect 8206 16652 8262 16688
rect 8206 16632 8208 16652
rect 8208 16632 8260 16652
rect 8260 16632 8262 16652
rect 8206 16360 8262 16416
rect 8022 15136 8078 15192
rect 8574 18808 8630 18864
rect 8574 16496 8630 16552
rect 8390 15680 8446 15736
rect 7930 12824 7986 12880
rect 8574 13232 8630 13288
rect 8758 17720 8814 17776
rect 8482 12280 8538 12336
rect 7562 11736 7618 11792
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 8298 5616 8354 5672
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5078 5072 5134 5128
rect 4066 4528 4122 4584
rect 3882 1400 3938 1456
rect 3238 856 3294 912
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 8298 3848 8354 3904
rect 9126 21684 9182 21720
rect 9126 21664 9128 21684
rect 9128 21664 9180 21684
rect 9180 21664 9182 21684
rect 9862 24520 9918 24576
rect 9954 24248 10010 24304
rect 9770 23316 9826 23352
rect 9770 23296 9772 23316
rect 9772 23296 9824 23316
rect 9824 23296 9826 23316
rect 9034 20576 9090 20632
rect 9126 15544 9182 15600
rect 9126 13796 9182 13832
rect 9126 13776 9128 13796
rect 9128 13776 9180 13796
rect 9180 13776 9182 13796
rect 9218 11872 9274 11928
rect 9770 21936 9826 21992
rect 9678 21292 9680 21312
rect 9680 21292 9732 21312
rect 9732 21292 9734 21312
rect 9678 21256 9734 21292
rect 9770 21120 9826 21176
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10138 23840 10194 23896
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10966 24556 10968 24576
rect 10968 24556 11020 24576
rect 11020 24556 11022 24576
rect 10966 24520 11022 24556
rect 10874 24384 10930 24440
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10138 19216 10194 19272
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10782 20052 10838 20088
rect 10782 20032 10784 20052
rect 10784 20032 10836 20052
rect 10836 20032 10838 20052
rect 9770 18536 9826 18592
rect 9954 18400 10010 18456
rect 9678 16360 9734 16416
rect 9770 15272 9826 15328
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 11518 23160 11574 23216
rect 12162 24248 12218 24304
rect 11702 21936 11758 21992
rect 10966 18944 11022 19000
rect 10782 17856 10838 17912
rect 10690 17196 10746 17232
rect 10690 17176 10692 17196
rect 10692 17176 10744 17196
rect 10744 17176 10746 17196
rect 10782 16904 10838 16960
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10690 16088 10746 16144
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10138 15680 10194 15736
rect 10322 15444 10324 15464
rect 10324 15444 10376 15464
rect 10376 15444 10378 15464
rect 10322 15408 10378 15444
rect 10046 14476 10102 14512
rect 10046 14456 10048 14476
rect 10048 14456 10100 14476
rect 10100 14456 10102 14476
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10690 13524 10746 13560
rect 10690 13504 10692 13524
rect 10692 13504 10744 13524
rect 10744 13504 10746 13524
rect 9954 12960 10010 13016
rect 11150 16088 11206 16144
rect 10966 14728 11022 14784
rect 11610 17448 11666 17504
rect 11334 16088 11390 16144
rect 11794 19624 11850 19680
rect 12898 24656 12954 24712
rect 12806 23704 12862 23760
rect 12438 21664 12494 21720
rect 12162 20204 12164 20224
rect 12164 20204 12216 20224
rect 12216 20204 12218 20224
rect 12162 20168 12218 20204
rect 12990 23840 13046 23896
rect 12622 21800 12678 21856
rect 12162 18672 12218 18728
rect 12438 20032 12494 20088
rect 12346 19080 12402 19136
rect 11702 14864 11758 14920
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10138 12280 10194 12336
rect 10690 11872 10746 11928
rect 10138 11464 10194 11520
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 11518 12416 11574 12472
rect 10690 11328 10746 11384
rect 9494 10648 9550 10704
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 9218 9968 9274 10024
rect 11978 14048 12034 14104
rect 11886 13640 11942 13696
rect 12622 15272 12678 15328
rect 12438 13948 12440 13968
rect 12440 13948 12492 13968
rect 12492 13948 12494 13968
rect 12438 13912 12494 13948
rect 12162 13776 12218 13832
rect 13266 25356 13322 25392
rect 13266 25336 13268 25356
rect 13268 25336 13320 25356
rect 13320 25336 13322 25356
rect 13266 23296 13322 23352
rect 13082 22208 13138 22264
rect 12806 20476 12808 20496
rect 12808 20476 12860 20496
rect 12860 20476 12862 20496
rect 12806 20440 12862 20476
rect 12806 20168 12862 20224
rect 13082 17992 13138 18048
rect 13082 16904 13138 16960
rect 12990 16768 13046 16824
rect 12898 15136 12954 15192
rect 12806 14764 12808 14784
rect 12808 14764 12860 14784
rect 12860 14764 12862 14784
rect 12806 14728 12862 14764
rect 11702 9424 11758 9480
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 9586 9016 9642 9072
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 9586 6160 9642 6216
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 8850 3576 8906 3632
rect 12806 11192 12862 11248
rect 12438 3440 12494 3496
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 8298 2896 8354 2952
rect 12438 2896 12494 2952
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 12714 2508 12770 2544
rect 12714 2488 12716 2508
rect 12716 2488 12768 2508
rect 12768 2488 12770 2508
rect 4066 312 4122 368
rect 12990 13640 13046 13696
rect 12990 12008 13046 12064
rect 13266 21256 13322 21312
rect 13634 24404 13690 24440
rect 13634 24384 13636 24404
rect 13636 24384 13688 24404
rect 13688 24384 13690 24404
rect 13542 24112 13598 24168
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14370 24676 14426 24712
rect 14370 24656 14372 24676
rect 14372 24656 14424 24676
rect 14424 24656 14426 24676
rect 13450 21936 13506 21992
rect 13358 21120 13414 21176
rect 13542 21664 13598 21720
rect 13358 20576 13414 20632
rect 13358 17604 13414 17640
rect 13358 17584 13360 17604
rect 13360 17584 13412 17604
rect 13412 17584 13414 17604
rect 13450 17332 13506 17368
rect 13450 17312 13452 17332
rect 13452 17312 13504 17332
rect 13504 17312 13506 17332
rect 13542 16652 13598 16688
rect 13542 16632 13544 16652
rect 13544 16632 13596 16652
rect 13596 16632 13598 16652
rect 13726 23024 13782 23080
rect 14186 23024 14242 23080
rect 14186 22616 14242 22672
rect 13910 21972 13912 21992
rect 13912 21972 13964 21992
rect 13964 21972 13966 21992
rect 13910 21936 13966 21972
rect 14922 24828 14924 24848
rect 14924 24828 14976 24848
rect 14976 24828 14978 24848
rect 14922 24792 14978 24828
rect 15106 24792 15162 24848
rect 14554 21800 14610 21856
rect 15198 24248 15254 24304
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15474 24404 15530 24440
rect 15474 24384 15476 24404
rect 15476 24384 15528 24404
rect 15528 24384 15530 24404
rect 16854 25744 16910 25800
rect 15750 24656 15806 24712
rect 15658 24112 15714 24168
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15290 22208 15346 22264
rect 14738 21936 14794 21992
rect 13910 20168 13966 20224
rect 14462 21256 14518 21312
rect 13726 17584 13782 17640
rect 13818 17176 13874 17232
rect 14094 17992 14150 18048
rect 14186 17720 14242 17776
rect 13818 16496 13874 16552
rect 13818 13676 13820 13696
rect 13820 13676 13872 13696
rect 13872 13676 13874 13696
rect 13818 13640 13874 13676
rect 13358 13504 13414 13560
rect 13818 13252 13874 13288
rect 13818 13232 13820 13252
rect 13820 13232 13872 13252
rect 13872 13232 13874 13252
rect 13266 12824 13322 12880
rect 13174 12008 13230 12064
rect 13082 11500 13084 11520
rect 13084 11500 13136 11520
rect 13136 11500 13138 11520
rect 13082 11464 13138 11500
rect 13082 11056 13138 11112
rect 12990 9560 13046 9616
rect 13726 11636 13728 11656
rect 13728 11636 13780 11656
rect 13780 11636 13782 11656
rect 13726 11600 13782 11636
rect 14002 14048 14058 14104
rect 14462 20712 14518 20768
rect 14370 20168 14426 20224
rect 14462 20032 14518 20088
rect 14462 19760 14518 19816
rect 14370 19488 14426 19544
rect 14462 18828 14518 18864
rect 14462 18808 14464 18828
rect 14464 18808 14516 18828
rect 14516 18808 14518 18828
rect 14370 18536 14426 18592
rect 14370 18128 14426 18184
rect 14462 17992 14518 18048
rect 14646 19216 14702 19272
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14738 18944 14794 19000
rect 15566 21936 15622 21992
rect 14646 18808 14702 18864
rect 14554 17856 14610 17912
rect 14462 16496 14518 16552
rect 15382 18672 15438 18728
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14738 17856 14794 17912
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15106 17196 15162 17232
rect 15106 17176 15108 17196
rect 15108 17176 15160 17196
rect 15160 17176 15162 17196
rect 15014 17060 15070 17096
rect 15014 17040 15016 17060
rect 15016 17040 15068 17060
rect 15068 17040 15070 17060
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14554 16088 14610 16144
rect 14554 15544 14610 15600
rect 14278 13504 14334 13560
rect 14094 12552 14150 12608
rect 15382 16224 15438 16280
rect 15842 21292 15844 21312
rect 15844 21292 15896 21312
rect 15896 21292 15898 21312
rect 15842 21256 15898 21292
rect 15842 20868 15898 20904
rect 15842 20848 15844 20868
rect 15844 20848 15896 20868
rect 15896 20848 15898 20868
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15290 14592 15346 14648
rect 16394 24384 16450 24440
rect 16854 24928 16910 24984
rect 16670 22380 16672 22400
rect 16672 22380 16724 22400
rect 16724 22380 16726 22400
rect 16670 22344 16726 22380
rect 17314 23976 17370 24032
rect 16302 19080 16358 19136
rect 16394 18944 16450 19000
rect 16394 18128 16450 18184
rect 16210 17856 16266 17912
rect 16118 17720 16174 17776
rect 16302 17740 16358 17776
rect 16302 17720 16304 17740
rect 16304 17720 16356 17740
rect 16356 17720 16358 17740
rect 16118 17312 16174 17368
rect 16210 17040 16266 17096
rect 16394 16768 16450 16824
rect 15750 15816 15806 15872
rect 15566 15408 15622 15464
rect 15750 15408 15806 15464
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14830 12416 14886 12472
rect 14738 11620 14794 11656
rect 14738 11600 14740 11620
rect 14740 11600 14792 11620
rect 14792 11600 14794 11620
rect 14278 11056 14334 11112
rect 13450 10104 13506 10160
rect 13266 5480 13322 5536
rect 13726 5072 13782 5128
rect 13726 3984 13782 4040
rect 13910 3576 13966 3632
rect 13082 3440 13138 3496
rect 14554 9560 14610 9616
rect 14370 5616 14426 5672
rect 14186 5480 14242 5536
rect 14554 5208 14610 5264
rect 14738 9016 14794 9072
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15750 11620 15806 11656
rect 15750 11600 15752 11620
rect 15752 11600 15804 11620
rect 15804 11600 15806 11620
rect 16946 17856 17002 17912
rect 16302 14340 16358 14376
rect 16302 14320 16304 14340
rect 16304 14320 16356 14340
rect 16356 14320 16358 14340
rect 16670 14456 16726 14512
rect 17130 16088 17186 16144
rect 17038 15156 17094 15192
rect 17038 15136 17040 15156
rect 17040 15136 17092 15156
rect 17092 15136 17094 15156
rect 16854 13640 16910 13696
rect 16210 12280 16266 12336
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 16762 12960 16818 13016
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 16854 11076 16910 11112
rect 16854 11056 16856 11076
rect 16856 11056 16908 11076
rect 16908 11056 16910 11076
rect 17222 15972 17278 16008
rect 17222 15952 17224 15972
rect 17224 15952 17276 15972
rect 17276 15952 17278 15972
rect 17406 22500 17462 22536
rect 17406 22480 17408 22500
rect 17408 22480 17460 22500
rect 17460 22480 17462 22500
rect 17866 23568 17922 23624
rect 18050 22228 18106 22264
rect 18050 22208 18052 22228
rect 18052 22208 18104 22228
rect 18104 22208 18106 22228
rect 17774 21564 17776 21584
rect 17776 21564 17828 21584
rect 17828 21564 17830 21584
rect 17774 21528 17830 21564
rect 17590 21120 17646 21176
rect 17774 20304 17830 20360
rect 17590 18536 17646 18592
rect 18510 21392 18566 21448
rect 18234 19216 18290 19272
rect 17682 15952 17738 16008
rect 17222 15408 17278 15464
rect 17774 15272 17830 15328
rect 17774 14592 17830 14648
rect 17498 13232 17554 13288
rect 18418 19080 18474 19136
rect 18326 17856 18382 17912
rect 18234 17584 18290 17640
rect 17866 13504 17922 13560
rect 18050 13096 18106 13152
rect 18602 20712 18658 20768
rect 18694 18944 18750 19000
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19430 24656 19486 24712
rect 20166 24928 20222 24984
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19246 24248 19302 24304
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 20258 23704 20314 23760
rect 19522 22480 19578 22536
rect 19338 22344 19394 22400
rect 19062 20168 19118 20224
rect 19338 20032 19394 20088
rect 19338 18400 19394 18456
rect 19246 18264 19302 18320
rect 19062 17584 19118 17640
rect 18878 16632 18934 16688
rect 18786 16088 18842 16144
rect 18786 15816 18842 15872
rect 18694 15000 18750 15056
rect 18510 13096 18566 13152
rect 17866 11736 17922 11792
rect 17130 10920 17186 10976
rect 18694 12588 18696 12608
rect 18696 12588 18748 12608
rect 18748 12588 18750 12608
rect 18694 12552 18750 12588
rect 17958 9424 18014 9480
rect 18602 9424 18658 9480
rect 17958 7656 18014 7712
rect 17130 6840 17186 6896
rect 17314 6840 17370 6896
rect 19154 16632 19210 16688
rect 19062 16496 19118 16552
rect 19062 16088 19118 16144
rect 19246 15680 19302 15736
rect 18970 15000 19026 15056
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 20074 20032 20130 20088
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 20994 23296 21050 23352
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19430 13640 19486 13696
rect 18970 11056 19026 11112
rect 19982 14356 19984 14376
rect 19984 14356 20036 14376
rect 20036 14356 20038 14376
rect 19982 14320 20038 14356
rect 20258 14320 20314 14376
rect 20718 17584 20774 17640
rect 20442 13640 20498 13696
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 20718 15680 20774 15736
rect 20902 18672 20958 18728
rect 20626 12552 20682 12608
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19798 12180 19800 12200
rect 19800 12180 19852 12200
rect 19852 12180 19854 12200
rect 19798 12144 19854 12180
rect 20626 12008 20682 12064
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19338 8880 19394 8936
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19246 7928 19302 7984
rect 21270 23568 21326 23624
rect 21086 22752 21142 22808
rect 21178 22344 21234 22400
rect 21362 20712 21418 20768
rect 21178 20168 21234 20224
rect 21086 19216 21142 19272
rect 21086 18536 21142 18592
rect 20810 13232 20866 13288
rect 21362 18536 21418 18592
rect 21822 23024 21878 23080
rect 21546 20304 21602 20360
rect 21546 16632 21602 16688
rect 22006 23296 22062 23352
rect 22006 23024 22062 23080
rect 22006 22616 22062 22672
rect 21822 20748 21824 20768
rect 21824 20748 21876 20768
rect 21876 20748 21878 20768
rect 21822 20712 21878 20748
rect 22006 19932 22008 19952
rect 22008 19932 22060 19952
rect 22060 19932 22062 19952
rect 22006 19896 22062 19932
rect 21730 19352 21786 19408
rect 21730 16224 21786 16280
rect 21454 14184 21510 14240
rect 21086 12416 21142 12472
rect 20902 9968 20958 10024
rect 20994 9016 21050 9072
rect 20718 7384 20774 7440
rect 19062 7248 19118 7304
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 17314 6296 17370 6352
rect 18786 6296 18842 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 21638 13524 21694 13560
rect 21638 13504 21640 13524
rect 21640 13504 21692 13524
rect 21692 13504 21694 13524
rect 21822 15952 21878 16008
rect 22006 14728 22062 14784
rect 22558 22516 22560 22536
rect 22560 22516 22612 22536
rect 22612 22516 22614 22536
rect 22558 22480 22614 22516
rect 22558 22072 22614 22128
rect 22466 21392 22522 21448
rect 22282 18264 22338 18320
rect 22190 14592 22246 14648
rect 22466 16904 22522 16960
rect 22650 20440 22706 20496
rect 22650 20032 22706 20088
rect 22650 19760 22706 19816
rect 23018 19624 23074 19680
rect 22926 19216 22982 19272
rect 22834 18400 22890 18456
rect 22742 17856 22798 17912
rect 22466 16088 22522 16144
rect 21822 13776 21878 13832
rect 21914 12724 21916 12744
rect 21916 12724 21968 12744
rect 21968 12724 21970 12744
rect 21914 12688 21970 12724
rect 22374 13504 22430 13560
rect 22374 13232 22430 13288
rect 22282 11756 22338 11792
rect 22282 11736 22284 11756
rect 22284 11736 22336 11756
rect 22336 11736 22338 11756
rect 22374 11600 22430 11656
rect 22650 14592 22706 14648
rect 22558 13504 22614 13560
rect 22650 12980 22706 13016
rect 22650 12960 22652 12980
rect 22652 12960 22704 12980
rect 22704 12960 22706 12980
rect 22926 17992 22982 18048
rect 22926 17620 22928 17640
rect 22928 17620 22980 17640
rect 22980 17620 22982 17640
rect 22926 17584 22982 17620
rect 22926 17312 22982 17368
rect 22926 16088 22982 16144
rect 22926 14728 22982 14784
rect 22466 10104 22522 10160
rect 23110 15680 23166 15736
rect 24674 26424 24730 26480
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 23754 24792 23810 24848
rect 24214 24792 24270 24848
rect 23938 24268 23994 24304
rect 23938 24248 23940 24268
rect 23940 24248 23992 24268
rect 23992 24248 23994 24268
rect 23478 23976 23534 24032
rect 24766 25880 24822 25936
rect 24766 25200 24822 25256
rect 24674 23976 24730 24032
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 23846 23024 23902 23080
rect 23294 18420 23350 18456
rect 23294 18400 23296 18420
rect 23296 18400 23348 18420
rect 23348 18400 23350 18420
rect 23570 17720 23626 17776
rect 23754 18264 23810 18320
rect 23754 17856 23810 17912
rect 23386 16632 23442 16688
rect 23294 15680 23350 15736
rect 23386 15136 23442 15192
rect 23478 14884 23534 14920
rect 23478 14864 23480 14884
rect 23480 14864 23532 14884
rect 23532 14864 23534 14884
rect 23386 12416 23442 12472
rect 23018 11892 23074 11928
rect 23018 11872 23020 11892
rect 23020 11872 23072 11892
rect 23072 11872 23074 11892
rect 23662 17332 23718 17368
rect 23662 17312 23664 17332
rect 23664 17312 23716 17332
rect 23716 17312 23718 17332
rect 23662 16768 23718 16824
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24398 22616 24454 22672
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24766 22208 24822 22264
rect 25318 23180 25374 23216
rect 25318 23160 25320 23180
rect 25320 23160 25372 23180
rect 25372 23160 25374 23180
rect 25134 22380 25136 22400
rect 25136 22380 25188 22400
rect 25188 22380 25190 22400
rect 25134 22344 25190 22380
rect 24674 21528 24730 21584
rect 24122 20712 24178 20768
rect 24122 19760 24178 19816
rect 23846 15952 23902 16008
rect 23754 15272 23810 15328
rect 23662 14220 23664 14240
rect 23664 14220 23716 14240
rect 23716 14220 23718 14240
rect 23662 14184 23718 14220
rect 24030 17176 24086 17232
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24950 20848 25006 20904
rect 24766 20304 24822 20360
rect 25226 21936 25282 21992
rect 25042 19216 25098 19272
rect 25042 18808 25098 18864
rect 25042 17992 25098 18048
rect 24398 17740 24454 17776
rect 24398 17720 24400 17740
rect 24400 17720 24452 17740
rect 24452 17720 24454 17740
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24306 17176 24362 17232
rect 24858 17584 24914 17640
rect 24766 17448 24822 17504
rect 24766 17312 24822 17368
rect 24674 16940 24676 16960
rect 24676 16940 24728 16960
rect 24728 16940 24730 16960
rect 24674 16904 24730 16940
rect 24306 16768 24362 16824
rect 24674 16768 24730 16824
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24950 16768 25006 16824
rect 24950 16496 25006 16552
rect 24858 16396 24860 16416
rect 24860 16396 24912 16416
rect 24912 16396 24914 16416
rect 24858 16360 24914 16396
rect 24766 16088 24822 16144
rect 24766 15408 24822 15464
rect 24030 14456 24086 14512
rect 23754 12688 23810 12744
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24214 13912 24270 13968
rect 24214 13368 24270 13424
rect 23478 10920 23534 10976
rect 22926 9288 22982 9344
rect 23662 11192 23718 11248
rect 23570 10512 23626 10568
rect 23478 8880 23534 8936
rect 21270 7792 21326 7848
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24122 12824 24178 12880
rect 24398 12416 24454 12472
rect 23938 10104 23994 10160
rect 23846 9560 23902 9616
rect 23662 5752 23718 5808
rect 20994 5072 21050 5128
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 16394 4528 16450 4584
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 19522 3984 19578 4040
rect 14830 3576 14886 3632
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14646 2488 14702 2544
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 14186 1400 14242 1456
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24582 11328 24638 11384
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24398 10668 24454 10704
rect 24398 10648 24400 10668
rect 24400 10648 24452 10668
rect 24452 10648 24454 10668
rect 24858 13912 24914 13968
rect 25502 27104 25558 27160
rect 25502 23316 25558 23352
rect 25502 23296 25504 23316
rect 25504 23296 25556 23316
rect 25556 23296 25558 23316
rect 25778 22480 25834 22536
rect 25502 21528 25558 21584
rect 25226 17076 25228 17096
rect 25228 17076 25280 17096
rect 25280 17076 25282 17096
rect 25226 17040 25282 17076
rect 25042 15408 25098 15464
rect 25226 15544 25282 15600
rect 25594 20032 25650 20088
rect 25594 18148 25650 18184
rect 25594 18128 25596 18148
rect 25596 18128 25648 18148
rect 25648 18128 25650 18148
rect 25410 13776 25466 13832
rect 25318 12588 25320 12608
rect 25320 12588 25372 12608
rect 25372 12588 25374 12608
rect 25318 12552 25374 12588
rect 25134 12416 25190 12472
rect 25686 12144 25742 12200
rect 25870 13504 25926 13560
rect 24766 10104 24822 10160
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24674 9424 24730 9480
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24122 3848 24178 3904
rect 23478 3576 23534 3632
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 12898 40 12954 96
rect 24674 3440 24730 3496
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24122 2624 24178 2680
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25134 9460 25136 9480
rect 25136 9460 25188 9480
rect 25188 9460 25190 9480
rect 25134 9424 25190 9460
rect 26238 24656 26294 24712
rect 26330 19080 26386 19136
rect 26238 17856 26294 17912
rect 26238 17176 26294 17232
rect 26238 13096 26294 13152
rect 26146 10376 26202 10432
rect 27618 24384 27674 24440
rect 26422 6840 26478 6896
rect 24766 3304 24822 3360
rect 24674 2080 24730 2136
rect 23478 312 23534 368
<< metal3 >>
rect 0 27706 480 27736
rect 3509 27706 3575 27709
rect 0 27704 3575 27706
rect 0 27648 3514 27704
rect 3570 27648 3575 27704
rect 0 27646 3575 27648
rect 0 27616 480 27646
rect 3509 27643 3575 27646
rect 25589 27706 25655 27709
rect 27520 27706 28000 27736
rect 25589 27704 28000 27706
rect 25589 27648 25594 27704
rect 25650 27648 28000 27704
rect 25589 27646 28000 27648
rect 25589 27643 25655 27646
rect 27520 27616 28000 27646
rect 0 27162 480 27192
rect 3785 27162 3851 27165
rect 0 27160 3851 27162
rect 0 27104 3790 27160
rect 3846 27104 3851 27160
rect 0 27102 3851 27104
rect 0 27072 480 27102
rect 3785 27099 3851 27102
rect 25497 27162 25563 27165
rect 27520 27162 28000 27192
rect 25497 27160 28000 27162
rect 25497 27104 25502 27160
rect 25558 27104 28000 27160
rect 25497 27102 28000 27104
rect 25497 27099 25563 27102
rect 27520 27072 28000 27102
rect 0 26482 480 26512
rect 4061 26482 4127 26485
rect 0 26480 4127 26482
rect 0 26424 4066 26480
rect 4122 26424 4127 26480
rect 0 26422 4127 26424
rect 0 26392 480 26422
rect 4061 26419 4127 26422
rect 24669 26482 24735 26485
rect 27520 26482 28000 26512
rect 24669 26480 28000 26482
rect 24669 26424 24674 26480
rect 24730 26424 28000 26480
rect 24669 26422 28000 26424
rect 24669 26419 24735 26422
rect 27520 26392 28000 26422
rect 0 25938 480 25968
rect 2773 25938 2839 25941
rect 0 25936 2839 25938
rect 0 25880 2778 25936
rect 2834 25880 2839 25936
rect 0 25878 2839 25880
rect 0 25848 480 25878
rect 2773 25875 2839 25878
rect 24761 25938 24827 25941
rect 27520 25938 28000 25968
rect 24761 25936 28000 25938
rect 24761 25880 24766 25936
rect 24822 25880 28000 25936
rect 24761 25878 28000 25880
rect 24761 25875 24827 25878
rect 27520 25848 28000 25878
rect 4153 25802 4219 25805
rect 16849 25802 16915 25805
rect 4153 25800 16915 25802
rect 4153 25744 4158 25800
rect 4214 25744 16854 25800
rect 16910 25744 16915 25800
rect 4153 25742 16915 25744
rect 4153 25739 4219 25742
rect 16849 25739 16915 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 13118 25332 13124 25396
rect 13188 25394 13194 25396
rect 13261 25394 13327 25397
rect 13188 25392 13327 25394
rect 13188 25336 13266 25392
rect 13322 25336 13327 25392
rect 13188 25334 13327 25336
rect 13188 25332 13194 25334
rect 13261 25331 13327 25334
rect 0 25258 480 25288
rect 2681 25258 2747 25261
rect 0 25256 2747 25258
rect 0 25200 2686 25256
rect 2742 25200 2747 25256
rect 0 25198 2747 25200
rect 0 25168 480 25198
rect 2681 25195 2747 25198
rect 24761 25258 24827 25261
rect 27520 25258 28000 25288
rect 24761 25256 28000 25258
rect 24761 25200 24766 25256
rect 24822 25200 28000 25256
rect 24761 25198 28000 25200
rect 24761 25195 24827 25198
rect 27520 25168 28000 25198
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 2497 24986 2563 24989
rect 16849 24986 16915 24989
rect 20161 24986 20227 24989
rect 2497 24984 5504 24986
rect 2497 24928 2502 24984
rect 2558 24928 5504 24984
rect 2497 24926 5504 24928
rect 2497 24923 2563 24926
rect 5444 24850 5504 24926
rect 16849 24984 20227 24986
rect 16849 24928 16854 24984
rect 16910 24928 20166 24984
rect 20222 24928 20227 24984
rect 16849 24926 20227 24928
rect 16849 24923 16915 24926
rect 20161 24923 20227 24926
rect 14917 24850 14983 24853
rect 5444 24848 14983 24850
rect 5444 24792 14922 24848
rect 14978 24792 14983 24848
rect 5444 24790 14983 24792
rect 14917 24787 14983 24790
rect 15101 24850 15167 24853
rect 15101 24848 23306 24850
rect 15101 24792 15106 24848
rect 15162 24792 23306 24848
rect 15101 24790 23306 24792
rect 15101 24787 15167 24790
rect 0 24714 480 24744
rect 1577 24714 1643 24717
rect 0 24712 1643 24714
rect 0 24656 1582 24712
rect 1638 24656 1643 24712
rect 0 24654 1643 24656
rect 0 24624 480 24654
rect 1577 24651 1643 24654
rect 12893 24714 12959 24717
rect 14365 24714 14431 24717
rect 12893 24712 14431 24714
rect 12893 24656 12898 24712
rect 12954 24656 14370 24712
rect 14426 24656 14431 24712
rect 12893 24654 14431 24656
rect 12893 24651 12959 24654
rect 14365 24651 14431 24654
rect 15745 24714 15811 24717
rect 19425 24714 19491 24717
rect 15745 24712 19491 24714
rect 15745 24656 15750 24712
rect 15806 24656 19430 24712
rect 19486 24656 19491 24712
rect 15745 24654 19491 24656
rect 15745 24651 15811 24654
rect 19425 24651 19491 24654
rect 6085 24578 6151 24581
rect 9857 24578 9923 24581
rect 6085 24576 9923 24578
rect 6085 24520 6090 24576
rect 6146 24520 9862 24576
rect 9918 24520 9923 24576
rect 6085 24518 9923 24520
rect 6085 24515 6151 24518
rect 9857 24515 9923 24518
rect 10961 24578 11027 24581
rect 10961 24576 13922 24578
rect 10961 24520 10966 24576
rect 11022 24520 13922 24576
rect 10961 24518 13922 24520
rect 10961 24515 11027 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 2589 24442 2655 24445
rect 6913 24442 6979 24445
rect 2589 24440 6979 24442
rect 2589 24384 2594 24440
rect 2650 24384 6918 24440
rect 6974 24384 6979 24440
rect 2589 24382 6979 24384
rect 2589 24379 2655 24382
rect 6913 24379 6979 24382
rect 10869 24442 10935 24445
rect 13629 24442 13695 24445
rect 10869 24440 13695 24442
rect 10869 24384 10874 24440
rect 10930 24384 13634 24440
rect 13690 24384 13695 24440
rect 10869 24382 13695 24384
rect 13862 24442 13922 24518
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 15469 24442 15535 24445
rect 16389 24442 16455 24445
rect 13862 24440 15535 24442
rect 13862 24384 15474 24440
rect 15530 24384 15535 24440
rect 13862 24382 15535 24384
rect 10869 24379 10935 24382
rect 13629 24379 13695 24382
rect 15469 24379 15535 24382
rect 16254 24440 16455 24442
rect 16254 24384 16394 24440
rect 16450 24384 16455 24440
rect 16254 24382 16455 24384
rect 23246 24442 23306 24790
rect 23422 24788 23428 24852
rect 23492 24850 23498 24852
rect 23749 24850 23815 24853
rect 23492 24848 23815 24850
rect 23492 24792 23754 24848
rect 23810 24792 23815 24848
rect 23492 24790 23815 24792
rect 23492 24788 23498 24790
rect 23749 24787 23815 24790
rect 23974 24788 23980 24852
rect 24044 24850 24050 24852
rect 24209 24850 24275 24853
rect 24044 24848 24275 24850
rect 24044 24792 24214 24848
rect 24270 24792 24275 24848
rect 24044 24790 24275 24792
rect 24044 24788 24050 24790
rect 24209 24787 24275 24790
rect 26233 24714 26299 24717
rect 27520 24714 28000 24744
rect 26233 24712 28000 24714
rect 26233 24656 26238 24712
rect 26294 24656 28000 24712
rect 26233 24654 28000 24656
rect 26233 24651 26299 24654
rect 27520 24624 28000 24654
rect 27613 24442 27679 24445
rect 23246 24440 27679 24442
rect 23246 24384 27618 24440
rect 27674 24384 27679 24440
rect 23246 24382 27679 24384
rect 3233 24306 3299 24309
rect 8293 24306 8359 24309
rect 3233 24304 8359 24306
rect 3233 24248 3238 24304
rect 3294 24248 8298 24304
rect 8354 24248 8359 24304
rect 3233 24246 8359 24248
rect 3233 24243 3299 24246
rect 8293 24243 8359 24246
rect 9949 24306 10015 24309
rect 10910 24306 10916 24308
rect 9949 24304 10916 24306
rect 9949 24248 9954 24304
rect 10010 24248 10916 24304
rect 9949 24246 10916 24248
rect 9949 24243 10015 24246
rect 10910 24244 10916 24246
rect 10980 24244 10986 24308
rect 12157 24306 12223 24309
rect 15193 24306 15259 24309
rect 12157 24304 15259 24306
rect 12157 24248 12162 24304
rect 12218 24248 15198 24304
rect 15254 24248 15259 24304
rect 12157 24246 15259 24248
rect 12157 24243 12223 24246
rect 15193 24243 15259 24246
rect 3049 24170 3115 24173
rect 8937 24170 9003 24173
rect 13537 24172 13603 24173
rect 13486 24170 13492 24172
rect 3049 24168 7850 24170
rect 3049 24112 3054 24168
rect 3110 24112 7850 24168
rect 3049 24110 7850 24112
rect 3049 24107 3115 24110
rect 0 24034 480 24064
rect 3785 24034 3851 24037
rect 0 24032 3851 24034
rect 0 23976 3790 24032
rect 3846 23976 3851 24032
rect 0 23974 3851 23976
rect 7790 24034 7850 24110
rect 8937 24168 13492 24170
rect 13556 24168 13603 24172
rect 15653 24170 15719 24173
rect 16254 24170 16314 24382
rect 16389 24379 16455 24382
rect 27613 24379 27679 24382
rect 19241 24306 19307 24309
rect 23933 24306 23999 24309
rect 19241 24304 23999 24306
rect 19241 24248 19246 24304
rect 19302 24248 23938 24304
rect 23994 24248 23999 24304
rect 19241 24246 23999 24248
rect 19241 24243 19307 24246
rect 23933 24243 23999 24246
rect 8937 24112 8942 24168
rect 8998 24112 13492 24168
rect 13598 24112 13603 24168
rect 8937 24110 13492 24112
rect 8937 24107 9003 24110
rect 13486 24108 13492 24110
rect 13556 24108 13603 24112
rect 13537 24107 13603 24108
rect 14782 24168 16314 24170
rect 14782 24112 15658 24168
rect 15714 24112 16314 24168
rect 14782 24110 16314 24112
rect 14782 24034 14842 24110
rect 15653 24107 15719 24110
rect 7790 23974 14842 24034
rect 17309 24034 17375 24037
rect 23473 24034 23539 24037
rect 17309 24032 23539 24034
rect 17309 23976 17314 24032
rect 17370 23976 23478 24032
rect 23534 23976 23539 24032
rect 17309 23974 23539 23976
rect 0 23944 480 23974
rect 3785 23971 3851 23974
rect 17309 23971 17375 23974
rect 23473 23971 23539 23974
rect 24669 24034 24735 24037
rect 27520 24034 28000 24064
rect 24669 24032 28000 24034
rect 24669 23976 24674 24032
rect 24730 23976 28000 24032
rect 24669 23974 28000 23976
rect 24669 23971 24735 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 27520 23944 28000 23974
rect 24277 23903 24597 23904
rect 6453 23898 6519 23901
rect 8293 23898 8359 23901
rect 6453 23896 8359 23898
rect 6453 23840 6458 23896
rect 6514 23840 8298 23896
rect 8354 23840 8359 23896
rect 6453 23838 8359 23840
rect 6453 23835 6519 23838
rect 8293 23835 8359 23838
rect 10133 23898 10199 23901
rect 12985 23898 13051 23901
rect 10133 23896 13051 23898
rect 10133 23840 10138 23896
rect 10194 23840 12990 23896
rect 13046 23840 13051 23896
rect 10133 23838 13051 23840
rect 10133 23835 10199 23838
rect 12985 23835 13051 23838
rect 8845 23762 8911 23765
rect 12801 23762 12867 23765
rect 20253 23762 20319 23765
rect 8845 23760 12867 23762
rect 8845 23704 8850 23760
rect 8906 23704 12806 23760
rect 12862 23704 12867 23760
rect 8845 23702 12867 23704
rect 8845 23699 8911 23702
rect 12801 23699 12867 23702
rect 15334 23760 20319 23762
rect 15334 23704 20258 23760
rect 20314 23704 20319 23760
rect 15334 23702 20319 23704
rect 2221 23626 2287 23629
rect 5165 23626 5231 23629
rect 2221 23624 5231 23626
rect 2221 23568 2226 23624
rect 2282 23568 5170 23624
rect 5226 23568 5231 23624
rect 2221 23566 5231 23568
rect 2221 23563 2287 23566
rect 5165 23563 5231 23566
rect 0 23490 480 23520
rect 4061 23490 4127 23493
rect 0 23488 4127 23490
rect 0 23432 4066 23488
rect 4122 23432 4127 23488
rect 0 23430 4127 23432
rect 0 23400 480 23430
rect 4061 23427 4127 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 2405 23354 2471 23357
rect 7097 23354 7163 23357
rect 2405 23352 7163 23354
rect 2405 23296 2410 23352
rect 2466 23296 7102 23352
rect 7158 23296 7163 23352
rect 2405 23294 7163 23296
rect 2405 23291 2471 23294
rect 7097 23291 7163 23294
rect 7741 23354 7807 23357
rect 9765 23354 9831 23357
rect 7741 23352 9831 23354
rect 7741 23296 7746 23352
rect 7802 23296 9770 23352
rect 9826 23296 9831 23352
rect 7741 23294 9831 23296
rect 7741 23291 7807 23294
rect 9765 23291 9831 23294
rect 13261 23354 13327 23357
rect 15334 23354 15394 23702
rect 20253 23699 20319 23702
rect 17861 23626 17927 23629
rect 21265 23626 21331 23629
rect 17861 23624 21331 23626
rect 17861 23568 17866 23624
rect 17922 23568 21270 23624
rect 21326 23568 21331 23624
rect 17861 23566 21331 23568
rect 17861 23563 17927 23566
rect 21265 23563 21331 23566
rect 27520 23490 28000 23520
rect 25638 23430 28000 23490
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 13261 23352 15394 23354
rect 13261 23296 13266 23352
rect 13322 23296 15394 23352
rect 13261 23294 15394 23296
rect 20989 23354 21055 23357
rect 22001 23354 22067 23357
rect 20989 23352 22067 23354
rect 20989 23296 20994 23352
rect 21050 23296 22006 23352
rect 22062 23296 22067 23352
rect 20989 23294 22067 23296
rect 13261 23291 13327 23294
rect 20989 23291 21055 23294
rect 22001 23291 22067 23294
rect 25497 23354 25563 23357
rect 25638 23354 25698 23430
rect 27520 23400 28000 23430
rect 25497 23352 25698 23354
rect 25497 23296 25502 23352
rect 25558 23296 25698 23352
rect 25497 23294 25698 23296
rect 25497 23291 25563 23294
rect 8569 23218 8635 23221
rect 11513 23218 11579 23221
rect 25313 23218 25379 23221
rect 8569 23216 11579 23218
rect 8569 23160 8574 23216
rect 8630 23160 11518 23216
rect 11574 23160 11579 23216
rect 8569 23158 11579 23160
rect 8569 23155 8635 23158
rect 11513 23155 11579 23158
rect 13862 23216 25379 23218
rect 13862 23160 25318 23216
rect 25374 23160 25379 23216
rect 13862 23158 25379 23160
rect 13721 23082 13787 23085
rect 13862 23082 13922 23158
rect 25313 23155 25379 23158
rect 13721 23080 13922 23082
rect 13721 23024 13726 23080
rect 13782 23024 13922 23080
rect 13721 23022 13922 23024
rect 14181 23082 14247 23085
rect 21817 23082 21883 23085
rect 14181 23080 21883 23082
rect 14181 23024 14186 23080
rect 14242 23024 21822 23080
rect 21878 23024 21883 23080
rect 14181 23022 21883 23024
rect 13721 23019 13787 23022
rect 14181 23019 14247 23022
rect 21817 23019 21883 23022
rect 22001 23082 22067 23085
rect 23841 23082 23907 23085
rect 22001 23080 23907 23082
rect 22001 23024 22006 23080
rect 22062 23024 23846 23080
rect 23902 23024 23907 23080
rect 22001 23022 23907 23024
rect 22001 23019 22067 23022
rect 23841 23019 23907 23022
rect 9121 22946 9187 22949
rect 9121 22944 14842 22946
rect 9121 22888 9126 22944
rect 9182 22888 14842 22944
rect 9121 22886 14842 22888
rect 9121 22883 9187 22886
rect 5610 22880 5930 22881
rect 0 22810 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 2773 22810 2839 22813
rect 0 22808 2839 22810
rect 0 22752 2778 22808
rect 2834 22752 2839 22808
rect 0 22750 2839 22752
rect 0 22720 480 22750
rect 2773 22747 2839 22750
rect 3325 22674 3391 22677
rect 14181 22674 14247 22677
rect 3325 22672 14247 22674
rect 3325 22616 3330 22672
rect 3386 22616 14186 22672
rect 14242 22616 14247 22672
rect 3325 22614 14247 22616
rect 14782 22674 14842 22886
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 21081 22810 21147 22813
rect 27520 22810 28000 22840
rect 16990 22808 21147 22810
rect 16990 22752 21086 22808
rect 21142 22752 21147 22808
rect 16990 22750 21147 22752
rect 16990 22674 17050 22750
rect 21081 22747 21147 22750
rect 24718 22750 28000 22810
rect 22001 22674 22067 22677
rect 14782 22614 17050 22674
rect 17174 22672 22067 22674
rect 17174 22616 22006 22672
rect 22062 22616 22067 22672
rect 17174 22614 22067 22616
rect 3325 22611 3391 22614
rect 14181 22611 14247 22614
rect 7281 22538 7347 22541
rect 17174 22538 17234 22614
rect 22001 22611 22067 22614
rect 24393 22674 24459 22677
rect 24718 22674 24778 22750
rect 27520 22720 28000 22750
rect 24393 22672 24778 22674
rect 24393 22616 24398 22672
rect 24454 22616 24778 22672
rect 24393 22614 24778 22616
rect 24393 22611 24459 22614
rect 7281 22536 17234 22538
rect 7281 22480 7286 22536
rect 7342 22480 17234 22536
rect 7281 22478 17234 22480
rect 17401 22538 17467 22541
rect 19517 22538 19583 22541
rect 17401 22536 19583 22538
rect 17401 22480 17406 22536
rect 17462 22480 19522 22536
rect 19578 22480 19583 22536
rect 17401 22478 19583 22480
rect 7281 22475 7347 22478
rect 17401 22475 17467 22478
rect 19517 22475 19583 22478
rect 22553 22538 22619 22541
rect 25773 22538 25839 22541
rect 22553 22536 25839 22538
rect 22553 22480 22558 22536
rect 22614 22480 25778 22536
rect 25834 22480 25839 22536
rect 22553 22478 25839 22480
rect 22553 22475 22619 22478
rect 25773 22475 25839 22478
rect 4889 22402 4955 22405
rect 7189 22402 7255 22405
rect 4889 22400 7255 22402
rect 4889 22344 4894 22400
rect 4950 22344 7194 22400
rect 7250 22344 7255 22400
rect 4889 22342 7255 22344
rect 4889 22339 4955 22342
rect 7189 22339 7255 22342
rect 16665 22402 16731 22405
rect 19333 22402 19399 22405
rect 16665 22400 19399 22402
rect 16665 22344 16670 22400
rect 16726 22344 19338 22400
rect 19394 22344 19399 22400
rect 16665 22342 19399 22344
rect 16665 22339 16731 22342
rect 19333 22339 19399 22342
rect 21173 22402 21239 22405
rect 25129 22402 25195 22405
rect 21173 22400 25195 22402
rect 21173 22344 21178 22400
rect 21234 22344 25134 22400
rect 25190 22344 25195 22400
rect 21173 22342 25195 22344
rect 21173 22339 21239 22342
rect 25129 22339 25195 22342
rect 10277 22336 10597 22337
rect 0 22266 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 1577 22266 1643 22269
rect 0 22264 1643 22266
rect 0 22208 1582 22264
rect 1638 22208 1643 22264
rect 0 22206 1643 22208
rect 0 22176 480 22206
rect 1577 22203 1643 22206
rect 2497 22266 2563 22269
rect 2773 22266 2839 22269
rect 5441 22266 5507 22269
rect 8385 22266 8451 22269
rect 2497 22264 5320 22266
rect 2497 22208 2502 22264
rect 2558 22208 2778 22264
rect 2834 22208 5320 22264
rect 2497 22206 5320 22208
rect 2497 22203 2563 22206
rect 2773 22203 2839 22206
rect 5260 22130 5320 22206
rect 5441 22264 8451 22266
rect 5441 22208 5446 22264
rect 5502 22208 8390 22264
rect 8446 22208 8451 22264
rect 5441 22206 8451 22208
rect 5441 22203 5507 22206
rect 8385 22203 8451 22206
rect 13077 22266 13143 22269
rect 13302 22266 13308 22268
rect 13077 22264 13308 22266
rect 13077 22208 13082 22264
rect 13138 22208 13308 22264
rect 13077 22206 13308 22208
rect 13077 22203 13143 22206
rect 13302 22204 13308 22206
rect 13372 22204 13378 22268
rect 15285 22266 15351 22269
rect 18045 22266 18111 22269
rect 15285 22264 18111 22266
rect 15285 22208 15290 22264
rect 15346 22208 18050 22264
rect 18106 22208 18111 22264
rect 15285 22206 18111 22208
rect 15285 22203 15351 22206
rect 18045 22203 18111 22206
rect 24761 22266 24827 22269
rect 27520 22266 28000 22296
rect 24761 22264 28000 22266
rect 24761 22208 24766 22264
rect 24822 22208 28000 22264
rect 24761 22206 28000 22208
rect 24761 22203 24827 22206
rect 27520 22176 28000 22206
rect 22553 22130 22619 22133
rect 5260 22128 22619 22130
rect 5260 22072 22558 22128
rect 22614 22072 22619 22128
rect 5260 22070 22619 22072
rect 22553 22067 22619 22070
rect 1485 21994 1551 21997
rect 3233 21994 3299 21997
rect 1485 21992 3299 21994
rect 1485 21936 1490 21992
rect 1546 21936 3238 21992
rect 3294 21936 3299 21992
rect 1485 21934 3299 21936
rect 1485 21931 1551 21934
rect 3233 21931 3299 21934
rect 3877 21994 3943 21997
rect 6085 21994 6151 21997
rect 3877 21992 6151 21994
rect 3877 21936 3882 21992
rect 3938 21936 6090 21992
rect 6146 21936 6151 21992
rect 3877 21934 6151 21936
rect 3877 21931 3943 21934
rect 6085 21931 6151 21934
rect 8109 21994 8175 21997
rect 8753 21994 8819 21997
rect 9765 21994 9831 21997
rect 8109 21992 9831 21994
rect 8109 21936 8114 21992
rect 8170 21936 8758 21992
rect 8814 21936 9770 21992
rect 9826 21936 9831 21992
rect 8109 21934 9831 21936
rect 8109 21931 8175 21934
rect 8753 21931 8819 21934
rect 9765 21931 9831 21934
rect 11697 21994 11763 21997
rect 13445 21994 13511 21997
rect 13905 21994 13971 21997
rect 14733 21994 14799 21997
rect 11697 21992 14799 21994
rect 11697 21936 11702 21992
rect 11758 21936 13450 21992
rect 13506 21936 13910 21992
rect 13966 21936 14738 21992
rect 14794 21936 14799 21992
rect 11697 21934 14799 21936
rect 11697 21931 11763 21934
rect 13445 21931 13511 21934
rect 13905 21931 13971 21934
rect 14733 21931 14799 21934
rect 15561 21994 15627 21997
rect 25221 21994 25287 21997
rect 15561 21992 25287 21994
rect 15561 21936 15566 21992
rect 15622 21936 25226 21992
rect 25282 21936 25287 21992
rect 15561 21934 25287 21936
rect 15561 21931 15627 21934
rect 25221 21931 25287 21934
rect 12617 21858 12683 21861
rect 14549 21858 14615 21861
rect 7606 21856 14615 21858
rect 7606 21800 12622 21856
rect 12678 21800 14554 21856
rect 14610 21800 14615 21856
rect 7606 21798 14615 21800
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 2405 21722 2471 21725
rect 5257 21722 5323 21725
rect 2405 21720 5323 21722
rect 2405 21664 2410 21720
rect 2466 21664 5262 21720
rect 5318 21664 5323 21720
rect 2405 21662 5323 21664
rect 2405 21659 2471 21662
rect 5257 21659 5323 21662
rect 0 21586 480 21616
rect 2681 21586 2747 21589
rect 0 21584 2747 21586
rect 0 21528 2686 21584
rect 2742 21528 2747 21584
rect 0 21526 2747 21528
rect 0 21496 480 21526
rect 2681 21523 2747 21526
rect 2589 21450 2655 21453
rect 7606 21450 7666 21798
rect 12617 21795 12683 21798
rect 14549 21795 14615 21798
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 9121 21722 9187 21725
rect 12433 21722 12499 21725
rect 9121 21720 12499 21722
rect 9121 21664 9126 21720
rect 9182 21664 12438 21720
rect 12494 21664 12499 21720
rect 9121 21662 12499 21664
rect 9121 21659 9187 21662
rect 12433 21659 12499 21662
rect 13302 21660 13308 21724
rect 13372 21722 13378 21724
rect 13537 21722 13603 21725
rect 13372 21720 13603 21722
rect 13372 21664 13542 21720
rect 13598 21664 13603 21720
rect 13372 21662 13603 21664
rect 13372 21660 13378 21662
rect 13537 21659 13603 21662
rect 17769 21586 17835 21589
rect 2589 21448 7666 21450
rect 2589 21392 2594 21448
rect 2650 21392 7666 21448
rect 2589 21390 7666 21392
rect 7790 21584 17835 21586
rect 7790 21528 17774 21584
rect 17830 21528 17835 21584
rect 7790 21526 17835 21528
rect 2589 21387 2655 21390
rect 3601 21314 3667 21317
rect 7790 21314 7850 21526
rect 17769 21523 17835 21526
rect 24669 21586 24735 21589
rect 25497 21586 25563 21589
rect 27520 21586 28000 21616
rect 24669 21584 25563 21586
rect 24669 21528 24674 21584
rect 24730 21528 25502 21584
rect 25558 21528 25563 21584
rect 24669 21526 25563 21528
rect 24669 21523 24735 21526
rect 25497 21523 25563 21526
rect 25638 21526 28000 21586
rect 8385 21450 8451 21453
rect 18505 21450 18571 21453
rect 8385 21448 18571 21450
rect 8385 21392 8390 21448
rect 8446 21392 18510 21448
rect 18566 21392 18571 21448
rect 8385 21390 18571 21392
rect 8385 21387 8451 21390
rect 18505 21387 18571 21390
rect 22461 21450 22527 21453
rect 25638 21450 25698 21526
rect 27520 21496 28000 21526
rect 22461 21448 25698 21450
rect 22461 21392 22466 21448
rect 22522 21392 25698 21448
rect 22461 21390 25698 21392
rect 22461 21387 22527 21390
rect 3601 21312 7850 21314
rect 3601 21256 3606 21312
rect 3662 21256 7850 21312
rect 3601 21254 7850 21256
rect 8017 21314 8083 21317
rect 9673 21314 9739 21317
rect 8017 21312 9739 21314
rect 8017 21256 8022 21312
rect 8078 21256 9678 21312
rect 9734 21256 9739 21312
rect 8017 21254 9739 21256
rect 3601 21251 3667 21254
rect 8017 21251 8083 21254
rect 9673 21251 9739 21254
rect 13118 21252 13124 21316
rect 13188 21314 13194 21316
rect 13261 21314 13327 21317
rect 13188 21312 13327 21314
rect 13188 21256 13266 21312
rect 13322 21256 13327 21312
rect 13188 21254 13327 21256
rect 13188 21252 13194 21254
rect 13261 21251 13327 21254
rect 14457 21314 14523 21317
rect 15837 21314 15903 21317
rect 14457 21312 15903 21314
rect 14457 21256 14462 21312
rect 14518 21256 15842 21312
rect 15898 21256 15903 21312
rect 14457 21254 15903 21256
rect 14457 21251 14523 21254
rect 15837 21251 15903 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 7741 21178 7807 21181
rect 9765 21178 9831 21181
rect 7741 21176 9831 21178
rect 7741 21120 7746 21176
rect 7802 21120 9770 21176
rect 9826 21120 9831 21176
rect 7741 21118 9831 21120
rect 7741 21115 7807 21118
rect 9765 21115 9831 21118
rect 13353 21178 13419 21181
rect 17585 21178 17651 21181
rect 13353 21176 17651 21178
rect 13353 21120 13358 21176
rect 13414 21120 17590 21176
rect 17646 21120 17651 21176
rect 13353 21118 17651 21120
rect 13353 21115 13419 21118
rect 17585 21115 17651 21118
rect 0 21042 480 21072
rect 1393 21042 1459 21045
rect 0 21040 1459 21042
rect 0 20984 1398 21040
rect 1454 20984 1459 21040
rect 0 20982 1459 20984
rect 0 20952 480 20982
rect 1393 20979 1459 20982
rect 7097 21042 7163 21045
rect 14774 21042 14780 21044
rect 7097 21040 14780 21042
rect 7097 20984 7102 21040
rect 7158 20984 14780 21040
rect 7097 20982 14780 20984
rect 7097 20979 7163 20982
rect 14774 20980 14780 20982
rect 14844 20980 14850 21044
rect 24710 20980 24716 21044
rect 24780 21042 24786 21044
rect 27520 21042 28000 21072
rect 24780 20982 28000 21042
rect 24780 20980 24786 20982
rect 27520 20952 28000 20982
rect 3141 20906 3207 20909
rect 8385 20906 8451 20909
rect 3141 20904 8451 20906
rect 3141 20848 3146 20904
rect 3202 20848 8390 20904
rect 8446 20848 8451 20904
rect 3141 20846 8451 20848
rect 3141 20843 3207 20846
rect 8385 20843 8451 20846
rect 15837 20906 15903 20909
rect 24945 20906 25011 20909
rect 15837 20904 25011 20906
rect 15837 20848 15842 20904
rect 15898 20848 24950 20904
rect 25006 20848 25011 20904
rect 15837 20846 25011 20848
rect 15837 20843 15903 20846
rect 24945 20843 25011 20846
rect 6637 20770 6703 20773
rect 14457 20770 14523 20773
rect 6637 20768 14523 20770
rect 6637 20712 6642 20768
rect 6698 20712 14462 20768
rect 14518 20712 14523 20768
rect 6637 20710 14523 20712
rect 6637 20707 6703 20710
rect 14457 20707 14523 20710
rect 18597 20770 18663 20773
rect 21357 20770 21423 20773
rect 18597 20768 21423 20770
rect 18597 20712 18602 20768
rect 18658 20712 21362 20768
rect 21418 20712 21423 20768
rect 18597 20710 21423 20712
rect 18597 20707 18663 20710
rect 21357 20707 21423 20710
rect 21817 20770 21883 20773
rect 24117 20770 24183 20773
rect 21817 20768 24183 20770
rect 21817 20712 21822 20768
rect 21878 20712 24122 20768
rect 24178 20712 24183 20768
rect 21817 20710 24183 20712
rect 21817 20707 21883 20710
rect 24117 20707 24183 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 5993 20634 6059 20637
rect 9029 20634 9095 20637
rect 5993 20632 9095 20634
rect 5993 20576 5998 20632
rect 6054 20576 9034 20632
rect 9090 20576 9095 20632
rect 5993 20574 9095 20576
rect 5993 20571 6059 20574
rect 3601 20498 3667 20501
rect 6134 20498 6194 20574
rect 9029 20571 9095 20574
rect 13353 20634 13419 20637
rect 13486 20634 13492 20636
rect 13353 20632 13492 20634
rect 13353 20576 13358 20632
rect 13414 20576 13492 20632
rect 13353 20574 13492 20576
rect 13353 20571 13419 20574
rect 13486 20572 13492 20574
rect 13556 20572 13562 20636
rect 3601 20496 6194 20498
rect 3601 20440 3606 20496
rect 3662 20440 6194 20496
rect 3601 20438 6194 20440
rect 7557 20498 7623 20501
rect 12014 20498 12020 20500
rect 7557 20496 12020 20498
rect 7557 20440 7562 20496
rect 7618 20440 12020 20496
rect 7557 20438 12020 20440
rect 3601 20435 3667 20438
rect 7557 20435 7623 20438
rect 12014 20436 12020 20438
rect 12084 20436 12090 20500
rect 12801 20498 12867 20501
rect 22645 20498 22711 20501
rect 12801 20496 22711 20498
rect 12801 20440 12806 20496
rect 12862 20440 22650 20496
rect 22706 20440 22711 20496
rect 12801 20438 22711 20440
rect 12801 20435 12867 20438
rect 22645 20435 22711 20438
rect 0 20362 480 20392
rect 1669 20362 1735 20365
rect 0 20360 1735 20362
rect 0 20304 1674 20360
rect 1730 20304 1735 20360
rect 0 20302 1735 20304
rect 0 20272 480 20302
rect 1669 20299 1735 20302
rect 4245 20362 4311 20365
rect 17769 20362 17835 20365
rect 4245 20360 17835 20362
rect 4245 20304 4250 20360
rect 4306 20304 17774 20360
rect 17830 20304 17835 20360
rect 4245 20302 17835 20304
rect 4245 20299 4311 20302
rect 17769 20299 17835 20302
rect 21541 20362 21607 20365
rect 24761 20362 24827 20365
rect 27520 20362 28000 20392
rect 21541 20360 24827 20362
rect 21541 20304 21546 20360
rect 21602 20304 24766 20360
rect 24822 20304 24827 20360
rect 21541 20302 24827 20304
rect 21541 20299 21607 20302
rect 24761 20299 24827 20302
rect 24902 20302 28000 20362
rect 2037 20226 2103 20229
rect 6637 20226 6703 20229
rect 2037 20224 6703 20226
rect 2037 20168 2042 20224
rect 2098 20168 6642 20224
rect 6698 20168 6703 20224
rect 2037 20166 6703 20168
rect 2037 20163 2103 20166
rect 6637 20163 6703 20166
rect 12157 20226 12223 20229
rect 12801 20226 12867 20229
rect 13905 20226 13971 20229
rect 12157 20224 13971 20226
rect 12157 20168 12162 20224
rect 12218 20168 12806 20224
rect 12862 20168 13910 20224
rect 13966 20168 13971 20224
rect 12157 20166 13971 20168
rect 12157 20163 12223 20166
rect 12801 20163 12867 20166
rect 13905 20163 13971 20166
rect 14365 20226 14431 20229
rect 19057 20226 19123 20229
rect 14365 20224 19123 20226
rect 14365 20168 14370 20224
rect 14426 20168 19062 20224
rect 19118 20168 19123 20224
rect 14365 20166 19123 20168
rect 14365 20163 14431 20166
rect 19057 20163 19123 20166
rect 21173 20226 21239 20229
rect 24902 20226 24962 20302
rect 27520 20272 28000 20302
rect 21173 20224 24962 20226
rect 21173 20168 21178 20224
rect 21234 20168 24962 20224
rect 21173 20166 24962 20168
rect 21173 20163 21239 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 10777 20090 10843 20093
rect 12433 20090 12499 20093
rect 10777 20088 12499 20090
rect 10777 20032 10782 20088
rect 10838 20032 12438 20088
rect 12494 20032 12499 20088
rect 10777 20030 12499 20032
rect 10777 20027 10843 20030
rect 12433 20027 12499 20030
rect 14457 20090 14523 20093
rect 19333 20090 19399 20093
rect 14457 20088 19399 20090
rect 14457 20032 14462 20088
rect 14518 20032 19338 20088
rect 19394 20032 19399 20088
rect 14457 20030 19399 20032
rect 14457 20027 14523 20030
rect 19333 20027 19399 20030
rect 20069 20090 20135 20093
rect 22645 20090 22711 20093
rect 25589 20090 25655 20093
rect 20069 20088 25655 20090
rect 20069 20032 20074 20088
rect 20130 20032 22650 20088
rect 22706 20032 25594 20088
rect 25650 20032 25655 20088
rect 20069 20030 25655 20032
rect 20069 20027 20135 20030
rect 22645 20027 22711 20030
rect 25589 20027 25655 20030
rect 3233 19954 3299 19957
rect 7189 19954 7255 19957
rect 22001 19954 22067 19957
rect 22686 19954 22692 19956
rect 3233 19952 7114 19954
rect 3233 19896 3238 19952
rect 3294 19896 7114 19952
rect 3233 19894 7114 19896
rect 3233 19891 3299 19894
rect 0 19818 480 19848
rect 1577 19818 1643 19821
rect 0 19816 1643 19818
rect 0 19760 1582 19816
rect 1638 19760 1643 19816
rect 0 19758 1643 19760
rect 0 19728 480 19758
rect 1577 19755 1643 19758
rect 3417 19818 3483 19821
rect 6913 19818 6979 19821
rect 3417 19816 6979 19818
rect 3417 19760 3422 19816
rect 3478 19760 6918 19816
rect 6974 19760 6979 19816
rect 3417 19758 6979 19760
rect 7054 19818 7114 19894
rect 7189 19952 17280 19954
rect 7189 19896 7194 19952
rect 7250 19896 17280 19952
rect 7189 19894 17280 19896
rect 7189 19891 7255 19894
rect 14457 19818 14523 19821
rect 7054 19816 14523 19818
rect 7054 19760 14462 19816
rect 14518 19760 14523 19816
rect 7054 19758 14523 19760
rect 3417 19755 3483 19758
rect 6913 19755 6979 19758
rect 14457 19755 14523 19758
rect 14774 19756 14780 19820
rect 14844 19818 14850 19820
rect 17220 19818 17280 19894
rect 22001 19952 22692 19954
rect 22001 19896 22006 19952
rect 22062 19896 22692 19952
rect 22001 19894 22692 19896
rect 22001 19891 22067 19894
rect 22686 19892 22692 19894
rect 22756 19892 22762 19956
rect 22645 19818 22711 19821
rect 14844 19758 15394 19818
rect 17220 19816 22711 19818
rect 17220 19760 22650 19816
rect 22706 19760 22711 19816
rect 17220 19758 22711 19760
rect 14844 19756 14850 19758
rect 11789 19682 11855 19685
rect 8388 19680 11855 19682
rect 8388 19624 11794 19680
rect 11850 19624 11855 19680
rect 8388 19622 11855 19624
rect 15334 19682 15394 19758
rect 22645 19755 22711 19758
rect 24117 19818 24183 19821
rect 27520 19818 28000 19848
rect 24117 19816 28000 19818
rect 24117 19760 24122 19816
rect 24178 19760 28000 19816
rect 24117 19758 28000 19760
rect 24117 19755 24183 19758
rect 27520 19728 28000 19758
rect 23013 19682 23079 19685
rect 15334 19680 23079 19682
rect 15334 19624 23018 19680
rect 23074 19624 23079 19680
rect 15334 19622 23079 19624
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 3693 19410 3759 19413
rect 7557 19410 7623 19413
rect 3693 19408 7623 19410
rect 3693 19352 3698 19408
rect 3754 19352 7562 19408
rect 7618 19352 7623 19408
rect 3693 19350 7623 19352
rect 3693 19347 3759 19350
rect 7557 19347 7623 19350
rect 1945 19274 2011 19277
rect 5993 19274 6059 19277
rect 1945 19272 6059 19274
rect 1945 19216 1950 19272
rect 2006 19216 5998 19272
rect 6054 19216 6059 19272
rect 1945 19214 6059 19216
rect 1945 19211 2011 19214
rect 5993 19211 6059 19214
rect 0 19138 480 19168
rect 3601 19138 3667 19141
rect 0 19136 3667 19138
rect 0 19080 3606 19136
rect 3662 19080 3667 19136
rect 0 19078 3667 19080
rect 0 19048 480 19078
rect 3601 19075 3667 19078
rect 3877 19138 3943 19141
rect 8388 19138 8448 19622
rect 11789 19619 11855 19622
rect 23013 19619 23079 19622
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 12014 19484 12020 19548
rect 12084 19546 12090 19548
rect 14365 19546 14431 19549
rect 12084 19544 14431 19546
rect 12084 19488 14370 19544
rect 14426 19488 14431 19544
rect 12084 19486 14431 19488
rect 12084 19484 12090 19486
rect 14365 19483 14431 19486
rect 8569 19410 8635 19413
rect 21725 19410 21791 19413
rect 8569 19408 21791 19410
rect 8569 19352 8574 19408
rect 8630 19352 21730 19408
rect 21786 19352 21791 19408
rect 8569 19350 21791 19352
rect 8569 19347 8635 19350
rect 21725 19347 21791 19350
rect 10133 19274 10199 19277
rect 14641 19274 14707 19277
rect 10133 19272 14707 19274
rect 10133 19216 10138 19272
rect 10194 19216 14646 19272
rect 14702 19216 14707 19272
rect 10133 19214 14707 19216
rect 10133 19211 10199 19214
rect 14641 19211 14707 19214
rect 18229 19274 18295 19277
rect 21081 19274 21147 19277
rect 18229 19272 21147 19274
rect 18229 19216 18234 19272
rect 18290 19216 21086 19272
rect 21142 19216 21147 19272
rect 18229 19214 21147 19216
rect 18229 19211 18295 19214
rect 21081 19211 21147 19214
rect 22921 19274 22987 19277
rect 25037 19274 25103 19277
rect 22921 19272 25103 19274
rect 22921 19216 22926 19272
rect 22982 19216 25042 19272
rect 25098 19216 25103 19272
rect 22921 19214 25103 19216
rect 22921 19211 22987 19214
rect 25037 19211 25103 19214
rect 3877 19136 8448 19138
rect 3877 19080 3882 19136
rect 3938 19080 8448 19136
rect 3877 19078 8448 19080
rect 12341 19138 12407 19141
rect 16297 19138 16363 19141
rect 18413 19138 18479 19141
rect 12341 19136 18479 19138
rect 12341 19080 12346 19136
rect 12402 19080 16302 19136
rect 16358 19080 18418 19136
rect 18474 19080 18479 19136
rect 12341 19078 18479 19080
rect 3877 19075 3943 19078
rect 12341 19075 12407 19078
rect 16297 19075 16363 19078
rect 18413 19075 18479 19078
rect 26325 19138 26391 19141
rect 27520 19138 28000 19168
rect 26325 19136 28000 19138
rect 26325 19080 26330 19136
rect 26386 19080 28000 19136
rect 26325 19078 28000 19080
rect 26325 19075 26391 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19078
rect 19610 19007 19930 19008
rect 10961 19002 11027 19005
rect 14733 19002 14799 19005
rect 10961 19000 14799 19002
rect 10961 18944 10966 19000
rect 11022 18944 14738 19000
rect 14794 18944 14799 19000
rect 10961 18942 14799 18944
rect 10961 18939 11027 18942
rect 14733 18939 14799 18942
rect 16389 19002 16455 19005
rect 18689 19002 18755 19005
rect 16389 19000 18755 19002
rect 16389 18944 16394 19000
rect 16450 18944 18694 19000
rect 18750 18944 18755 19000
rect 16389 18942 18755 18944
rect 16389 18939 16455 18942
rect 18689 18939 18755 18942
rect 8569 18866 8635 18869
rect 14457 18866 14523 18869
rect 8569 18864 14523 18866
rect 8569 18808 8574 18864
rect 8630 18808 14462 18864
rect 14518 18808 14523 18864
rect 8569 18806 14523 18808
rect 8569 18803 8635 18806
rect 14457 18803 14523 18806
rect 14641 18866 14707 18869
rect 25037 18866 25103 18869
rect 14641 18864 25103 18866
rect 14641 18808 14646 18864
rect 14702 18808 25042 18864
rect 25098 18808 25103 18864
rect 14641 18806 25103 18808
rect 14641 18803 14707 18806
rect 25037 18803 25103 18806
rect 7281 18730 7347 18733
rect 12157 18730 12223 18733
rect 7281 18728 12223 18730
rect 7281 18672 7286 18728
rect 7342 18672 12162 18728
rect 12218 18672 12223 18728
rect 7281 18670 12223 18672
rect 7281 18667 7347 18670
rect 12157 18667 12223 18670
rect 15377 18730 15443 18733
rect 20897 18730 20963 18733
rect 15377 18728 20963 18730
rect 15377 18672 15382 18728
rect 15438 18672 20902 18728
rect 20958 18672 20963 18728
rect 15377 18670 20963 18672
rect 15377 18667 15443 18670
rect 20897 18667 20963 18670
rect 0 18594 480 18624
rect 4245 18594 4311 18597
rect 0 18592 4311 18594
rect 0 18536 4250 18592
rect 4306 18536 4311 18592
rect 0 18534 4311 18536
rect 0 18504 480 18534
rect 4245 18531 4311 18534
rect 9765 18594 9831 18597
rect 14365 18594 14431 18597
rect 9765 18592 14431 18594
rect 9765 18536 9770 18592
rect 9826 18536 14370 18592
rect 14426 18536 14431 18592
rect 9765 18534 14431 18536
rect 9765 18531 9831 18534
rect 14365 18531 14431 18534
rect 17585 18594 17651 18597
rect 21081 18594 21147 18597
rect 21357 18594 21423 18597
rect 27520 18594 28000 18624
rect 17585 18592 21423 18594
rect 17585 18536 17590 18592
rect 17646 18536 21086 18592
rect 21142 18536 21362 18592
rect 21418 18536 21423 18592
rect 17585 18534 21423 18536
rect 17585 18531 17651 18534
rect 21081 18531 21147 18534
rect 21357 18531 21423 18534
rect 24718 18534 28000 18594
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 7925 18458 7991 18461
rect 9949 18458 10015 18461
rect 7925 18456 10015 18458
rect 7925 18400 7930 18456
rect 7986 18400 9954 18456
rect 10010 18400 10015 18456
rect 7925 18398 10015 18400
rect 7925 18395 7991 18398
rect 9949 18395 10015 18398
rect 19333 18458 19399 18461
rect 22829 18458 22895 18461
rect 23289 18458 23355 18461
rect 19333 18456 23355 18458
rect 19333 18400 19338 18456
rect 19394 18400 22834 18456
rect 22890 18400 23294 18456
rect 23350 18400 23355 18456
rect 19333 18398 23355 18400
rect 19333 18395 19399 18398
rect 22829 18395 22895 18398
rect 23289 18395 23355 18398
rect 2957 18322 3023 18325
rect 6821 18322 6887 18325
rect 2957 18320 6887 18322
rect 2957 18264 2962 18320
rect 3018 18264 6826 18320
rect 6882 18264 6887 18320
rect 2957 18262 6887 18264
rect 2957 18259 3023 18262
rect 6821 18259 6887 18262
rect 19241 18322 19307 18325
rect 22277 18322 22343 18325
rect 19241 18320 22343 18322
rect 19241 18264 19246 18320
rect 19302 18264 22282 18320
rect 22338 18264 22343 18320
rect 19241 18262 22343 18264
rect 19241 18259 19307 18262
rect 22277 18259 22343 18262
rect 23749 18322 23815 18325
rect 24718 18322 24778 18534
rect 27520 18504 28000 18534
rect 23749 18320 24778 18322
rect 23749 18264 23754 18320
rect 23810 18264 24778 18320
rect 23749 18262 24778 18264
rect 23749 18259 23815 18262
rect 2497 18186 2563 18189
rect 6085 18186 6151 18189
rect 2497 18184 6151 18186
rect 2497 18128 2502 18184
rect 2558 18128 6090 18184
rect 6146 18128 6151 18184
rect 2497 18126 6151 18128
rect 2497 18123 2563 18126
rect 6085 18123 6151 18126
rect 8017 18186 8083 18189
rect 14365 18186 14431 18189
rect 8017 18184 14431 18186
rect 8017 18128 8022 18184
rect 8078 18128 14370 18184
rect 14426 18128 14431 18184
rect 8017 18126 14431 18128
rect 8017 18123 8083 18126
rect 14365 18123 14431 18126
rect 16389 18186 16455 18189
rect 25589 18186 25655 18189
rect 16389 18184 25655 18186
rect 16389 18128 16394 18184
rect 16450 18128 25594 18184
rect 25650 18128 25655 18184
rect 16389 18126 25655 18128
rect 16389 18123 16455 18126
rect 25589 18123 25655 18126
rect 4061 18050 4127 18053
rect 7097 18050 7163 18053
rect 4061 18048 7163 18050
rect 4061 17992 4066 18048
rect 4122 17992 7102 18048
rect 7158 17992 7163 18048
rect 4061 17990 7163 17992
rect 4061 17987 4127 17990
rect 7097 17987 7163 17990
rect 13077 18050 13143 18053
rect 14089 18050 14155 18053
rect 14457 18050 14523 18053
rect 13077 18048 14523 18050
rect 13077 17992 13082 18048
rect 13138 17992 14094 18048
rect 14150 17992 14462 18048
rect 14518 17992 14523 18048
rect 13077 17990 14523 17992
rect 13077 17987 13143 17990
rect 14089 17987 14155 17990
rect 14457 17987 14523 17990
rect 22921 18050 22987 18053
rect 25037 18050 25103 18053
rect 22921 18048 25103 18050
rect 22921 17992 22926 18048
rect 22982 17992 25042 18048
rect 25098 17992 25103 18048
rect 22921 17990 25103 17992
rect 22921 17987 22987 17990
rect 25037 17987 25103 17990
rect 10277 17984 10597 17985
rect 0 17914 480 17944
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 3693 17914 3759 17917
rect 0 17912 3759 17914
rect 0 17856 3698 17912
rect 3754 17856 3759 17912
rect 0 17854 3759 17856
rect 0 17824 480 17854
rect 3693 17851 3759 17854
rect 10777 17914 10843 17917
rect 14549 17914 14615 17917
rect 10777 17912 14615 17914
rect 10777 17856 10782 17912
rect 10838 17856 14554 17912
rect 14610 17856 14615 17912
rect 10777 17854 14615 17856
rect 10777 17851 10843 17854
rect 14549 17851 14615 17854
rect 14733 17914 14799 17917
rect 16205 17914 16271 17917
rect 14733 17912 16271 17914
rect 14733 17856 14738 17912
rect 14794 17856 16210 17912
rect 16266 17856 16271 17912
rect 14733 17854 16271 17856
rect 14733 17851 14799 17854
rect 16205 17851 16271 17854
rect 16941 17914 17007 17917
rect 18321 17914 18387 17917
rect 16941 17912 18387 17914
rect 16941 17856 16946 17912
rect 17002 17856 18326 17912
rect 18382 17856 18387 17912
rect 16941 17854 18387 17856
rect 16941 17851 17007 17854
rect 18321 17851 18387 17854
rect 22737 17914 22803 17917
rect 23749 17914 23815 17917
rect 22737 17912 23815 17914
rect 22737 17856 22742 17912
rect 22798 17856 23754 17912
rect 23810 17856 23815 17912
rect 22737 17854 23815 17856
rect 22737 17851 22803 17854
rect 23749 17851 23815 17854
rect 26233 17914 26299 17917
rect 27520 17914 28000 17944
rect 26233 17912 28000 17914
rect 26233 17856 26238 17912
rect 26294 17856 28000 17912
rect 26233 17854 28000 17856
rect 26233 17851 26299 17854
rect 27520 17824 28000 17854
rect 8753 17778 8819 17781
rect 14181 17778 14247 17781
rect 16113 17778 16179 17781
rect 8753 17776 14247 17778
rect 8753 17720 8758 17776
rect 8814 17720 14186 17776
rect 14242 17720 14247 17776
rect 8753 17718 14247 17720
rect 8753 17715 8819 17718
rect 14181 17715 14247 17718
rect 14414 17776 16179 17778
rect 14414 17720 16118 17776
rect 16174 17720 16179 17776
rect 14414 17718 16179 17720
rect 3417 17642 3483 17645
rect 13353 17642 13419 17645
rect 3417 17640 13419 17642
rect 3417 17584 3422 17640
rect 3478 17584 13358 17640
rect 13414 17584 13419 17640
rect 3417 17582 13419 17584
rect 3417 17579 3483 17582
rect 13353 17579 13419 17582
rect 13721 17642 13787 17645
rect 14414 17642 14474 17718
rect 16113 17715 16179 17718
rect 16297 17778 16363 17781
rect 23565 17778 23631 17781
rect 16297 17776 23631 17778
rect 16297 17720 16302 17776
rect 16358 17720 23570 17776
rect 23626 17720 23631 17776
rect 16297 17718 23631 17720
rect 16297 17715 16363 17718
rect 23565 17715 23631 17718
rect 23974 17716 23980 17780
rect 24044 17778 24050 17780
rect 24393 17778 24459 17781
rect 24044 17776 24459 17778
rect 24044 17720 24398 17776
rect 24454 17720 24459 17776
rect 24044 17718 24459 17720
rect 24044 17716 24050 17718
rect 24393 17715 24459 17718
rect 18229 17642 18295 17645
rect 13721 17640 14474 17642
rect 13721 17584 13726 17640
rect 13782 17584 14474 17640
rect 13721 17582 14474 17584
rect 14782 17640 18295 17642
rect 14782 17584 18234 17640
rect 18290 17584 18295 17640
rect 14782 17582 18295 17584
rect 13721 17579 13787 17582
rect 11605 17506 11671 17509
rect 14782 17506 14842 17582
rect 18229 17579 18295 17582
rect 19057 17642 19123 17645
rect 20713 17642 20779 17645
rect 19057 17640 20779 17642
rect 19057 17584 19062 17640
rect 19118 17584 20718 17640
rect 20774 17584 20779 17640
rect 19057 17582 20779 17584
rect 19057 17579 19123 17582
rect 20713 17579 20779 17582
rect 22921 17642 22987 17645
rect 24853 17642 24919 17645
rect 22921 17640 24919 17642
rect 22921 17584 22926 17640
rect 22982 17584 24858 17640
rect 24914 17584 24919 17640
rect 22921 17582 24919 17584
rect 22921 17579 22987 17582
rect 24853 17579 24919 17582
rect 2638 17446 5412 17506
rect 0 17370 480 17400
rect 2638 17370 2698 17446
rect 0 17310 2698 17370
rect 0 17280 480 17310
rect 5352 17234 5412 17446
rect 11605 17504 14842 17506
rect 11605 17448 11610 17504
rect 11666 17448 14842 17504
rect 11605 17446 14842 17448
rect 24761 17506 24827 17509
rect 24894 17506 24900 17508
rect 24761 17504 24900 17506
rect 24761 17448 24766 17504
rect 24822 17448 24900 17504
rect 24761 17446 24900 17448
rect 11605 17443 11671 17446
rect 24761 17443 24827 17446
rect 24894 17444 24900 17446
rect 24964 17444 24970 17508
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 6637 17370 6703 17373
rect 13445 17370 13511 17373
rect 6637 17368 13511 17370
rect 6637 17312 6642 17368
rect 6698 17312 13450 17368
rect 13506 17312 13511 17368
rect 6637 17310 13511 17312
rect 6637 17307 6703 17310
rect 13445 17307 13511 17310
rect 16113 17370 16179 17373
rect 22921 17370 22987 17373
rect 16113 17368 22987 17370
rect 16113 17312 16118 17368
rect 16174 17312 22926 17368
rect 22982 17312 22987 17368
rect 16113 17310 22987 17312
rect 16113 17307 16179 17310
rect 22921 17307 22987 17310
rect 23054 17308 23060 17372
rect 23124 17370 23130 17372
rect 23657 17370 23723 17373
rect 23124 17368 23723 17370
rect 23124 17312 23662 17368
rect 23718 17312 23723 17368
rect 23124 17310 23723 17312
rect 23124 17308 23130 17310
rect 23657 17307 23723 17310
rect 24761 17370 24827 17373
rect 27520 17370 28000 17400
rect 24761 17368 28000 17370
rect 24761 17312 24766 17368
rect 24822 17312 28000 17368
rect 24761 17310 28000 17312
rect 24761 17307 24827 17310
rect 27520 17280 28000 17310
rect 6913 17234 6979 17237
rect 5352 17232 6979 17234
rect 5352 17176 6918 17232
rect 6974 17176 6979 17232
rect 5352 17174 6979 17176
rect 6913 17171 6979 17174
rect 10685 17234 10751 17237
rect 13813 17234 13879 17237
rect 10685 17232 13879 17234
rect 10685 17176 10690 17232
rect 10746 17176 13818 17232
rect 13874 17176 13879 17232
rect 10685 17174 13879 17176
rect 10685 17171 10751 17174
rect 13813 17171 13879 17174
rect 15101 17234 15167 17237
rect 24025 17234 24091 17237
rect 15101 17232 24091 17234
rect 15101 17176 15106 17232
rect 15162 17176 24030 17232
rect 24086 17176 24091 17232
rect 15101 17174 24091 17176
rect 15101 17171 15167 17174
rect 24025 17171 24091 17174
rect 24301 17234 24367 17237
rect 26233 17234 26299 17237
rect 24301 17232 26299 17234
rect 24301 17176 24306 17232
rect 24362 17176 26238 17232
rect 26294 17176 26299 17232
rect 24301 17174 26299 17176
rect 24301 17171 24367 17174
rect 26233 17171 26299 17174
rect 1669 17098 1735 17101
rect 6085 17098 6151 17101
rect 1669 17096 6151 17098
rect 1669 17040 1674 17096
rect 1730 17040 6090 17096
rect 6146 17040 6151 17096
rect 1669 17038 6151 17040
rect 1669 17035 1735 17038
rect 6085 17035 6151 17038
rect 15009 17098 15075 17101
rect 15510 17098 15516 17100
rect 15009 17096 15516 17098
rect 15009 17040 15014 17096
rect 15070 17040 15516 17096
rect 15009 17038 15516 17040
rect 15009 17035 15075 17038
rect 15510 17036 15516 17038
rect 15580 17036 15586 17100
rect 16205 17098 16271 17101
rect 25221 17098 25287 17101
rect 16205 17096 25287 17098
rect 16205 17040 16210 17096
rect 16266 17040 25226 17096
rect 25282 17040 25287 17096
rect 16205 17038 25287 17040
rect 16205 17035 16271 17038
rect 25221 17035 25287 17038
rect 4337 16962 4403 16965
rect 7649 16962 7715 16965
rect 4337 16960 7715 16962
rect 4337 16904 4342 16960
rect 4398 16904 7654 16960
rect 7710 16904 7715 16960
rect 4337 16902 7715 16904
rect 4337 16899 4403 16902
rect 7649 16899 7715 16902
rect 10777 16962 10843 16965
rect 13077 16962 13143 16965
rect 10777 16960 13143 16962
rect 10777 16904 10782 16960
rect 10838 16904 13082 16960
rect 13138 16904 13143 16960
rect 10777 16902 13143 16904
rect 10777 16899 10843 16902
rect 13077 16899 13143 16902
rect 22461 16964 22527 16965
rect 22461 16960 22508 16964
rect 22572 16962 22578 16964
rect 22461 16904 22466 16960
rect 22461 16900 22508 16904
rect 22572 16902 22618 16962
rect 22572 16900 22578 16902
rect 23974 16900 23980 16964
rect 24044 16962 24050 16964
rect 24669 16962 24735 16965
rect 24044 16960 24735 16962
rect 24044 16904 24674 16960
rect 24730 16904 24735 16960
rect 24044 16902 24735 16904
rect 24044 16900 24050 16902
rect 22461 16899 22527 16900
rect 24669 16899 24735 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 3325 16826 3391 16829
rect 6453 16826 6519 16829
rect 3325 16824 6519 16826
rect 3325 16768 3330 16824
rect 3386 16768 6458 16824
rect 6514 16768 6519 16824
rect 3325 16766 6519 16768
rect 3325 16763 3391 16766
rect 6453 16763 6519 16766
rect 12985 16826 13051 16829
rect 16389 16826 16455 16829
rect 12985 16824 16455 16826
rect 12985 16768 12990 16824
rect 13046 16768 16394 16824
rect 16450 16768 16455 16824
rect 12985 16766 16455 16768
rect 12985 16763 13051 16766
rect 16389 16763 16455 16766
rect 23657 16826 23723 16829
rect 24301 16826 24367 16829
rect 23657 16824 24367 16826
rect 23657 16768 23662 16824
rect 23718 16768 24306 16824
rect 24362 16768 24367 16824
rect 23657 16766 24367 16768
rect 23657 16763 23723 16766
rect 24301 16763 24367 16766
rect 24669 16826 24735 16829
rect 24945 16826 25011 16829
rect 24669 16824 25011 16826
rect 24669 16768 24674 16824
rect 24730 16768 24950 16824
rect 25006 16768 25011 16824
rect 24669 16766 25011 16768
rect 24669 16763 24735 16766
rect 24945 16763 25011 16766
rect 0 16690 480 16720
rect 1577 16690 1643 16693
rect 0 16688 1643 16690
rect 0 16632 1582 16688
rect 1638 16632 1643 16688
rect 0 16630 1643 16632
rect 0 16600 480 16630
rect 1577 16627 1643 16630
rect 1853 16690 1919 16693
rect 6729 16690 6795 16693
rect 1853 16688 6795 16690
rect 1853 16632 1858 16688
rect 1914 16632 6734 16688
rect 6790 16632 6795 16688
rect 1853 16630 6795 16632
rect 1853 16627 1919 16630
rect 6729 16627 6795 16630
rect 8201 16690 8267 16693
rect 13537 16690 13603 16693
rect 18873 16690 18939 16693
rect 8201 16688 13603 16690
rect 8201 16632 8206 16688
rect 8262 16632 13542 16688
rect 13598 16632 13603 16688
rect 8201 16630 13603 16632
rect 8201 16627 8267 16630
rect 13537 16627 13603 16630
rect 13678 16688 18939 16690
rect 13678 16632 18878 16688
rect 18934 16632 18939 16688
rect 13678 16630 18939 16632
rect 6269 16554 6335 16557
rect 8569 16554 8635 16557
rect 13678 16554 13738 16630
rect 18873 16627 18939 16630
rect 19149 16690 19215 16693
rect 21541 16690 21607 16693
rect 19149 16688 21607 16690
rect 19149 16632 19154 16688
rect 19210 16632 21546 16688
rect 21602 16632 21607 16688
rect 19149 16630 21607 16632
rect 19149 16627 19215 16630
rect 21541 16627 21607 16630
rect 23381 16690 23447 16693
rect 27520 16690 28000 16720
rect 23381 16688 28000 16690
rect 23381 16632 23386 16688
rect 23442 16632 28000 16688
rect 23381 16630 28000 16632
rect 23381 16627 23447 16630
rect 27520 16600 28000 16630
rect 6269 16552 8635 16554
rect 6269 16496 6274 16552
rect 6330 16496 8574 16552
rect 8630 16496 8635 16552
rect 6269 16494 8635 16496
rect 6269 16491 6335 16494
rect 8569 16491 8635 16494
rect 12206 16494 13738 16554
rect 13813 16554 13879 16557
rect 14457 16554 14523 16557
rect 19057 16554 19123 16557
rect 24945 16554 25011 16557
rect 13813 16552 19123 16554
rect 13813 16496 13818 16552
rect 13874 16496 14462 16552
rect 14518 16496 19062 16552
rect 19118 16496 19123 16552
rect 13813 16494 19123 16496
rect 8201 16418 8267 16421
rect 9673 16418 9739 16421
rect 8201 16416 9739 16418
rect 8201 16360 8206 16416
rect 8262 16360 9678 16416
rect 9734 16360 9739 16416
rect 8201 16358 9739 16360
rect 8201 16355 8267 16358
rect 9673 16355 9739 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 2313 16282 2379 16285
rect 4613 16282 4679 16285
rect 12206 16282 12266 16494
rect 13813 16491 13879 16494
rect 14457 16491 14523 16494
rect 19057 16491 19123 16494
rect 24120 16552 25011 16554
rect 24120 16496 24950 16552
rect 25006 16496 25011 16552
rect 24120 16494 25011 16496
rect 24120 16418 24180 16494
rect 24945 16491 25011 16494
rect 24853 16420 24919 16421
rect 24853 16418 24900 16420
rect 19014 16358 24180 16418
rect 24808 16416 24900 16418
rect 24808 16360 24858 16416
rect 24808 16358 24900 16360
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 2313 16280 4679 16282
rect 2313 16224 2318 16280
rect 2374 16224 4618 16280
rect 4674 16224 4679 16280
rect 9768 16248 12266 16282
rect 2313 16222 4679 16224
rect 2313 16219 2379 16222
rect 4613 16219 4679 16222
rect 9492 16222 12266 16248
rect 15377 16282 15443 16285
rect 19014 16282 19074 16358
rect 24853 16356 24900 16358
rect 24964 16356 24970 16420
rect 24853 16355 24919 16356
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 15377 16280 19074 16282
rect 15377 16224 15382 16280
rect 15438 16224 19074 16280
rect 15377 16222 19074 16224
rect 21725 16282 21791 16285
rect 21725 16280 24042 16282
rect 21725 16224 21730 16280
rect 21786 16224 24042 16280
rect 21725 16222 24042 16224
rect 9492 16188 9828 16222
rect 15377 16219 15443 16222
rect 21725 16219 21791 16222
rect 0 16146 480 16176
rect 1393 16146 1459 16149
rect 0 16144 1459 16146
rect 0 16088 1398 16144
rect 1454 16088 1459 16144
rect 0 16086 1459 16088
rect 0 16056 480 16086
rect 1393 16083 1459 16086
rect 4061 16146 4127 16149
rect 6361 16146 6427 16149
rect 4061 16144 6427 16146
rect 4061 16088 4066 16144
rect 4122 16088 6366 16144
rect 6422 16088 6427 16144
rect 4061 16086 6427 16088
rect 4061 16083 4127 16086
rect 6361 16083 6427 16086
rect 6913 16146 6979 16149
rect 9492 16146 9552 16188
rect 6913 16144 9552 16146
rect 6913 16088 6918 16144
rect 6974 16088 9552 16144
rect 6913 16086 9552 16088
rect 10685 16146 10751 16149
rect 11145 16146 11211 16149
rect 10685 16144 11211 16146
rect 10685 16088 10690 16144
rect 10746 16088 11150 16144
rect 11206 16088 11211 16144
rect 10685 16086 11211 16088
rect 6913 16083 6979 16086
rect 10685 16083 10751 16086
rect 11145 16083 11211 16086
rect 11329 16146 11395 16149
rect 14549 16146 14615 16149
rect 17125 16146 17191 16149
rect 18781 16146 18847 16149
rect 11329 16144 14474 16146
rect 11329 16088 11334 16144
rect 11390 16088 14474 16144
rect 11329 16086 14474 16088
rect 11329 16083 11395 16086
rect 749 16010 815 16013
rect 14414 16010 14474 16086
rect 14549 16144 18847 16146
rect 14549 16088 14554 16144
rect 14610 16088 17130 16144
rect 17186 16088 18786 16144
rect 18842 16088 18847 16144
rect 14549 16086 18847 16088
rect 14549 16083 14615 16086
rect 17125 16083 17191 16086
rect 18781 16083 18847 16086
rect 19057 16146 19123 16149
rect 22461 16146 22527 16149
rect 22921 16148 22987 16149
rect 19057 16144 22527 16146
rect 19057 16088 19062 16144
rect 19118 16088 22466 16144
rect 22522 16088 22527 16144
rect 19057 16086 22527 16088
rect 19057 16083 19123 16086
rect 22461 16083 22527 16086
rect 22870 16084 22876 16148
rect 22940 16146 22987 16148
rect 23982 16146 24042 16222
rect 24761 16146 24827 16149
rect 27520 16146 28000 16176
rect 22940 16144 23032 16146
rect 22982 16088 23032 16144
rect 22940 16086 23032 16088
rect 23982 16144 24827 16146
rect 23982 16088 24766 16144
rect 24822 16088 24827 16144
rect 23982 16086 24827 16088
rect 22940 16084 22987 16086
rect 22921 16083 22987 16084
rect 24761 16083 24827 16086
rect 24902 16086 28000 16146
rect 17217 16010 17283 16013
rect 749 16008 14336 16010
rect 749 15952 754 16008
rect 810 15952 14336 16008
rect 749 15950 14336 15952
rect 14414 16008 17283 16010
rect 14414 15952 17222 16008
rect 17278 15952 17283 16008
rect 14414 15950 17283 15952
rect 749 15947 815 15950
rect 4153 15874 4219 15877
rect 7557 15874 7623 15877
rect 4153 15872 7623 15874
rect 4153 15816 4158 15872
rect 4214 15816 7562 15872
rect 7618 15816 7623 15872
rect 4153 15814 7623 15816
rect 14276 15874 14336 15950
rect 17217 15947 17283 15950
rect 17677 16010 17743 16013
rect 21817 16010 21883 16013
rect 17677 16008 21883 16010
rect 17677 15952 17682 16008
rect 17738 15952 21822 16008
rect 21878 15952 21883 16008
rect 17677 15950 21883 15952
rect 17677 15947 17743 15950
rect 21817 15947 21883 15950
rect 23841 16010 23907 16013
rect 24902 16010 24962 16086
rect 27520 16056 28000 16086
rect 23841 16008 24962 16010
rect 23841 15952 23846 16008
rect 23902 15952 24962 16008
rect 23841 15950 24962 15952
rect 23841 15947 23907 15950
rect 15745 15874 15811 15877
rect 14276 15872 15811 15874
rect 14276 15816 15750 15872
rect 15806 15816 15811 15872
rect 14276 15814 15811 15816
rect 17220 15874 17280 15947
rect 18781 15874 18847 15877
rect 17220 15872 18847 15874
rect 17220 15816 18786 15872
rect 18842 15816 18847 15872
rect 17220 15814 18847 15816
rect 4153 15811 4219 15814
rect 7557 15811 7623 15814
rect 15745 15811 15811 15814
rect 18781 15811 18847 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 4705 15738 4771 15741
rect 8385 15738 8451 15741
rect 10133 15738 10199 15741
rect 19241 15738 19307 15741
rect 20713 15738 20779 15741
rect 4705 15736 8451 15738
rect 4705 15680 4710 15736
rect 4766 15680 8390 15736
rect 8446 15680 8451 15736
rect 4705 15678 8451 15680
rect 4705 15675 4771 15678
rect 8385 15675 8451 15678
rect 8526 15736 10199 15738
rect 8526 15680 10138 15736
rect 10194 15680 10199 15736
rect 8526 15678 10199 15680
rect 4245 15602 4311 15605
rect 8526 15602 8586 15678
rect 10133 15675 10199 15678
rect 14414 15736 19307 15738
rect 14414 15680 19246 15736
rect 19302 15680 19307 15736
rect 14414 15678 19307 15680
rect 4245 15600 8586 15602
rect 4245 15544 4250 15600
rect 4306 15544 8586 15600
rect 4245 15542 8586 15544
rect 9121 15602 9187 15605
rect 14414 15602 14474 15678
rect 19241 15675 19307 15678
rect 20670 15736 20779 15738
rect 20670 15680 20718 15736
rect 20774 15680 20779 15736
rect 20670 15675 20779 15680
rect 23105 15738 23171 15741
rect 23289 15738 23355 15741
rect 23105 15736 23355 15738
rect 23105 15680 23110 15736
rect 23166 15680 23294 15736
rect 23350 15680 23355 15736
rect 23105 15678 23355 15680
rect 23105 15675 23171 15678
rect 23289 15675 23355 15678
rect 9121 15600 14474 15602
rect 9121 15544 9126 15600
rect 9182 15544 14474 15600
rect 9121 15542 14474 15544
rect 14549 15602 14615 15605
rect 20670 15602 20730 15675
rect 25221 15602 25287 15605
rect 14549 15600 25287 15602
rect 14549 15544 14554 15600
rect 14610 15544 25226 15600
rect 25282 15544 25287 15600
rect 14549 15542 25287 15544
rect 4245 15539 4311 15542
rect 9121 15539 9187 15542
rect 14549 15539 14615 15542
rect 25221 15539 25287 15542
rect 0 15466 480 15496
rect 3509 15466 3575 15469
rect 0 15464 3575 15466
rect 0 15408 3514 15464
rect 3570 15408 3575 15464
rect 0 15406 3575 15408
rect 0 15376 480 15406
rect 3509 15403 3575 15406
rect 3877 15466 3943 15469
rect 5533 15466 5599 15469
rect 3877 15464 5599 15466
rect 3877 15408 3882 15464
rect 3938 15408 5538 15464
rect 5594 15408 5599 15464
rect 3877 15406 5599 15408
rect 3877 15403 3943 15406
rect 5533 15403 5599 15406
rect 10317 15466 10383 15469
rect 15561 15466 15627 15469
rect 10317 15464 15627 15466
rect 10317 15408 10322 15464
rect 10378 15408 15566 15464
rect 15622 15408 15627 15464
rect 10317 15406 15627 15408
rect 10317 15403 10383 15406
rect 15561 15403 15627 15406
rect 15745 15466 15811 15469
rect 17217 15466 17283 15469
rect 15745 15464 17283 15466
rect 15745 15408 15750 15464
rect 15806 15408 17222 15464
rect 17278 15408 17283 15464
rect 15745 15406 17283 15408
rect 15745 15403 15811 15406
rect 17217 15403 17283 15406
rect 24761 15466 24827 15469
rect 25037 15466 25103 15469
rect 27520 15466 28000 15496
rect 24761 15464 28000 15466
rect 24761 15408 24766 15464
rect 24822 15408 25042 15464
rect 25098 15408 28000 15464
rect 24761 15406 28000 15408
rect 24761 15403 24827 15406
rect 25037 15403 25103 15406
rect 27520 15376 28000 15406
rect 6177 15330 6243 15333
rect 6545 15330 6611 15333
rect 6177 15328 6611 15330
rect 6177 15272 6182 15328
rect 6238 15272 6550 15328
rect 6606 15272 6611 15328
rect 6177 15270 6611 15272
rect 6177 15267 6243 15270
rect 6545 15267 6611 15270
rect 9765 15330 9831 15333
rect 12617 15330 12683 15333
rect 9765 15328 12683 15330
rect 9765 15272 9770 15328
rect 9826 15272 12622 15328
rect 12678 15272 12683 15328
rect 9765 15270 12683 15272
rect 9765 15267 9831 15270
rect 12617 15267 12683 15270
rect 17769 15330 17835 15333
rect 23749 15330 23815 15333
rect 17769 15328 23815 15330
rect 17769 15272 17774 15328
rect 17830 15272 23754 15328
rect 23810 15272 23815 15328
rect 17769 15270 23815 15272
rect 17769 15267 17835 15270
rect 23749 15267 23815 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 1669 15194 1735 15197
rect 5165 15194 5231 15197
rect 1669 15192 5231 15194
rect 1669 15136 1674 15192
rect 1730 15136 5170 15192
rect 5226 15136 5231 15192
rect 1669 15134 5231 15136
rect 1669 15131 1735 15134
rect 5165 15131 5231 15134
rect 8017 15194 8083 15197
rect 12893 15194 12959 15197
rect 8017 15192 12959 15194
rect 8017 15136 8022 15192
rect 8078 15136 12898 15192
rect 12954 15136 12959 15192
rect 8017 15134 12959 15136
rect 8017 15131 8083 15134
rect 12893 15131 12959 15134
rect 17033 15194 17099 15197
rect 23381 15194 23447 15197
rect 17033 15192 23447 15194
rect 17033 15136 17038 15192
rect 17094 15136 23386 15192
rect 23442 15136 23447 15192
rect 17033 15134 23447 15136
rect 17033 15131 17099 15134
rect 23381 15131 23447 15134
rect 4521 15058 4587 15061
rect 6269 15058 6335 15061
rect 4521 15056 6335 15058
rect 4521 15000 4526 15056
rect 4582 15000 6274 15056
rect 6330 15000 6335 15056
rect 4521 14998 6335 15000
rect 4521 14995 4587 14998
rect 6269 14995 6335 14998
rect 7373 15058 7439 15061
rect 18689 15058 18755 15061
rect 18965 15058 19031 15061
rect 7373 15056 19031 15058
rect 7373 15000 7378 15056
rect 7434 15000 18694 15056
rect 18750 15000 18970 15056
rect 19026 15000 19031 15056
rect 7373 14998 19031 15000
rect 7373 14995 7439 14998
rect 18689 14995 18755 14998
rect 18965 14995 19031 14998
rect 22686 14996 22692 15060
rect 22756 15058 22762 15060
rect 22756 14998 23674 15058
rect 22756 14996 22762 14998
rect 0 14922 480 14952
rect 3785 14922 3851 14925
rect 0 14920 3851 14922
rect 0 14864 3790 14920
rect 3846 14864 3851 14920
rect 0 14862 3851 14864
rect 0 14832 480 14862
rect 3785 14859 3851 14862
rect 11697 14922 11763 14925
rect 23473 14922 23539 14925
rect 11697 14920 23539 14922
rect 11697 14864 11702 14920
rect 11758 14864 23478 14920
rect 23534 14864 23539 14920
rect 11697 14862 23539 14864
rect 23614 14922 23674 14998
rect 27520 14922 28000 14952
rect 23614 14862 28000 14922
rect 11697 14859 11763 14862
rect 23473 14859 23539 14862
rect 27520 14832 28000 14862
rect 3877 14786 3943 14789
rect 5257 14786 5323 14789
rect 5625 14786 5691 14789
rect 3877 14784 5691 14786
rect 3877 14728 3882 14784
rect 3938 14728 5262 14784
rect 5318 14728 5630 14784
rect 5686 14728 5691 14784
rect 3877 14726 5691 14728
rect 3877 14723 3943 14726
rect 5257 14723 5323 14726
rect 5625 14723 5691 14726
rect 10961 14786 11027 14789
rect 12801 14786 12867 14789
rect 10961 14784 12867 14786
rect 10961 14728 10966 14784
rect 11022 14728 12806 14784
rect 12862 14728 12867 14784
rect 10961 14726 12867 14728
rect 10961 14723 11027 14726
rect 12801 14723 12867 14726
rect 22001 14786 22067 14789
rect 22921 14786 22987 14789
rect 22001 14784 22987 14786
rect 22001 14728 22006 14784
rect 22062 14728 22926 14784
rect 22982 14728 22987 14784
rect 22001 14726 22987 14728
rect 22001 14723 22067 14726
rect 22921 14723 22987 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 2773 14650 2839 14653
rect 3325 14650 3391 14653
rect 4429 14650 4495 14653
rect 2773 14648 4495 14650
rect 2773 14592 2778 14648
rect 2834 14592 3330 14648
rect 3386 14592 4434 14648
rect 4490 14592 4495 14648
rect 2773 14590 4495 14592
rect 2773 14587 2839 14590
rect 3325 14587 3391 14590
rect 4429 14587 4495 14590
rect 5349 14650 5415 14653
rect 6637 14650 6703 14653
rect 5349 14648 6703 14650
rect 5349 14592 5354 14648
rect 5410 14592 6642 14648
rect 6698 14592 6703 14648
rect 5349 14590 6703 14592
rect 5349 14587 5415 14590
rect 6637 14587 6703 14590
rect 15285 14650 15351 14653
rect 17769 14650 17835 14653
rect 22185 14652 22251 14653
rect 22134 14650 22140 14652
rect 15285 14648 17835 14650
rect 15285 14592 15290 14648
rect 15346 14592 17774 14648
rect 17830 14592 17835 14648
rect 15285 14590 17835 14592
rect 22094 14590 22140 14650
rect 22204 14648 22251 14652
rect 22246 14592 22251 14648
rect 15285 14587 15351 14590
rect 17769 14587 17835 14590
rect 22134 14588 22140 14590
rect 22204 14588 22251 14592
rect 22502 14588 22508 14652
rect 22572 14650 22578 14652
rect 22645 14650 22711 14653
rect 22572 14648 22711 14650
rect 22572 14592 22650 14648
rect 22706 14592 22711 14648
rect 22572 14590 22711 14592
rect 22572 14588 22578 14590
rect 22185 14587 22251 14588
rect 22645 14587 22711 14590
rect 22870 14588 22876 14652
rect 22940 14650 22946 14652
rect 22940 14590 24226 14650
rect 22940 14588 22946 14590
rect 10041 14514 10107 14517
rect 16665 14514 16731 14517
rect 10041 14512 16731 14514
rect 10041 14456 10046 14512
rect 10102 14456 16670 14512
rect 16726 14456 16731 14512
rect 10041 14454 16731 14456
rect 10041 14451 10107 14454
rect 16665 14451 16731 14454
rect 19374 14452 19380 14516
rect 19444 14514 19450 14516
rect 24025 14514 24091 14517
rect 19444 14512 24091 14514
rect 19444 14456 24030 14512
rect 24086 14456 24091 14512
rect 19444 14454 24091 14456
rect 19444 14452 19450 14454
rect 24025 14451 24091 14454
rect 0 14378 480 14408
rect 3233 14378 3299 14381
rect 0 14376 3299 14378
rect 0 14320 3238 14376
rect 3294 14320 3299 14376
rect 0 14318 3299 14320
rect 0 14288 480 14318
rect 3233 14315 3299 14318
rect 5165 14378 5231 14381
rect 6453 14378 6519 14381
rect 7465 14378 7531 14381
rect 5165 14376 7531 14378
rect 5165 14320 5170 14376
rect 5226 14320 6458 14376
rect 6514 14320 7470 14376
rect 7526 14320 7531 14376
rect 5165 14318 7531 14320
rect 5165 14315 5231 14318
rect 6453 14315 6519 14318
rect 7465 14315 7531 14318
rect 16297 14378 16363 14381
rect 19977 14378 20043 14381
rect 16297 14376 20043 14378
rect 16297 14320 16302 14376
rect 16358 14320 19982 14376
rect 20038 14320 20043 14376
rect 16297 14318 20043 14320
rect 16297 14315 16363 14318
rect 19977 14315 20043 14318
rect 20253 14378 20319 14381
rect 23974 14378 23980 14380
rect 20253 14376 23980 14378
rect 20253 14320 20258 14376
rect 20314 14320 23980 14376
rect 20253 14318 23980 14320
rect 20253 14315 20319 14318
rect 23974 14316 23980 14318
rect 24044 14316 24050 14380
rect 24166 14378 24226 14590
rect 27520 14378 28000 14408
rect 24166 14318 28000 14378
rect 27520 14288 28000 14318
rect 21449 14242 21515 14245
rect 23657 14242 23723 14245
rect 21449 14240 23723 14242
rect 21449 14184 21454 14240
rect 21510 14184 23662 14240
rect 23718 14184 23723 14240
rect 21449 14182 23723 14184
rect 21449 14179 21515 14182
rect 23657 14179 23723 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 11973 14106 12039 14109
rect 13997 14106 14063 14109
rect 11973 14104 14063 14106
rect 11973 14048 11978 14104
rect 12034 14048 14002 14104
rect 14058 14048 14063 14104
rect 11973 14046 14063 14048
rect 11973 14043 12039 14046
rect 13997 14043 14063 14046
rect 12433 13970 12499 13973
rect 24209 13970 24275 13973
rect 24853 13970 24919 13973
rect 12433 13968 24919 13970
rect 12433 13912 12438 13968
rect 12494 13912 24214 13968
rect 24270 13912 24858 13968
rect 24914 13912 24919 13968
rect 12433 13910 24919 13912
rect 12433 13907 12499 13910
rect 24209 13907 24275 13910
rect 24853 13907 24919 13910
rect 9121 13834 9187 13837
rect 12157 13834 12223 13837
rect 9121 13832 12223 13834
rect 9121 13776 9126 13832
rect 9182 13776 12162 13832
rect 12218 13776 12223 13832
rect 9121 13774 12223 13776
rect 9121 13771 9187 13774
rect 12157 13771 12223 13774
rect 21817 13834 21883 13837
rect 25405 13834 25471 13837
rect 21817 13832 25471 13834
rect 21817 13776 21822 13832
rect 21878 13776 25410 13832
rect 25466 13776 25471 13832
rect 21817 13774 25471 13776
rect 21817 13771 21883 13774
rect 25405 13771 25471 13774
rect 0 13698 480 13728
rect 3417 13698 3483 13701
rect 0 13696 3483 13698
rect 0 13640 3422 13696
rect 3478 13640 3483 13696
rect 0 13638 3483 13640
rect 0 13608 480 13638
rect 3417 13635 3483 13638
rect 11881 13698 11947 13701
rect 12985 13698 13051 13701
rect 13813 13698 13879 13701
rect 11881 13696 13879 13698
rect 11881 13640 11886 13696
rect 11942 13640 12990 13696
rect 13046 13640 13818 13696
rect 13874 13640 13879 13696
rect 11881 13638 13879 13640
rect 11881 13635 11947 13638
rect 12985 13635 13051 13638
rect 13813 13635 13879 13638
rect 16849 13698 16915 13701
rect 19425 13698 19491 13701
rect 16849 13696 19491 13698
rect 16849 13640 16854 13696
rect 16910 13640 19430 13696
rect 19486 13640 19491 13696
rect 16849 13638 19491 13640
rect 16849 13635 16915 13638
rect 19425 13635 19491 13638
rect 20437 13698 20503 13701
rect 27520 13698 28000 13728
rect 20437 13696 28000 13698
rect 20437 13640 20442 13696
rect 20498 13640 28000 13696
rect 20437 13638 28000 13640
rect 20437 13635 20503 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 27520 13608 28000 13638
rect 19610 13567 19930 13568
rect 10685 13562 10751 13565
rect 13353 13562 13419 13565
rect 10685 13560 13419 13562
rect 10685 13504 10690 13560
rect 10746 13504 13358 13560
rect 13414 13504 13419 13560
rect 10685 13502 13419 13504
rect 10685 13499 10751 13502
rect 13353 13499 13419 13502
rect 14273 13562 14339 13565
rect 17861 13562 17927 13565
rect 14273 13560 17927 13562
rect 14273 13504 14278 13560
rect 14334 13504 17866 13560
rect 17922 13504 17927 13560
rect 14273 13502 17927 13504
rect 14273 13499 14339 13502
rect 17861 13499 17927 13502
rect 21633 13562 21699 13565
rect 22369 13562 22435 13565
rect 21633 13560 22435 13562
rect 21633 13504 21638 13560
rect 21694 13504 22374 13560
rect 22430 13504 22435 13560
rect 21633 13502 22435 13504
rect 21633 13499 21699 13502
rect 22369 13499 22435 13502
rect 22553 13562 22619 13565
rect 25865 13562 25931 13565
rect 22553 13560 25931 13562
rect 22553 13504 22558 13560
rect 22614 13504 25870 13560
rect 25926 13504 25931 13560
rect 22553 13502 25931 13504
rect 22553 13499 22619 13502
rect 25865 13499 25931 13502
rect 6361 13426 6427 13429
rect 24209 13426 24275 13429
rect 6361 13424 24275 13426
rect 6361 13368 6366 13424
rect 6422 13368 24214 13424
rect 24270 13368 24275 13424
rect 6361 13366 24275 13368
rect 6361 13363 6427 13366
rect 24209 13363 24275 13366
rect 2773 13290 2839 13293
rect 3877 13290 3943 13293
rect 2773 13288 3943 13290
rect 2773 13232 2778 13288
rect 2834 13232 3882 13288
rect 3938 13232 3943 13288
rect 2773 13230 3943 13232
rect 2773 13227 2839 13230
rect 3877 13227 3943 13230
rect 6177 13290 6243 13293
rect 8569 13290 8635 13293
rect 13813 13290 13879 13293
rect 17493 13290 17559 13293
rect 20805 13290 20871 13293
rect 6177 13288 17418 13290
rect 6177 13232 6182 13288
rect 6238 13232 8574 13288
rect 8630 13232 13818 13288
rect 13874 13232 17418 13288
rect 6177 13230 17418 13232
rect 6177 13227 6243 13230
rect 8569 13227 8635 13230
rect 13813 13227 13879 13230
rect 0 13154 480 13184
rect 3417 13154 3483 13157
rect 0 13152 3483 13154
rect 0 13096 3422 13152
rect 3478 13096 3483 13152
rect 0 13094 3483 13096
rect 17358 13154 17418 13230
rect 17493 13288 20871 13290
rect 17493 13232 17498 13288
rect 17554 13232 20810 13288
rect 20866 13232 20871 13288
rect 17493 13230 20871 13232
rect 17493 13227 17559 13230
rect 20805 13227 20871 13230
rect 22369 13290 22435 13293
rect 23606 13290 23612 13292
rect 22369 13288 23612 13290
rect 22369 13232 22374 13288
rect 22430 13232 23612 13288
rect 22369 13230 23612 13232
rect 22369 13227 22435 13230
rect 23606 13228 23612 13230
rect 23676 13228 23682 13292
rect 18045 13154 18111 13157
rect 17358 13152 18111 13154
rect 17358 13096 18050 13152
rect 18106 13096 18111 13152
rect 17358 13094 18111 13096
rect 0 13064 480 13094
rect 3417 13091 3483 13094
rect 18045 13091 18111 13094
rect 18505 13154 18571 13157
rect 26233 13154 26299 13157
rect 27520 13154 28000 13184
rect 18505 13152 24042 13154
rect 18505 13096 18510 13152
rect 18566 13096 24042 13152
rect 18505 13094 24042 13096
rect 18505 13091 18571 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 7189 13018 7255 13021
rect 9949 13018 10015 13021
rect 7189 13016 10015 13018
rect 7189 12960 7194 13016
rect 7250 12960 9954 13016
rect 10010 12960 10015 13016
rect 7189 12958 10015 12960
rect 7189 12955 7255 12958
rect 9949 12955 10015 12958
rect 16757 13018 16823 13021
rect 19374 13018 19380 13020
rect 16757 13016 19380 13018
rect 16757 12960 16762 13016
rect 16818 12960 19380 13016
rect 16757 12958 19380 12960
rect 16757 12955 16823 12958
rect 19374 12956 19380 12958
rect 19444 12956 19450 13020
rect 22645 13018 22711 13021
rect 23422 13018 23428 13020
rect 22645 13016 23428 13018
rect 22645 12960 22650 13016
rect 22706 12960 23428 13016
rect 22645 12958 23428 12960
rect 22645 12955 22711 12958
rect 23422 12956 23428 12958
rect 23492 12956 23498 13020
rect 4705 12882 4771 12885
rect 5165 12882 5231 12885
rect 7925 12882 7991 12885
rect 4705 12880 7991 12882
rect 4705 12824 4710 12880
rect 4766 12824 5170 12880
rect 5226 12824 7930 12880
rect 7986 12824 7991 12880
rect 4705 12822 7991 12824
rect 4705 12819 4771 12822
rect 5165 12819 5231 12822
rect 7925 12819 7991 12822
rect 13261 12882 13327 12885
rect 23790 12882 23796 12884
rect 13261 12880 23796 12882
rect 13261 12824 13266 12880
rect 13322 12824 23796 12880
rect 13261 12822 23796 12824
rect 13261 12819 13327 12822
rect 23790 12820 23796 12822
rect 23860 12820 23866 12884
rect 3509 12746 3575 12749
rect 21909 12746 21975 12749
rect 3509 12744 21975 12746
rect 3509 12688 3514 12744
rect 3570 12688 21914 12744
rect 21970 12688 21975 12744
rect 3509 12686 21975 12688
rect 3509 12683 3575 12686
rect 21909 12683 21975 12686
rect 23606 12684 23612 12748
rect 23676 12746 23682 12748
rect 23749 12746 23815 12749
rect 23676 12744 23815 12746
rect 23676 12688 23754 12744
rect 23810 12688 23815 12744
rect 23676 12686 23815 12688
rect 23982 12746 24042 13094
rect 26233 13152 28000 13154
rect 26233 13096 26238 13152
rect 26294 13096 28000 13152
rect 26233 13094 28000 13096
rect 26233 13091 26299 13094
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13094
rect 24277 13023 24597 13024
rect 24117 12882 24183 12885
rect 24710 12882 24716 12884
rect 24117 12880 24716 12882
rect 24117 12824 24122 12880
rect 24178 12824 24716 12880
rect 24117 12822 24716 12824
rect 24117 12819 24183 12822
rect 24710 12820 24716 12822
rect 24780 12820 24786 12884
rect 23982 12686 25514 12746
rect 23676 12684 23682 12686
rect 23749 12683 23815 12686
rect 14089 12610 14155 12613
rect 18689 12610 18755 12613
rect 14089 12608 18755 12610
rect 14089 12552 14094 12608
rect 14150 12552 18694 12608
rect 18750 12552 18755 12608
rect 14089 12550 18755 12552
rect 14089 12547 14155 12550
rect 18689 12547 18755 12550
rect 20621 12610 20687 12613
rect 25313 12610 25379 12613
rect 20621 12608 25379 12610
rect 20621 12552 20626 12608
rect 20682 12552 25318 12608
rect 25374 12552 25379 12608
rect 20621 12550 25379 12552
rect 20621 12547 20687 12550
rect 25313 12547 25379 12550
rect 10277 12544 10597 12545
rect 0 12474 480 12504
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 6913 12474 6979 12477
rect 0 12472 6979 12474
rect 0 12416 6918 12472
rect 6974 12416 6979 12472
rect 0 12414 6979 12416
rect 0 12384 480 12414
rect 6913 12411 6979 12414
rect 11513 12474 11579 12477
rect 14825 12474 14891 12477
rect 11513 12472 14891 12474
rect 11513 12416 11518 12472
rect 11574 12416 14830 12472
rect 14886 12416 14891 12472
rect 11513 12414 14891 12416
rect 11513 12411 11579 12414
rect 14825 12411 14891 12414
rect 21081 12474 21147 12477
rect 23381 12474 23447 12477
rect 21081 12472 23447 12474
rect 21081 12416 21086 12472
rect 21142 12416 23386 12472
rect 23442 12416 23447 12472
rect 21081 12414 23447 12416
rect 21081 12411 21147 12414
rect 23381 12411 23447 12414
rect 23790 12412 23796 12476
rect 23860 12474 23866 12476
rect 24393 12474 24459 12477
rect 25129 12474 25195 12477
rect 23860 12472 25195 12474
rect 23860 12416 24398 12472
rect 24454 12416 25134 12472
rect 25190 12416 25195 12472
rect 23860 12414 25195 12416
rect 25454 12474 25514 12686
rect 27520 12474 28000 12504
rect 25454 12414 28000 12474
rect 23860 12412 23866 12414
rect 24393 12411 24459 12414
rect 25129 12411 25195 12414
rect 27520 12384 28000 12414
rect 4705 12338 4771 12341
rect 8477 12338 8543 12341
rect 4705 12336 8543 12338
rect 4705 12280 4710 12336
rect 4766 12280 8482 12336
rect 8538 12280 8543 12336
rect 4705 12278 8543 12280
rect 4705 12275 4771 12278
rect 8477 12275 8543 12278
rect 10133 12338 10199 12341
rect 16205 12338 16271 12341
rect 10133 12336 25882 12338
rect 10133 12280 10138 12336
rect 10194 12280 16210 12336
rect 16266 12280 25882 12336
rect 10133 12278 25882 12280
rect 10133 12275 10199 12278
rect 16205 12275 16271 12278
rect 3417 12202 3483 12205
rect 19793 12202 19859 12205
rect 25681 12202 25747 12205
rect 3417 12200 12220 12202
rect 3417 12144 3422 12200
rect 3478 12168 12220 12200
rect 12344 12168 15394 12202
rect 3478 12144 15394 12168
rect 3417 12142 15394 12144
rect 3417 12139 3483 12142
rect 12160 12108 12404 12142
rect 12985 12066 13051 12069
rect 13169 12066 13235 12069
rect 15334 12066 15394 12142
rect 19793 12200 25747 12202
rect 19793 12144 19798 12200
rect 19854 12144 25686 12200
rect 25742 12144 25747 12200
rect 19793 12142 25747 12144
rect 19793 12139 19859 12142
rect 25681 12139 25747 12142
rect 20621 12066 20687 12069
rect 12985 12064 14842 12066
rect 12985 12008 12990 12064
rect 13046 12008 13174 12064
rect 13230 12008 14842 12064
rect 12985 12006 14842 12008
rect 15334 12064 20687 12066
rect 15334 12008 20626 12064
rect 20682 12008 20687 12064
rect 15334 12006 20687 12008
rect 12985 12003 13051 12006
rect 13169 12003 13235 12006
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 4061 11930 4127 11933
rect 0 11928 4127 11930
rect 0 11872 4066 11928
rect 4122 11872 4127 11928
rect 0 11870 4127 11872
rect 0 11840 480 11870
rect 4061 11867 4127 11870
rect 9213 11930 9279 11933
rect 10685 11930 10751 11933
rect 9213 11928 10751 11930
rect 9213 11872 9218 11928
rect 9274 11872 10690 11928
rect 10746 11872 10751 11928
rect 9213 11870 10751 11872
rect 9213 11867 9279 11870
rect 10685 11867 10751 11870
rect 7557 11794 7623 11797
rect 14782 11794 14842 12006
rect 20621 12003 20687 12006
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 23013 11930 23079 11933
rect 15334 11928 23079 11930
rect 15334 11872 23018 11928
rect 23074 11872 23079 11928
rect 15334 11870 23079 11872
rect 25822 11930 25882 12278
rect 27520 11930 28000 11960
rect 25822 11870 28000 11930
rect 15334 11794 15394 11870
rect 23013 11867 23079 11870
rect 27520 11840 28000 11870
rect 7557 11792 14658 11794
rect 7557 11736 7562 11792
rect 7618 11736 14658 11792
rect 7557 11734 14658 11736
rect 14782 11734 15394 11794
rect 17861 11794 17927 11797
rect 22277 11794 22343 11797
rect 17861 11792 22343 11794
rect 17861 11736 17866 11792
rect 17922 11736 22282 11792
rect 22338 11736 22343 11792
rect 17861 11734 22343 11736
rect 7557 11731 7623 11734
rect 13721 11658 13787 11661
rect 2868 11656 13787 11658
rect 2868 11600 13726 11656
rect 13782 11600 13787 11656
rect 2868 11598 13787 11600
rect 14598 11658 14658 11734
rect 17861 11731 17927 11734
rect 22277 11731 22343 11734
rect 14733 11658 14799 11661
rect 15745 11658 15811 11661
rect 22369 11658 22435 11661
rect 14598 11656 14799 11658
rect 14598 11600 14738 11656
rect 14794 11600 14799 11656
rect 14598 11598 14799 11600
rect 0 11250 480 11280
rect 2868 11250 2928 11598
rect 13721 11595 13787 11598
rect 14733 11595 14799 11598
rect 14966 11656 22435 11658
rect 14966 11600 15750 11656
rect 15806 11600 22374 11656
rect 22430 11600 22435 11656
rect 14966 11598 22435 11600
rect 4613 11522 4679 11525
rect 10133 11522 10199 11525
rect 4613 11520 10199 11522
rect 4613 11464 4618 11520
rect 4674 11464 10138 11520
rect 10194 11464 10199 11520
rect 4613 11462 10199 11464
rect 4613 11459 4679 11462
rect 10133 11459 10199 11462
rect 13077 11522 13143 11525
rect 14966 11522 15026 11598
rect 15745 11595 15811 11598
rect 22369 11595 22435 11598
rect 13077 11520 15026 11522
rect 13077 11464 13082 11520
rect 13138 11464 15026 11520
rect 13077 11462 15026 11464
rect 13077 11459 13143 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 10685 11386 10751 11389
rect 24577 11386 24643 11389
rect 10685 11384 17234 11386
rect 10685 11328 10690 11384
rect 10746 11328 17234 11384
rect 10685 11326 17234 11328
rect 10685 11323 10751 11326
rect 0 11190 2928 11250
rect 4061 11250 4127 11253
rect 12801 11250 12867 11253
rect 4061 11248 12867 11250
rect 4061 11192 4066 11248
rect 4122 11192 12806 11248
rect 12862 11192 12867 11248
rect 4061 11190 12867 11192
rect 17174 11250 17234 11326
rect 23430 11384 24643 11386
rect 23430 11328 24582 11384
rect 24638 11328 24643 11384
rect 23430 11326 24643 11328
rect 23430 11250 23490 11326
rect 24577 11323 24643 11326
rect 23657 11252 23723 11253
rect 23606 11250 23612 11252
rect 17174 11190 23490 11250
rect 23566 11190 23612 11250
rect 23676 11248 23723 11252
rect 27520 11250 28000 11280
rect 23718 11192 23723 11248
rect 0 11160 480 11190
rect 4061 11187 4127 11190
rect 12801 11187 12867 11190
rect 23606 11188 23612 11190
rect 23676 11188 23723 11192
rect 23657 11187 23723 11188
rect 24902 11190 28000 11250
rect 3877 11114 3943 11117
rect 13077 11114 13143 11117
rect 3877 11112 13143 11114
rect 3877 11056 3882 11112
rect 3938 11056 13082 11112
rect 13138 11056 13143 11112
rect 3877 11054 13143 11056
rect 3877 11051 3943 11054
rect 13077 11051 13143 11054
rect 14273 11114 14339 11117
rect 16849 11114 16915 11117
rect 14273 11112 16915 11114
rect 14273 11056 14278 11112
rect 14334 11056 16854 11112
rect 16910 11056 16915 11112
rect 14273 11054 16915 11056
rect 14273 11051 14339 11054
rect 16849 11051 16915 11054
rect 18965 11114 19031 11117
rect 24902 11114 24962 11190
rect 27520 11160 28000 11190
rect 18965 11112 24962 11114
rect 18965 11056 18970 11112
rect 19026 11056 24962 11112
rect 18965 11054 24962 11056
rect 18965 11051 19031 11054
rect 17125 10978 17191 10981
rect 23473 10978 23539 10981
rect 17125 10976 23539 10978
rect 17125 10920 17130 10976
rect 17186 10920 23478 10976
rect 23534 10920 23539 10976
rect 17125 10918 23539 10920
rect 17125 10915 17191 10918
rect 23473 10915 23539 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 0 10706 480 10736
rect 1393 10706 1459 10709
rect 0 10704 1459 10706
rect 0 10648 1398 10704
rect 1454 10648 1459 10704
rect 0 10646 1459 10648
rect 0 10616 480 10646
rect 1393 10643 1459 10646
rect 9489 10706 9555 10709
rect 24393 10706 24459 10709
rect 27520 10706 28000 10736
rect 9489 10704 24459 10706
rect 9489 10648 9494 10704
rect 9550 10648 24398 10704
rect 24454 10648 24459 10704
rect 9489 10646 24459 10648
rect 9489 10643 9555 10646
rect 24393 10643 24459 10646
rect 24534 10646 28000 10706
rect 1577 10570 1643 10573
rect 23565 10570 23631 10573
rect 24534 10570 24594 10646
rect 27520 10616 28000 10646
rect 1577 10568 20178 10570
rect 1577 10512 1582 10568
rect 1638 10512 20178 10568
rect 1577 10510 20178 10512
rect 1577 10507 1643 10510
rect 20118 10434 20178 10510
rect 23565 10568 24594 10570
rect 23565 10512 23570 10568
rect 23626 10512 24594 10568
rect 23565 10510 24594 10512
rect 23565 10507 23631 10510
rect 26141 10434 26207 10437
rect 20118 10432 26207 10434
rect 20118 10376 26146 10432
rect 26202 10376 26207 10432
rect 20118 10374 26207 10376
rect 26141 10371 26207 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 13445 10162 13511 10165
rect 22461 10162 22527 10165
rect 23933 10162 23999 10165
rect 13445 10160 23999 10162
rect 13445 10104 13450 10160
rect 13506 10104 22466 10160
rect 22522 10104 23938 10160
rect 23994 10104 23999 10160
rect 13445 10102 23999 10104
rect 13445 10099 13511 10102
rect 22461 10099 22527 10102
rect 23933 10099 23999 10102
rect 24761 10162 24827 10165
rect 24894 10162 24900 10164
rect 24761 10160 24900 10162
rect 24761 10104 24766 10160
rect 24822 10104 24900 10160
rect 24761 10102 24900 10104
rect 24761 10099 24827 10102
rect 24894 10100 24900 10102
rect 24964 10100 24970 10164
rect 0 10026 480 10056
rect 9213 10026 9279 10029
rect 0 10024 9279 10026
rect 0 9968 9218 10024
rect 9274 9968 9279 10024
rect 0 9966 9279 9968
rect 0 9936 480 9966
rect 9213 9963 9279 9966
rect 20897 10026 20963 10029
rect 27520 10026 28000 10056
rect 20897 10024 28000 10026
rect 20897 9968 20902 10024
rect 20958 9968 28000 10024
rect 20897 9966 28000 9968
rect 20897 9963 20963 9966
rect 27520 9936 28000 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 4061 9618 4127 9621
rect 12985 9618 13051 9621
rect 4061 9616 13051 9618
rect 4061 9560 4066 9616
rect 4122 9560 12990 9616
rect 13046 9560 13051 9616
rect 4061 9558 13051 9560
rect 4061 9555 4127 9558
rect 12985 9555 13051 9558
rect 14549 9618 14615 9621
rect 23841 9618 23907 9621
rect 14549 9616 23907 9618
rect 14549 9560 14554 9616
rect 14610 9560 23846 9616
rect 23902 9560 23907 9616
rect 14549 9558 23907 9560
rect 14549 9555 14615 9558
rect 23841 9555 23907 9558
rect 0 9482 480 9512
rect 11697 9482 11763 9485
rect 0 9480 11763 9482
rect 0 9424 11702 9480
rect 11758 9424 11763 9480
rect 0 9422 11763 9424
rect 0 9392 480 9422
rect 11697 9419 11763 9422
rect 17953 9482 18019 9485
rect 18597 9482 18663 9485
rect 24669 9482 24735 9485
rect 25129 9482 25195 9485
rect 27520 9482 28000 9512
rect 17953 9480 25195 9482
rect 17953 9424 17958 9480
rect 18014 9424 18602 9480
rect 18658 9424 24674 9480
rect 24730 9424 25134 9480
rect 25190 9424 25195 9480
rect 17953 9422 25195 9424
rect 17953 9419 18019 9422
rect 18597 9419 18663 9422
rect 24669 9419 24735 9422
rect 25129 9419 25195 9422
rect 25270 9422 28000 9482
rect 22921 9346 22987 9349
rect 25270 9346 25330 9422
rect 27520 9392 28000 9422
rect 22921 9344 25330 9346
rect 22921 9288 22926 9344
rect 22982 9288 25330 9344
rect 22921 9286 25330 9288
rect 22921 9283 22987 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 12206 9150 14474 9210
rect 9581 9074 9647 9077
rect 12206 9074 12266 9150
rect 9581 9072 12266 9074
rect 9581 9016 9586 9072
rect 9642 9016 12266 9072
rect 9581 9014 12266 9016
rect 9581 9011 9647 9014
rect 14414 8938 14474 9150
rect 14733 9074 14799 9077
rect 20989 9074 21055 9077
rect 14733 9072 21055 9074
rect 14733 9016 14738 9072
rect 14794 9016 20994 9072
rect 21050 9016 21055 9072
rect 14733 9014 21055 9016
rect 14733 9011 14799 9014
rect 20989 9011 21055 9014
rect 19333 8938 19399 8941
rect 14414 8936 19399 8938
rect 14414 8880 19338 8936
rect 19394 8880 19399 8936
rect 14414 8878 19399 8880
rect 19333 8875 19399 8878
rect 23473 8938 23539 8941
rect 23473 8936 24778 8938
rect 23473 8880 23478 8936
rect 23534 8880 24778 8936
rect 23473 8878 24778 8880
rect 23473 8875 23539 8878
rect 0 8802 480 8832
rect 4061 8802 4127 8805
rect 0 8800 4127 8802
rect 0 8744 4066 8800
rect 4122 8744 4127 8800
rect 0 8742 4127 8744
rect 24718 8802 24778 8878
rect 27520 8802 28000 8832
rect 24718 8742 28000 8802
rect 0 8712 480 8742
rect 4061 8739 4127 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 27520 8712 28000 8742
rect 24277 8671 24597 8672
rect 1393 8394 1459 8397
rect 1350 8392 1459 8394
rect 1350 8336 1398 8392
rect 1454 8336 1459 8392
rect 1350 8331 1459 8336
rect 0 8258 480 8288
rect 1350 8258 1410 8331
rect 27520 8258 28000 8288
rect 0 8198 1410 8258
rect 24902 8198 28000 8258
rect 0 8168 480 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 19241 7986 19307 7989
rect 24902 7986 24962 8198
rect 27520 8168 28000 8198
rect 3926 7926 16866 7986
rect 0 7578 480 7608
rect 3926 7578 3986 7926
rect 4061 7850 4127 7853
rect 16806 7850 16866 7926
rect 19241 7984 24962 7986
rect 19241 7928 19246 7984
rect 19302 7928 24962 7984
rect 19241 7926 24962 7928
rect 19241 7923 19307 7926
rect 21265 7850 21331 7853
rect 4061 7848 16682 7850
rect 4061 7792 4066 7848
rect 4122 7792 16682 7848
rect 4061 7790 16682 7792
rect 16806 7848 21331 7850
rect 16806 7792 21270 7848
rect 21326 7792 21331 7848
rect 16806 7790 21331 7792
rect 4061 7787 4127 7790
rect 16622 7714 16682 7790
rect 21265 7787 21331 7790
rect 17953 7714 18019 7717
rect 16622 7712 18019 7714
rect 16622 7656 17958 7712
rect 18014 7656 18019 7712
rect 16622 7654 18019 7656
rect 17953 7651 18019 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 27520 7578 28000 7608
rect 0 7518 3986 7578
rect 24902 7518 28000 7578
rect 0 7488 480 7518
rect 20713 7442 20779 7445
rect 24902 7442 24962 7518
rect 27520 7488 28000 7518
rect 20713 7440 24962 7442
rect 20713 7384 20718 7440
rect 20774 7384 24962 7440
rect 20713 7382 24962 7384
rect 20713 7379 20779 7382
rect 19057 7306 19123 7309
rect 19057 7304 24962 7306
rect 19057 7248 19062 7304
rect 19118 7248 24962 7304
rect 19057 7246 24962 7248
rect 19057 7243 19123 7246
rect 10277 7104 10597 7105
rect 0 7034 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 4061 7034 4127 7037
rect 0 7032 4127 7034
rect 0 6976 4066 7032
rect 4122 6976 4127 7032
rect 0 6974 4127 6976
rect 24902 7034 24962 7246
rect 27520 7034 28000 7064
rect 24902 6974 28000 7034
rect 0 6944 480 6974
rect 4061 6971 4127 6974
rect 27520 6944 28000 6974
rect 17125 6898 17191 6901
rect 614 6896 17191 6898
rect 614 6840 17130 6896
rect 17186 6840 17191 6896
rect 614 6838 17191 6840
rect 0 6354 480 6384
rect 614 6354 674 6838
rect 17125 6835 17191 6838
rect 17309 6898 17375 6901
rect 26417 6898 26483 6901
rect 17309 6896 26483 6898
rect 17309 6840 17314 6896
rect 17370 6840 26422 6896
rect 26478 6840 26483 6896
rect 17309 6838 26483 6840
rect 17309 6835 17375 6838
rect 26417 6835 26483 6838
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 9622 6428 9628 6492
rect 9692 6490 9698 6492
rect 9692 6430 12634 6490
rect 9692 6428 9698 6430
rect 0 6294 674 6354
rect 12574 6354 12634 6430
rect 17309 6354 17375 6357
rect 12574 6352 17375 6354
rect 12574 6296 17314 6352
rect 17370 6296 17375 6352
rect 12574 6294 17375 6296
rect 0 6264 480 6294
rect 17309 6291 17375 6294
rect 18781 6354 18847 6357
rect 27520 6354 28000 6384
rect 18781 6352 28000 6354
rect 18781 6296 18786 6352
rect 18842 6296 28000 6352
rect 18781 6294 28000 6296
rect 18781 6291 18847 6294
rect 27520 6264 28000 6294
rect 9581 6220 9647 6221
rect 9581 6216 9628 6220
rect 9692 6218 9698 6220
rect 9581 6160 9586 6216
rect 9581 6156 9628 6160
rect 9692 6158 9774 6218
rect 9692 6156 9698 6158
rect 9581 6155 9647 6156
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 0 5810 480 5840
rect 1393 5810 1459 5813
rect 0 5808 1459 5810
rect 0 5752 1398 5808
rect 1454 5752 1459 5808
rect 0 5750 1459 5752
rect 0 5720 480 5750
rect 1393 5747 1459 5750
rect 23657 5810 23723 5813
rect 27520 5810 28000 5840
rect 23657 5808 28000 5810
rect 23657 5752 23662 5808
rect 23718 5752 28000 5808
rect 23657 5750 28000 5752
rect 23657 5747 23723 5750
rect 27520 5720 28000 5750
rect 8293 5674 8359 5677
rect 14365 5674 14431 5677
rect 8293 5672 14431 5674
rect 8293 5616 8298 5672
rect 8354 5616 14370 5672
rect 14426 5616 14431 5672
rect 8293 5614 14431 5616
rect 8293 5611 8359 5614
rect 14365 5611 14431 5614
rect 13261 5538 13327 5541
rect 14181 5538 14247 5541
rect 13261 5536 14247 5538
rect 13261 5480 13266 5536
rect 13322 5480 14186 5536
rect 14242 5480 14247 5536
rect 13261 5478 14247 5480
rect 13261 5475 13327 5478
rect 14181 5475 14247 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 4061 5266 4127 5269
rect 14549 5266 14615 5269
rect 4061 5264 14615 5266
rect 4061 5208 4066 5264
rect 4122 5208 14554 5264
rect 14610 5208 14615 5264
rect 4061 5206 14615 5208
rect 4061 5203 4127 5206
rect 14549 5203 14615 5206
rect 0 5130 480 5160
rect 3877 5130 3943 5133
rect 0 5128 3943 5130
rect 0 5072 3882 5128
rect 3938 5072 3943 5128
rect 0 5070 3943 5072
rect 0 5040 480 5070
rect 3877 5067 3943 5070
rect 5073 5130 5139 5133
rect 13721 5130 13787 5133
rect 5073 5128 13787 5130
rect 5073 5072 5078 5128
rect 5134 5072 13726 5128
rect 13782 5072 13787 5128
rect 5073 5070 13787 5072
rect 5073 5067 5139 5070
rect 13721 5067 13787 5070
rect 20989 5130 21055 5133
rect 27520 5130 28000 5160
rect 20989 5128 28000 5130
rect 20989 5072 20994 5128
rect 21050 5072 28000 5128
rect 20989 5070 28000 5072
rect 20989 5067 21055 5070
rect 27520 5040 28000 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 0 4586 480 4616
rect 4061 4586 4127 4589
rect 0 4584 4127 4586
rect 0 4528 4066 4584
rect 4122 4528 4127 4584
rect 0 4526 4127 4528
rect 0 4496 480 4526
rect 4061 4523 4127 4526
rect 16389 4586 16455 4589
rect 27520 4586 28000 4616
rect 16389 4584 28000 4586
rect 16389 4528 16394 4584
rect 16450 4528 28000 4584
rect 16389 4526 28000 4528
rect 16389 4523 16455 4526
rect 27520 4496 28000 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 13721 4042 13787 4045
rect 19517 4042 19583 4045
rect 13721 4040 19583 4042
rect 13721 3984 13726 4040
rect 13782 3984 19522 4040
rect 19578 3984 19583 4040
rect 13721 3982 19583 3984
rect 13721 3979 13787 3982
rect 19517 3979 19583 3982
rect 0 3906 480 3936
rect 8293 3906 8359 3909
rect 0 3904 8359 3906
rect 0 3848 8298 3904
rect 8354 3848 8359 3904
rect 0 3846 8359 3848
rect 0 3816 480 3846
rect 8293 3843 8359 3846
rect 24117 3906 24183 3909
rect 27520 3906 28000 3936
rect 24117 3904 28000 3906
rect 24117 3848 24122 3904
rect 24178 3848 28000 3904
rect 24117 3846 28000 3848
rect 24117 3843 24183 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 27520 3816 28000 3846
rect 19610 3775 19930 3776
rect 8845 3634 8911 3637
rect 13905 3634 13971 3637
rect 8845 3632 13971 3634
rect 8845 3576 8850 3632
rect 8906 3576 13910 3632
rect 13966 3576 13971 3632
rect 8845 3574 13971 3576
rect 8845 3571 8911 3574
rect 13905 3571 13971 3574
rect 14825 3634 14891 3637
rect 23473 3634 23539 3637
rect 14825 3632 23539 3634
rect 14825 3576 14830 3632
rect 14886 3576 23478 3632
rect 23534 3576 23539 3632
rect 14825 3574 23539 3576
rect 14825 3571 14891 3574
rect 23473 3571 23539 3574
rect 2773 3498 2839 3501
rect 12433 3498 12499 3501
rect 2773 3496 12499 3498
rect 2773 3440 2778 3496
rect 2834 3440 12438 3496
rect 12494 3440 12499 3496
rect 2773 3438 12499 3440
rect 2773 3435 2839 3438
rect 12433 3435 12499 3438
rect 13077 3498 13143 3501
rect 24669 3498 24735 3501
rect 13077 3496 24735 3498
rect 13077 3440 13082 3496
rect 13138 3440 24674 3496
rect 24730 3440 24735 3496
rect 13077 3438 24735 3440
rect 13077 3435 13143 3438
rect 24669 3435 24735 3438
rect 0 3362 480 3392
rect 2865 3362 2931 3365
rect 0 3360 2931 3362
rect 0 3304 2870 3360
rect 2926 3304 2931 3360
rect 0 3302 2931 3304
rect 0 3272 480 3302
rect 2865 3299 2931 3302
rect 24761 3362 24827 3365
rect 27520 3362 28000 3392
rect 24761 3360 28000 3362
rect 24761 3304 24766 3360
rect 24822 3304 28000 3360
rect 24761 3302 28000 3304
rect 24761 3299 24827 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 27520 3272 28000 3302
rect 24277 3231 24597 3232
rect 8293 2954 8359 2957
rect 12433 2954 12499 2957
rect 8293 2952 12499 2954
rect 8293 2896 8298 2952
rect 8354 2896 12438 2952
rect 12494 2896 12499 2952
rect 8293 2894 12499 2896
rect 8293 2891 8359 2894
rect 12433 2891 12499 2894
rect 10277 2752 10597 2753
rect 0 2682 480 2712
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 565 2682 631 2685
rect 0 2680 631 2682
rect 0 2624 570 2680
rect 626 2624 631 2680
rect 0 2622 631 2624
rect 0 2592 480 2622
rect 565 2619 631 2622
rect 24117 2682 24183 2685
rect 27520 2682 28000 2712
rect 24117 2680 28000 2682
rect 24117 2624 24122 2680
rect 24178 2624 28000 2680
rect 24117 2622 28000 2624
rect 24117 2619 24183 2622
rect 27520 2592 28000 2622
rect 12709 2546 12775 2549
rect 14641 2546 14707 2549
rect 12709 2544 14707 2546
rect 12709 2488 12714 2544
rect 12770 2488 14646 2544
rect 14702 2488 14707 2544
rect 12709 2486 14707 2488
rect 12709 2483 12775 2486
rect 14641 2483 14707 2486
rect 5610 2208 5930 2209
rect 0 2138 480 2168
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 3509 2138 3575 2141
rect 0 2136 3575 2138
rect 0 2080 3514 2136
rect 3570 2080 3575 2136
rect 0 2078 3575 2080
rect 0 2048 480 2078
rect 3509 2075 3575 2078
rect 24669 2138 24735 2141
rect 27520 2138 28000 2168
rect 24669 2136 28000 2138
rect 24669 2080 24674 2136
rect 24730 2080 28000 2136
rect 24669 2078 28000 2080
rect 24669 2075 24735 2078
rect 27520 2048 28000 2078
rect 0 1458 480 1488
rect 3877 1458 3943 1461
rect 0 1456 3943 1458
rect 0 1400 3882 1456
rect 3938 1400 3943 1456
rect 0 1398 3943 1400
rect 0 1368 480 1398
rect 3877 1395 3943 1398
rect 14181 1458 14247 1461
rect 27520 1458 28000 1488
rect 14181 1456 28000 1458
rect 14181 1400 14186 1456
rect 14242 1400 28000 1456
rect 14181 1398 28000 1400
rect 14181 1395 14247 1398
rect 27520 1368 28000 1398
rect 0 914 480 944
rect 3233 914 3299 917
rect 27520 914 28000 944
rect 0 912 3299 914
rect 0 856 3238 912
rect 3294 856 3299 912
rect 0 854 3299 856
rect 0 824 480 854
rect 3233 851 3299 854
rect 27478 824 28000 914
rect 27478 642 27538 824
rect 26926 582 27538 642
rect 26926 506 26986 582
rect 21406 446 26986 506
rect 0 370 480 400
rect 4061 370 4127 373
rect 0 368 4127 370
rect 0 312 4066 368
rect 4122 312 4127 368
rect 0 310 4127 312
rect 0 280 480 310
rect 4061 307 4127 310
rect 12893 98 12959 101
rect 21406 98 21466 446
rect 23473 370 23539 373
rect 27520 370 28000 400
rect 23473 368 28000 370
rect 23473 312 23478 368
rect 23534 312 28000 368
rect 23473 310 28000 312
rect 23473 307 23539 310
rect 27520 280 28000 310
rect 12893 96 21466 98
rect 12893 40 12898 96
rect 12954 40 21466 96
rect 12893 38 21466 40
rect 12893 35 12959 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 13124 25332 13188 25396
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 23428 24788 23492 24852
rect 23980 24788 24044 24852
rect 10916 24244 10980 24308
rect 13492 24168 13556 24172
rect 13492 24112 13542 24168
rect 13542 24112 13556 24168
rect 13492 24108 13556 24112
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 13308 22204 13372 22268
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 13308 21660 13372 21724
rect 13124 21252 13188 21316
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 14780 20980 14844 21044
rect 24716 20980 24780 21044
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 13492 20572 13556 20636
rect 12020 20436 12084 20500
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 14780 19756 14844 19820
rect 22692 19892 22756 19956
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 12020 19484 12084 19548
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 23980 17716 24044 17780
rect 24900 17444 24964 17508
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 23060 17308 23124 17372
rect 15516 17036 15580 17100
rect 22508 16960 22572 16964
rect 22508 16904 22522 16960
rect 22522 16904 22572 16960
rect 22508 16900 22572 16904
rect 23980 16900 24044 16964
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 24900 16416 24964 16420
rect 24900 16360 24914 16416
rect 24914 16360 24964 16416
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24900 16356 24964 16360
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 22876 16144 22940 16148
rect 22876 16088 22926 16144
rect 22926 16088 22940 16144
rect 22876 16084 22940 16088
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 22692 14996 22756 15060
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 22140 14648 22204 14652
rect 22140 14592 22190 14648
rect 22190 14592 22204 14648
rect 22140 14588 22204 14592
rect 22508 14588 22572 14652
rect 22876 14588 22940 14652
rect 19380 14452 19444 14516
rect 23980 14316 24044 14380
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 23612 13228 23676 13292
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 19380 12956 19444 13020
rect 23428 12956 23492 13020
rect 23796 12820 23860 12884
rect 23612 12684 23676 12748
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 24716 12820 24780 12884
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 23796 12412 23860 12476
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 23612 11248 23676 11252
rect 23612 11192 23662 11248
rect 23662 11192 23676 11248
rect 23612 11188 23676 11192
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 24900 10100 24964 10164
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 9628 6428 9692 6492
rect 9628 6216 9692 6220
rect 9628 6160 9642 6216
rect 9642 6160 9692 6216
rect 9628 6156 9692 6160
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 13123 25396 13189 25397
rect 13123 25332 13124 25396
rect 13188 25332 13189 25396
rect 13123 25331 13189 25332
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10915 24308 10981 24309
rect 10915 24244 10916 24308
rect 10980 24244 10981 24308
rect 10915 24243 10981 24244
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10918 14738 10978 24243
rect 13126 21317 13186 25331
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 13491 24172 13557 24173
rect 13491 24108 13492 24172
rect 13556 24108 13557 24172
rect 13491 24107 13557 24108
rect 13307 22268 13373 22269
rect 13307 22204 13308 22268
rect 13372 22204 13373 22268
rect 13307 22203 13373 22204
rect 13310 21725 13370 22203
rect 13307 21724 13373 21725
rect 13307 21660 13308 21724
rect 13372 21660 13373 21724
rect 13307 21659 13373 21660
rect 13123 21316 13189 21317
rect 13123 21252 13124 21316
rect 13188 21252 13189 21316
rect 13123 21251 13189 21252
rect 13494 20637 13554 24107
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14779 21044 14845 21045
rect 14779 20980 14780 21044
rect 14844 20980 14845 21044
rect 14779 20979 14845 20980
rect 13491 20636 13557 20637
rect 13491 20572 13492 20636
rect 13556 20572 13557 20636
rect 13491 20571 13557 20572
rect 12019 20500 12085 20501
rect 12019 20436 12020 20500
rect 12084 20436 12085 20500
rect 12019 20435 12085 20436
rect 12022 19549 12082 20435
rect 14782 19821 14842 20979
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14779 19820 14845 19821
rect 14779 19756 14780 19820
rect 14844 19756 14845 19820
rect 14779 19755 14845 19756
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 12019 19548 12085 19549
rect 12019 19484 12020 19548
rect 12084 19484 12085 19548
rect 12019 19483 12085 19484
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 23427 24852 23493 24853
rect 23427 24788 23428 24852
rect 23492 24788 23493 24852
rect 23427 24787 23493 24788
rect 23979 24852 24045 24853
rect 23979 24788 23980 24852
rect 24044 24788 24045 24852
rect 23979 24787 24045 24788
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 22691 19956 22757 19957
rect 22691 19892 22692 19956
rect 22756 19892 22757 19956
rect 22691 19891 22757 19892
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 15518 17101 15578 17222
rect 15515 17100 15581 17101
rect 15515 17036 15516 17100
rect 15580 17036 15581 17100
rect 15515 17035 15581 17036
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 9627 6492 9693 6493
rect 9627 6428 9628 6492
rect 9692 6428 9693 6492
rect 9627 6427 9693 6428
rect 9630 6221 9690 6427
rect 9627 6220 9693 6221
rect 9627 6156 9628 6220
rect 9692 6156 9693 6220
rect 9627 6155 9693 6156
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 14176 15264 15200
rect 19610 16896 19930 17920
rect 22507 16964 22573 16965
rect 22507 16900 22508 16964
rect 22572 16900 22573 16964
rect 22507 16899 22573 16900
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19379 14516 19445 14517
rect 19379 14452 19380 14516
rect 19444 14452 19445 14516
rect 19379 14451 19445 14452
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 19382 13021 19442 14451
rect 19610 13632 19930 14656
rect 22510 14653 22570 16899
rect 22694 15061 22754 19891
rect 22875 16148 22941 16149
rect 22875 16084 22876 16148
rect 22940 16084 22941 16148
rect 22875 16083 22941 16084
rect 22691 15060 22757 15061
rect 22691 14996 22692 15060
rect 22756 14996 22757 15060
rect 22691 14995 22757 14996
rect 22878 14653 22938 16083
rect 22507 14652 22573 14653
rect 22507 14588 22508 14652
rect 22572 14588 22573 14652
rect 22507 14587 22573 14588
rect 22875 14652 22941 14653
rect 22875 14588 22876 14652
rect 22940 14588 22941 14652
rect 22875 14587 22941 14588
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19379 13020 19445 13021
rect 19379 12956 19380 13020
rect 19444 12956 19445 13020
rect 19379 12955 19445 12956
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 12544 19930 13568
rect 23430 13021 23490 24787
rect 23982 18730 24042 24787
rect 23614 18670 24042 18730
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24715 21044 24781 21045
rect 24715 20980 24716 21044
rect 24780 20980 24781 21044
rect 24715 20979 24781 20980
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 23614 13293 23674 18670
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 23979 17780 24045 17781
rect 23979 17716 23980 17780
rect 24044 17716 24045 17780
rect 23979 17715 24045 17716
rect 23982 16965 24042 17715
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 23979 16964 24045 16965
rect 23979 16900 23980 16964
rect 24044 16900 24045 16964
rect 23979 16899 24045 16900
rect 23982 14381 24042 16899
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 23979 14380 24045 14381
rect 23979 14316 23980 14380
rect 24044 14316 24045 14380
rect 23979 14315 24045 14316
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 23611 13292 23677 13293
rect 23611 13228 23612 13292
rect 23676 13228 23677 13292
rect 23611 13227 23677 13228
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 23427 13020 23493 13021
rect 23427 12956 23428 13020
rect 23492 12956 23493 13020
rect 23427 12955 23493 12956
rect 23795 12884 23861 12885
rect 23795 12820 23796 12884
rect 23860 12820 23861 12884
rect 23795 12819 23861 12820
rect 23611 12748 23677 12749
rect 23611 12684 23612 12748
rect 23676 12684 23677 12748
rect 23611 12683 23677 12684
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 23614 11253 23674 12683
rect 23798 12477 23858 12819
rect 23795 12476 23861 12477
rect 23795 12412 23796 12476
rect 23860 12412 23861 12476
rect 23795 12411 23861 12412
rect 24277 12000 24597 13024
rect 24718 12885 24778 20979
rect 24899 17508 24965 17509
rect 24899 17444 24900 17508
rect 24964 17444 24965 17508
rect 24899 17443 24965 17444
rect 24902 16421 24962 17443
rect 24899 16420 24965 16421
rect 24899 16356 24900 16420
rect 24964 16356 24965 16420
rect 24899 16355 24965 16356
rect 24715 12884 24781 12885
rect 24715 12820 24716 12884
rect 24780 12820 24781 12884
rect 24715 12819 24781 12820
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 23611 11252 23677 11253
rect 23611 11188 23612 11252
rect 23676 11188 23677 11252
rect 23611 11187 23677 11188
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24902 10165 24962 16355
rect 24899 10164 24965 10165
rect 24899 10100 24900 10164
rect 24964 10100 24965 10164
rect 24899 10099 24965 10100
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 15430 17222 15666 17458
rect 10830 14502 11066 14738
rect 22054 14652 22290 14738
rect 22974 17372 23210 17458
rect 22974 17308 23060 17372
rect 23060 17308 23124 17372
rect 23124 17308 23210 17372
rect 22974 17222 23210 17308
rect 22054 14588 22140 14652
rect 22140 14588 22204 14652
rect 22204 14588 22290 14652
rect 22054 14502 22290 14588
<< metal5 >>
rect 15388 17458 23252 17500
rect 15388 17222 15430 17458
rect 15666 17222 22974 17458
rect 23210 17222 23252 17458
rect 15388 17180 23252 17222
rect 10788 14738 22332 14780
rect 10788 14502 10830 14738
rect 11066 14502 22054 14738
rect 22290 14502 22332 14738
rect 10788 14460 22332 14502
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12696 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_0_142
timestamp 1604681595
transform 1 0 14168 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604681595
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1604681595
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604681595
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604681595
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _057_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1604681595
transform 1 0 24380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1604681595
transform 1 0 25484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604681595
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604681595
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1604681595
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604681595
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_7
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_19
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_31
timestamp 1604681595
transform 1 0 3956 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_43
timestamp 1604681595
transform 1 0 5060 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_55
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604681595
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_7
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_19
timestamp 1604681595
transform 1 0 2852 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604681595
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604681595
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604681595
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604681595
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604681595
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1604681595
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1604681595
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1604681595
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1604681595
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1604681595
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604681595
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1604681595
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_23
timestamp 1604681595
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_35
timestamp 1604681595
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_47
timestamp 1604681595
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1604681595
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1604681595
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1604681595
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1604681595
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1604681595
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1604681595
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1604681595
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1604681595
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 24564 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 24564 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_259
timestamp 1604681595
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_263
timestamp 1604681595
transform 1 0 25300 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_259
timestamp 1604681595
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_275
timestamp 1604681595
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1604681595
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_7
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_11
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_16
timestamp 1604681595
transform 1 0 2576 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_28
timestamp 1604681595
transform 1 0 3680 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_40
timestamp 1604681595
transform 1 0 4784 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_52
timestamp 1604681595
transform 1 0 5888 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1604681595
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 12972 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 13340 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_131
timestamp 1604681595
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_135
timestamp 1604681595
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_139
timestamp 1604681595
transform 1 0 13892 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_149
timestamp 1604681595
transform 1 0 14812 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_153
timestamp 1604681595
transform 1 0 15180 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_156
timestamp 1604681595
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_160
timestamp 1604681595
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_164
timestamp 1604681595
transform 1 0 16192 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_176
timestamp 1604681595
transform 1 0 17296 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1604681595
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_228
timestamp 1604681595
transform 1 0 22080 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 23828 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_233
timestamp 1604681595
transform 1 0 22540 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_241
timestamp 1604681595
transform 1 0 23276 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_249
timestamp 1604681595
transform 1 0 24012 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_259
timestamp 1604681595
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_263
timestamp 1604681595
transform 1 0 25300 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_275
timestamp 1604681595
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_7
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_12
timestamp 1604681595
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_16
timestamp 1604681595
transform 1 0 2576 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_20
timestamp 1604681595
transform 1 0 2944 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11408 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_105
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_111
timestamp 1604681595
transform 1 0 11316 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_114
timestamp 1604681595
transform 1 0 11592 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_124
timestamp 1604681595
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_128
timestamp 1604681595
transform 1 0 12880 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_138
timestamp 1604681595
transform 1 0 13800 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_144
timestamp 1604681595
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_148
timestamp 1604681595
transform 1 0 14720 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17204 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_167
timestamp 1604681595
transform 1 0 16468 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_173
timestamp 1604681595
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1604681595
transform 1 0 17388 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_189
timestamp 1604681595
transform 1 0 18492 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1604681595
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604681595
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 23460 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 22356 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24012 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_235
timestamp 1604681595
transform 1 0 22724 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_247
timestamp 1604681595
transform 1 0 23828 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 24564 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_259
timestamp 1604681595
transform 1 0 24932 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_271
timestamp 1604681595
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_12
timestamp 1604681595
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_16
timestamp 1604681595
transform 1 0 2576 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 3036 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_30
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_34
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_38
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_42
timestamp 1604681595
transform 1 0 4968 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_54
timestamp 1604681595
transform 1 0 6072 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1604681595
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_98
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_106
timestamp 1604681595
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12696 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1604681595
transform 1 0 13892 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_143
timestamp 1604681595
transform 1 0 14260 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16100 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 14536 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1604681595
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_159
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1604681595
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_176
timestamp 1604681595
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1604681595
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 18584 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1604681595
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_192
timestamp 1604681595
transform 1 0 18768 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_204
timestamp 1604681595
transform 1 0 19872 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _030_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 21436 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 21896 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_216
timestamp 1604681595
transform 1 0 20976 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_224
timestamp 1604681595
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_228
timestamp 1604681595
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604681595
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 22448 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604681595
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23828 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24012 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 25576 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_258
timestamp 1604681595
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_262
timestamp 1604681595
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_7
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp 1604681595
transform 1 0 2116 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_45
timestamp 1604681595
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_49
timestamp 1604681595
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_53
timestamp 1604681595
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_61
timestamp 1604681595
transform 1 0 6716 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_57
timestamp 1604681595
transform 1 0 6348 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8280 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 8648 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_64
timestamp 1604681595
transform 1 0 6992 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_72
timestamp 1604681595
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_76
timestamp 1604681595
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 10396 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_97
timestamp 1604681595
transform 1 0 10028 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_103
timestamp 1604681595
transform 1 0 10580 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11408 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_107
timestamp 1604681595
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_111
timestamp 1604681595
transform 1 0 11316 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1604681595
transform 1 0 12236 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_125
timestamp 1604681595
transform 1 0 12604 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12972 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_128
timestamp 1604681595
transform 1 0 12880 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1604681595
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_142
timestamp 1604681595
transform 1 0 14168 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_148
timestamp 1604681595
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 17848 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1604681595
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_180
timestamp 1604681595
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_184
timestamp 1604681595
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1604681595
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_188
timestamp 1604681595
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_193
timestamp 1604681595
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1604681595
transform 1 0 19228 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_201
timestamp 1604681595
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_206
timestamp 1604681595
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 21620 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_227
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 22724 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23828 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_239
timestamp 1604681595
transform 1 0 23092 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 25392 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24840 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_256
timestamp 1604681595
transform 1 0 24656 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_260
timestamp 1604681595
transform 1 0 25024 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_267
timestamp 1604681595
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_7
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_10
timestamp 1604681595
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_16
timestamp 1604681595
transform 1 0 2576 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_12
timestamp 1604681595
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2668 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_30
timestamp 1604681595
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_26
timestamp 1604681595
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4232 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_41
timestamp 1604681595
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_46
timestamp 1604681595
transform 1 0 5336 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_52
timestamp 1604681595
transform 1 0 5888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_47
timestamp 1604681595
transform 1 0 5428 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1604681595
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 5704 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1604681595
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_66
timestamp 1604681595
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_71
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_76
timestamp 1604681595
transform 1 0 8096 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7912 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 8648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_83
timestamp 1604681595
transform 1 0 8740 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_90
timestamp 1604681595
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_85
timestamp 1604681595
transform 1 0 8924 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_97
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 9752 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_122
timestamp 1604681595
transform 1 0 12328 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_118
timestamp 1604681595
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12972 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12696 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_128
timestamp 1604681595
transform 1 0 12880 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_145
timestamp 1604681595
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_150
timestamp 1604681595
transform 1 0 14904 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_146
timestamp 1604681595
transform 1 0 14536 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_149
timestamp 1604681595
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15180 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1604681595
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1604681595
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1604681595
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_174
timestamp 1604681595
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_167
timestamp 1604681595
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_173
timestamp 1604681595
transform 1 0 17020 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17296 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 16744 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1604681595
transform 1 0 16836 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_178
timestamp 1604681595
transform 1 0 17480 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 17848 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_185
timestamp 1604681595
transform 1 0 18124 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18216 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_195
timestamp 1604681595
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_189
timestamp 1604681595
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18860 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_199
timestamp 1604681595
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_202
timestamp 1604681595
transform 1 0 19688 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 19872 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 19780 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_206
timestamp 1604681595
transform 1 0 20056 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604681595
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_210
timestamp 1604681595
transform 1 0 20424 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 20516 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_225
timestamp 1604681595
transform 1 0 21804 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_224
timestamp 1604681595
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 21896 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 21436 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_228
timestamp 1604681595
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_237
timestamp 1604681595
transform 1 0 22908 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 22540 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_247
timestamp 1604681595
transform 1 0 23828 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24012 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 25300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_261
timestamp 1604681595
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_265
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_255
timestamp 1604681595
transform 1 0 24564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_259
timestamp 1604681595
transform 1 0 24932 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_267
timestamp 1604681595
transform 1 0 25668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2852 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_9
timestamp 1604681595
transform 1 0 1932 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_13
timestamp 1604681595
transform 1 0 2300 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_16
timestamp 1604681595
transform 1 0 2576 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4876 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_35
timestamp 1604681595
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_39
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_43
timestamp 1604681595
transform 1 0 5060 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_78
timestamp 1604681595
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_82
timestamp 1604681595
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_102
timestamp 1604681595
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_106
timestamp 1604681595
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1604681595
transform 1 0 11500 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14352 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_143
timestamp 1604681595
transform 1 0 14260 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_160
timestamp 1604681595
transform 1 0 15824 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_164
timestamp 1604681595
transform 1 0 16192 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_167
timestamp 1604681595
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 19596 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1604681595
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_197
timestamp 1604681595
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 21896 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21712 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_210
timestamp 1604681595
transform 1 0 20424 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_214
timestamp 1604681595
transform 1 0 20792 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_217
timestamp 1604681595
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1604681595
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_230
timestamp 1604681595
transform 1 0 22264 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1604681595
transform 1 0 25116 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_273
timestamp 1604681595
transform 1 0 26220 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_6
timestamp 1604681595
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_10
timestamp 1604681595
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4232 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5796 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_43
timestamp 1604681595
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_47
timestamp 1604681595
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_67
timestamp 1604681595
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_71
timestamp 1604681595
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9752 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_100
timestamp 1604681595
transform 1 0 10304 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_104
timestamp 1604681595
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11040 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_124
timestamp 1604681595
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13248 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_128
timestamp 1604681595
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_161
timestamp 1604681595
transform 1 0 15916 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_157
timestamp 1604681595
transform 1 0 15548 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 15732 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16284 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17848 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_174
timestamp 1604681595
transform 1 0 17112 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_180
timestamp 1604681595
transform 1 0 17664 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 19596 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19964 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_198
timestamp 1604681595
transform 1 0 19320 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_203
timestamp 1604681595
transform 1 0 19780 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_207
timestamp 1604681595
transform 1 0 20148 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20332 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 21896 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_219
timestamp 1604681595
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_223
timestamp 1604681595
transform 1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_228
timestamp 1604681595
transform 1 0 22080 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22632 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22264 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 24012 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_232
timestamp 1604681595
transform 1 0 22448 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_243
timestamp 1604681595
transform 1 0 23460 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_247
timestamp 1604681595
transform 1 0 23828 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24932 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_257
timestamp 1604681595
transform 1 0 24748 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_261
timestamp 1604681595
transform 1 0 25116 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_273
timestamp 1604681595
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2760 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_9
timestamp 1604681595
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_13
timestamp 1604681595
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_17
timestamp 1604681595
transform 1 0 2668 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_34
timestamp 1604681595
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_38
timestamp 1604681595
transform 1 0 4600 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 8556 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6992 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_73
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_77
timestamp 1604681595
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9752 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_84
timestamp 1604681595
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_88
timestamp 1604681595
transform 1 0 9200 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_136
timestamp 1604681595
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 1604681595
transform 1 0 13984 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_144
timestamp 1604681595
transform 1 0 14352 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_163
timestamp 1604681595
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_167
timestamp 1604681595
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18124 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20148 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_201
timestamp 1604681595
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_205
timestamp 1604681595
transform 1 0 19964 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20332 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21896 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 1604681595
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1604681595
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 22632 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604681595
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 25208 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_254
timestamp 1604681595
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_258
timestamp 1604681595
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_266
timestamp 1604681595
transform 1 0 25576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_270
timestamp 1604681595
transform 1 0 25944 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_276
timestamp 1604681595
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1932 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1604681595
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_18
timestamp 1604681595
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_22
timestamp 1604681595
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_26
timestamp 1604681595
transform 1 0 3496 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6072 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 5704 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_48
timestamp 1604681595
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_52
timestamp 1604681595
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_65
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_69
timestamp 1604681595
transform 1 0 7452 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_88
timestamp 1604681595
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 9752 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1604681595
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_101
timestamp 1604681595
transform 1 0 10396 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_121
timestamp 1604681595
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_125
timestamp 1604681595
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1604681595
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_142
timestamp 1604681595
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14720 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_146
timestamp 1604681595
transform 1 0 14536 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1604681595
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 16928 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17296 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 1604681595
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_174
timestamp 1604681595
transform 1 0 17112 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1604681595
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1604681595
transform 1 0 18216 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18400 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1604681595
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_224
timestamp 1604681595
transform 1 0 21712 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_229
timestamp 1604681595
transform 1 0 22172 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 22448 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 24104 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_248
timestamp 1604681595
transform 1 0 23920 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24656 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 24472 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_252
timestamp 1604681595
transform 1 0 24288 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_265
timestamp 1604681595
transform 1 0 25484 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_273
timestamp 1604681595
transform 1 0 26220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2852 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_9
timestamp 1604681595
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_13
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_28
timestamp 1604681595
transform 1 0 3680 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_34
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7728 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_65
timestamp 1604681595
transform 1 0 7084 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_70
timestamp 1604681595
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_90
timestamp 1604681595
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_94
timestamp 1604681595
transform 1 0 9752 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1604681595
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 13984 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1604681595
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_136
timestamp 1604681595
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15548 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_149
timestamp 1604681595
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_153
timestamp 1604681595
transform 1 0 15180 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1604681595
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_174
timestamp 1604681595
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_170
timestamp 1604681595
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1604681595
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_178
timestamp 1604681595
transform 1 0 17480 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17664 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 19872 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_200
timestamp 1604681595
transform 1 0 19504 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_206
timestamp 1604681595
transform 1 0 20056 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1604681595
transform 1 0 20424 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_219
timestamp 1604681595
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_223
timestamp 1604681595
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 25208 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_254
timestamp 1604681595
transform 1 0 24472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_258
timestamp 1604681595
transform 1 0 24840 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_261
timestamp 1604681595
transform 1 0 25116 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_266
timestamp 1604681595
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_270
timestamp 1604681595
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 26128 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_274
timestamp 1604681595
transform 1 0 26312 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1840 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1748 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_17
timestamp 1604681595
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_16
timestamp 1604681595
transform 1 0 2576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 3404 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_21
timestamp 1604681595
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_25
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_21
timestamp 1604681595
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1604681595
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_33
timestamp 1604681595
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_40
timestamp 1604681595
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_36
timestamp 1604681595
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4600 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_53
timestamp 1604681595
transform 1 0 5980 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_53
timestamp 1604681595
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 6716 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6532 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_57
timestamp 1604681595
transform 1 0 6348 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1604681595
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_71
timestamp 1604681595
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_67
timestamp 1604681595
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_69
timestamp 1604681595
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_65
timestamp 1604681595
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 6992 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1604681595
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8004 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1604681595
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_86
timestamp 1604681595
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_95
timestamp 1604681595
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1604681595
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9844 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10212 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_112
timestamp 1604681595
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1604681595
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_116
timestamp 1604681595
transform 1 0 11776 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_125
timestamp 1604681595
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 11132 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13340 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 14444 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13156 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_142
timestamp 1604681595
transform 1 0 14168 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_139
timestamp 1604681595
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_143
timestamp 1604681595
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_156
timestamp 1604681595
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_146
timestamp 1604681595
transform 1 0 14536 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 14628 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_160
timestamp 1604681595
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15456 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_173
timestamp 1604681595
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1604681595
transform 1 0 17296 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_172
timestamp 1604681595
transform 1 0 16928 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17112 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_177
timestamp 1604681595
transform 1 0 17388 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 17664 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 18308 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_193
timestamp 1604681595
transform 1 0 18860 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_189
timestamp 1604681595
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_193
timestamp 1604681595
transform 1 0 18860 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_189
timestamp 1604681595
transform 1 0 18492 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19044 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 18676 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 18676 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1604681595
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18952 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_27_217
timestamp 1604681595
transform 1 0 21068 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_214
timestamp 1604681595
transform 1 0 20792 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_210
timestamp 1604681595
transform 1 0 20424 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1604681595
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_228
timestamp 1604681595
transform 1 0 22080 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_224
timestamp 1604681595
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21160 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 22724 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22448 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_234
timestamp 1604681595
transform 1 0 22632 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_234
timestamp 1604681595
transform 1 0 22632 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604681595
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_258
timestamp 1604681595
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1604681595
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_255
timestamp 1604681595
transform 1 0 24564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 24380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_267
timestamp 1604681595
transform 1 0 25668 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 24932 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_268
timestamp 1604681595
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 26312 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_272
timestamp 1604681595
transform 1 0 26128 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_276
timestamp 1604681595
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_36
timestamp 1604681595
transform 1 0 4416 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_40
timestamp 1604681595
transform 1 0 4784 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_3_
timestamp 1604681595
transform 1 0 5244 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6440 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_43
timestamp 1604681595
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1604681595
transform 1 0 6072 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_60
timestamp 1604681595
transform 1 0 6624 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_64
timestamp 1604681595
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9844 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10580 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_101
timestamp 1604681595
transform 1 0 10396 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11132 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 10948 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_125
timestamp 1604681595
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13340 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_142
timestamp 1604681595
transform 1 0 14168 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_150
timestamp 1604681595
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_146
timestamp 1604681595
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14720 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 15364 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_159
timestamp 1604681595
transform 1 0 15732 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_163
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 16192 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16468 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18124 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_183
timestamp 1604681595
transform 1 0 17940 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_187
timestamp 1604681595
transform 1 0 18308 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18676 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 18492 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_200
timestamp 1604681595
transform 1 0 19504 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_204
timestamp 1604681595
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1604681595
transform 1 0 20240 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_224
timestamp 1604681595
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1604681595
transform 1 0 22080 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 24012 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 23644 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22264 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_241
timestamp 1604681595
transform 1 0 23276 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_247
timestamp 1604681595
transform 1 0 23828 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 25392 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_258
timestamp 1604681595
transform 1 0 24840 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_262
timestamp 1604681595
transform 1 0 25208 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_266
timestamp 1604681595
transform 1 0 25576 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_270
timestamp 1604681595
transform 1 0 25944 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_274
timestamp 1604681595
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 2116 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4324 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 3772 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_31
timestamp 1604681595
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6440 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_56
timestamp 1604681595
transform 1 0 6256 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_60
timestamp 1604681595
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8280 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7728 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_68
timestamp 1604681595
transform 1 0 7360 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10488 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10304 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_94
timestamp 1604681595
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12604 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_111
timestamp 1604681595
transform 1 0 11316 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_115
timestamp 1604681595
transform 1 0 11684 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 14352 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12788 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_136
timestamp 1604681595
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_140
timestamp 1604681595
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_153
timestamp 1604681595
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_157
timestamp 1604681595
transform 1 0 15548 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_162
timestamp 1604681595
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1604681595
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1604681595
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19596 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_193
timestamp 1604681595
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_197
timestamp 1604681595
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21804 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_217
timestamp 1604681595
transform 1 0 21068 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1604681595
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 22908 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23276 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_234
timestamp 1604681595
transform 1 0 22632 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_239
timestamp 1604681595
transform 1 0 23092 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_243
timestamp 1604681595
transform 1 0 23460 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 25300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 25668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_261
timestamp 1604681595
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_265
timestamp 1604681595
transform 1 0 25484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 26036 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_273
timestamp 1604681595
transform 1 0 26220 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1932 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1604681595
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_26
timestamp 1604681595
transform 1 0 3496 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_22
timestamp 1604681595
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_39
timestamp 1604681595
transform 1 0 4692 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_36
timestamp 1604681595
transform 1 0 4416 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 4508 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4876 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6440 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_50
timestamp 1604681595
transform 1 0 5704 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_54
timestamp 1604681595
transform 1 0 6072 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_67
timestamp 1604681595
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_71
timestamp 1604681595
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11868 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 12236 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_109
timestamp 1604681595
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_113
timestamp 1604681595
transform 1 0 11500 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_119
timestamp 1604681595
transform 1 0 12052 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_139
timestamp 1604681595
transform 1 0 13892 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_143
timestamp 1604681595
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15364 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_147
timestamp 1604681595
transform 1 0 14628 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_161
timestamp 1604681595
transform 1 0 15916 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_165
timestamp 1604681595
transform 1 0 16284 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 16652 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_168
timestamp 1604681595
transform 1 0 16560 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_185
timestamp 1604681595
transform 1 0 18124 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18860 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_189
timestamp 1604681595
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_210
timestamp 1604681595
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_224
timestamp 1604681595
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_228
timestamp 1604681595
transform 1 0 22080 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22908 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23920 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22724 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22264 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_232
timestamp 1604681595
transform 1 0 22448 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_246
timestamp 1604681595
transform 1 0 23736 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1604681595
transform 1 0 24104 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 24472 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25484 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 24288 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_267
timestamp 1604681595
transform 1 0 25668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_271
timestamp 1604681595
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2944 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_12
timestamp 1604681595
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_16
timestamp 1604681595
transform 1 0 2576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4508 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3956 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4324 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_29
timestamp 1604681595
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_33
timestamp 1604681595
transform 1 0 4140 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_53
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8556 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_77
timestamp 1604681595
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_90
timestamp 1604681595
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_94
timestamp 1604681595
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11868 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_107
timestamp 1604681595
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_111
timestamp 1604681595
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_115
timestamp 1604681595
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1604681595
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13340 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12972 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_127
timestamp 1604681595
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_131
timestamp 1604681595
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 15824 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_151
timestamp 1604681595
transform 1 0 14996 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_156
timestamp 1604681595
transform 1 0 15456 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_163
timestamp 1604681595
transform 1 0 16100 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17480 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_175
timestamp 1604681595
transform 1 0 17204 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1604681595
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_188
timestamp 1604681595
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_192
timestamp 1604681595
transform 1 0 18768 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 20792 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_212
timestamp 1604681595
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_216
timestamp 1604681595
transform 1 0 20976 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_229
timestamp 1604681595
transform 1 0 22172 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 22356 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 22724 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_233
timestamp 1604681595
transform 1 0 22540 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_237
timestamp 1604681595
transform 1 0 22908 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_241
timestamp 1604681595
transform 1 0 23276 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 25300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 25668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_261
timestamp 1604681595
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_265
timestamp 1604681595
transform 1 0 25484 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 1840 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_6
timestamp 1604681595
transform 1 0 1656 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_10
timestamp 1604681595
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4692 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4232 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_36
timestamp 1604681595
transform 1 0 4416 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6440 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_55
timestamp 1604681595
transform 1 0 6164 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_60
timestamp 1604681595
transform 1 0 6624 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1604681595
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_72
timestamp 1604681595
transform 1 0 7728 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_77
timestamp 1604681595
transform 1 0 8188 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10304 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_88
timestamp 1604681595
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_97
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11684 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_109
timestamp 1604681595
transform 1 0 11132 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_113
timestamp 1604681595
transform 1 0 11500 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13432 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 13248 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_126
timestamp 1604681595
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_130
timestamp 1604681595
transform 1 0 13064 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_143
timestamp 1604681595
transform 1 0 14260 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_147
timestamp 1604681595
transform 1 0 14628 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17296 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16928 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_170
timestamp 1604681595
transform 1 0 16744 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_174
timestamp 1604681595
transform 1 0 17112 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_187
timestamp 1604681595
transform 1 0 18308 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604681595
transform 1 0 18492 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 20240 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1604681595
transform 1 0 18676 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21896 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_210
timestamp 1604681595
transform 1 0 20424 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_224
timestamp 1604681595
transform 1 0 21712 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_228
timestamp 1604681595
transform 1 0 22080 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 22632 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22264 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_232
timestamp 1604681595
transform 1 0 22448 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1604681595
transform 1 0 24104 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24840 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24288 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 24656 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_254
timestamp 1604681595
transform 1 0 24472 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_267
timestamp 1604681595
transform 1 0 25668 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_6
timestamp 1604681595
transform 1 0 1656 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 1840 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604681595
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_10
timestamp 1604681595
transform 1 0 2024 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_23
timestamp 1604681595
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_28
timestamp 1604681595
transform 1 0 3680 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_24
timestamp 1604681595
transform 1 0 3312 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1604681595
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_32
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4508 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_34_49
timestamp 1604681595
transform 1 0 5612 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_45
timestamp 1604681595
transform 1 0 5244 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5428 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5060 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_60
timestamp 1604681595
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1604681595
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_53
timestamp 1604681595
transform 1 0 5980 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 5980 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6440 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6164 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7636 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_66
timestamp 1604681595
transform 1 0 7176 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_67
timestamp 1604681595
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_71
timestamp 1604681595
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_84
timestamp 1604681595
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_87
timestamp 1604681595
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_88
timestamp 1604681595
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_91
timestamp 1604681595
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 9844 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9844 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10028 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_34_113
timestamp 1604681595
transform 1 0 11500 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_111
timestamp 1604681595
transform 1 0 11316 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 11500 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_118
timestamp 1604681595
transform 1 0 11960 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_115
timestamp 1604681595
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 11776 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12144 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12328 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_135
timestamp 1604681595
transform 1 0 13524 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_131
timestamp 1604681595
transform 1 0 13156 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_132
timestamp 1604681595
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 13340 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_140
timestamp 1604681595
transform 1 0 13984 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_136
timestamp 1604681595
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14076 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 1604681595
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_34_163
timestamp 1604681595
transform 1 0 16100 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_161
timestamp 1604681595
transform 1 0 15916 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_157
timestamp 1604681595
transform 1 0 15548 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15732 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16100 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16284 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_177
timestamp 1604681595
transform 1 0 17388 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_172
timestamp 1604681595
transform 1 0 16928 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_168
timestamp 1604681595
transform 1 0 16560 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_174
timestamp 1604681595
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17296 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17204 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_187
timestamp 1604681595
transform 1 0 18308 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_178
timestamp 1604681595
transform 1 0 17480 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17572 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17756 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19044 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 19964 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 19596 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 18492 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_191
timestamp 1604681595
transform 1 0 18676 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1604681595
transform 1 0 19228 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_203
timestamp 1604681595
transform 1 0 19780 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_208
timestamp 1604681595
transform 1 0 20240 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1604681595
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_211
timestamp 1604681595
transform 1 0 20516 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20700 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21068 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_223
timestamp 1604681595
transform 1 0 21620 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_219
timestamp 1604681595
transform 1 0 21252 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21436 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21804 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21252 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_34_238
timestamp 1604681595
transform 1 0 23000 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_234
timestamp 1604681595
transform 1 0 22632 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_235
timestamp 1604681595
transform 1 0 22724 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 22816 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604681595
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23184 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 23368 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_34_258
timestamp 1604681595
transform 1 0 24840 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_258
timestamp 1604681595
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_254
timestamp 1604681595
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_266
timestamp 1604681595
transform 1 0 25576 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_262
timestamp 1604681595
transform 1 0 25208 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25024 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_268
timestamp 1604681595
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_272
timestamp 1604681595
transform 1 0 26128 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_276
timestamp 1604681595
transform 1 0 26496 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1604681595
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2760 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_10
timestamp 1604681595
transform 1 0 2024 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_16
timestamp 1604681595
transform 1 0 2576 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_34
timestamp 1604681595
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_38
timestamp 1604681595
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4968 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1604681595
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7360 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_66
timestamp 1604681595
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10212 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_84
timestamp 1604681595
transform 1 0 8832 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_88
timestamp 1604681595
transform 1 0 9200 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_92
timestamp 1604681595
transform 1 0 9568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_95
timestamp 1604681595
transform 1 0 9844 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_108
timestamp 1604681595
transform 1 0 11040 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_112
timestamp 1604681595
transform 1 0 11408 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13892 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_129
timestamp 1604681595
transform 1 0 12972 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_134
timestamp 1604681595
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_138
timestamp 1604681595
transform 1 0 13800 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16100 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15916 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 15548 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_155
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_159
timestamp 1604681595
transform 1 0 15732 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_172
timestamp 1604681595
transform 1 0 16928 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_176
timestamp 1604681595
transform 1 0 17296 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1604681595
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_3_
timestamp 1604681595
transform 1 0 19596 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_193
timestamp 1604681595
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_197
timestamp 1604681595
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21160 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22172 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_210
timestamp 1604681595
transform 1 0 20424 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_214
timestamp 1604681595
transform 1 0 20792 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_217
timestamp 1604681595
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_227
timestamp 1604681595
transform 1 0 21988 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 22724 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_231
timestamp 1604681595
transform 1 0 22356 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1604681595
transform 1 0 22908 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_241
timestamp 1604681595
transform 1 0 23276 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 25668 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_261
timestamp 1604681595
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_265
timestamp 1604681595
transform 1 0 25484 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_7
timestamp 1604681595
transform 1 0 1748 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_11
timestamp 1604681595
transform 1 0 2116 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_23
timestamp 1604681595
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6624 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5704 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6440 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_48
timestamp 1604681595
transform 1 0 5520 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_52
timestamp 1604681595
transform 1 0 5888 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8280 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8004 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_69
timestamp 1604681595
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_73
timestamp 1604681595
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_77
timestamp 1604681595
transform 1 0 8188 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10396 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_84
timestamp 1604681595
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_88
timestamp 1604681595
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_99
timestamp 1604681595
transform 1 0 10212 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_103
timestamp 1604681595
transform 1 0 10580 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11040 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_107
timestamp 1604681595
transform 1 0 10948 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_124
timestamp 1604681595
transform 1 0 12512 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13248 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14260 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13064 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12696 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_128
timestamp 1604681595
transform 1 0 12880 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1604681595
transform 1 0 14076 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_145
timestamp 1604681595
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_149
timestamp 1604681595
transform 1 0 14812 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604681595
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_165
timestamp 1604681595
transform 1 0 16284 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_162
timestamp 1604681595
transform 1 0 16008 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_158
timestamp 1604681595
transform 1 0 15640 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16100 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16376 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 18032 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_182
timestamp 1604681595
transform 1 0 17848 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_186
timestamp 1604681595
transform 1 0 18216 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18584 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 19596 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18400 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 19964 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_199
timestamp 1604681595
transform 1 0 19412 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1604681595
transform 1 0 19780 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_207
timestamp 1604681595
transform 1 0 20148 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_211
timestamp 1604681595
transform 1 0 20516 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_224
timestamp 1604681595
transform 1 0 21712 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_229
timestamp 1604681595
transform 1 0 22172 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 22724 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22356 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_233
timestamp 1604681595
transform 1 0 22540 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24932 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24748 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_255
timestamp 1604681595
transform 1 0 24564 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_265
timestamp 1604681595
transform 1 0 25484 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_273
timestamp 1604681595
transform 1 0 26220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2668 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_9
timestamp 1604681595
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_13
timestamp 1604681595
transform 1 0 2300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_33
timestamp 1604681595
transform 1 0 4140 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_37
timestamp 1604681595
transform 1 0 4508 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_40
timestamp 1604681595
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1604681595
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604681595
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_71
timestamp 1604681595
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_75
timestamp 1604681595
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10304 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9384 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_88
timestamp 1604681595
transform 1 0 9200 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_92
timestamp 1604681595
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_96
timestamp 1604681595
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11684 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_109
timestamp 1604681595
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1604681595
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_117
timestamp 1604681595
transform 1 0 11868 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14076 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13892 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_132
timestamp 1604681595
transform 1 0 13248 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_137
timestamp 1604681595
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16284 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16100 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15732 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_157
timestamp 1604681595
transform 1 0 15548 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_161
timestamp 1604681595
transform 1 0 15916 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17296 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_174
timestamp 1604681595
transform 1 0 17112 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_178
timestamp 1604681595
transform 1 0 17480 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20148 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19780 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_193
timestamp 1604681595
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_197
timestamp 1604681595
transform 1 0 19228 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_201
timestamp 1604681595
transform 1 0 19596 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_205
timestamp 1604681595
transform 1 0 19964 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20332 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21988 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21804 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 21436 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_218
timestamp 1604681595
transform 1 0 21160 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_223
timestamp 1604681595
transform 1 0 21620 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23736 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_236
timestamp 1604681595
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_240
timestamp 1604681595
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25300 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25116 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_255
timestamp 1604681595
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_259
timestamp 1604681595
transform 1 0 24932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_269
timestamp 1604681595
transform 1 0 25852 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 26036 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_273
timestamp 1604681595
transform 1 0 26220 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 2944 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2392 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 2760 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_12
timestamp 1604681595
transform 1 0 2208 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_16
timestamp 1604681595
transform 1 0 2576 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604681595
transform 1 0 4600 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_23
timestamp 1604681595
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_36
timestamp 1604681595
transform 1 0 4416 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_40
timestamp 1604681595
transform 1 0 4784 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_60
timestamp 1604681595
transform 1 0 6624 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7176 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_64
timestamp 1604681595
transform 1 0 6992 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_84
timestamp 1604681595
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_88
timestamp 1604681595
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_102
timestamp 1604681595
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11316 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11132 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_106
timestamp 1604681595
transform 1 0 10856 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13524 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_127
timestamp 1604681595
transform 1 0 12788 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_131
timestamp 1604681595
transform 1 0 13156 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_134
timestamp 1604681595
transform 1 0 13432 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_144
timestamp 1604681595
transform 1 0 14352 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_148
timestamp 1604681595
transform 1 0 14720 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_161
timestamp 1604681595
transform 1 0 15916 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_157
timestamp 1604681595
transform 1 0 15548 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16100 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15732 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16284 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18032 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_181
timestamp 1604681595
transform 1 0 17756 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_186
timestamp 1604681595
transform 1 0 18216 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18584 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18400 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_206
timestamp 1604681595
transform 1 0 20056 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21528 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21068 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 20332 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_211
timestamp 1604681595
transform 1 0 20516 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_219
timestamp 1604681595
transform 1 0 21252 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23736 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23184 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23552 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_238
timestamp 1604681595
transform 1 0 23000 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_242
timestamp 1604681595
transform 1 0 23368 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 25300 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24748 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_255
timestamp 1604681595
transform 1 0 24564 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_259
timestamp 1604681595
transform 1 0 24932 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_267
timestamp 1604681595
transform 1 0 25668 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_7
timestamp 1604681595
transform 1 0 1748 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_7
timestamp 1604681595
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 1932 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604681595
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1604681595
transform 1 0 2116 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_11
timestamp 1604681595
transform 1 0 2116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604681595
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_19
timestamp 1604681595
transform 1 0 2852 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_19
timestamp 1604681595
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_23
timestamp 1604681595
transform 1 0 3220 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_23
timestamp 1604681595
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1604681595
transform 1 0 3036 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604681595
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_36
timestamp 1604681595
transform 1 0 4416 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_35
timestamp 1604681595
transform 1 0 4324 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_31
timestamp 1604681595
transform 1 0 3956 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1604681595
transform 1 0 4508 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1604681595
transform 1 0 4140 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_39
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4784 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_46
timestamp 1604681595
transform 1 0 5336 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_42
timestamp 1604681595
transform 1 0 4968 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1604681595
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_53
timestamp 1604681595
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5612 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_40_69
timestamp 1604681595
transform 1 0 7452 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_65
timestamp 1604681595
transform 1 0 7084 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_71
timestamp 1604681595
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7268 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7636 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1604681595
transform 1 0 8648 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_75
timestamp 1604681595
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_90
timestamp 1604681595
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_86
timestamp 1604681595
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_92
timestamp 1604681595
transform 1 0 9568 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_88
timestamp 1604681595
transform 1 0 9200 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9200 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_102
timestamp 1604681595
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_95
timestamp 1604681595
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_111
timestamp 1604681595
transform 1 0 11316 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_106
timestamp 1604681595
transform 1 0 10856 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_106
timestamp 1604681595
transform 1 0 10856 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11132 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11500 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_124
timestamp 1604681595
transform 1 0 12512 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11684 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_40_131
timestamp 1604681595
transform 1 0 13156 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_128
timestamp 1604681595
transform 1 0 12880 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13248 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_143
timestamp 1604681595
transform 1 0 14260 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_139
timestamp 1604681595
transform 1 0 13892 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604681595
transform 1 0 14260 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 14076 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_145
timestamp 1604681595
transform 1 0 14444 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 14444 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_154
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_149
timestamp 1604681595
transform 1 0 14812 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_147
timestamp 1604681595
transform 1 0 14628 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14996 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_165
timestamp 1604681595
transform 1 0 16284 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15180 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_40_176
timestamp 1604681595
transform 1 0 17296 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1604681595
transform 1 0 16652 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_173
timestamp 1604681595
transform 1 0 17020 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1604681595
transform 1 0 16652 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16836 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16836 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16468 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 17020 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_180
timestamp 1604681595
transform 1 0 17664 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1604681595
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17480 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17848 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1604681595
transform 1 0 19228 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_193
timestamp 1604681595
transform 1 0 18860 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_201
timestamp 1604681595
transform 1 0 19596 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_200
timestamp 1604681595
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 19412 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 19688 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_206
timestamp 1604681595
transform 1 0 20056 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_204
timestamp 1604681595
transform 1 0 19872 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_210
timestamp 1604681595
transform 1 0 20424 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_228
timestamp 1604681595
transform 1 0 22080 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_224
timestamp 1604681595
transform 1 0 21712 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_229
timestamp 1604681595
transform 1 0 22172 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1604681595
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 21896 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21988 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 20332 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1604681595
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 22264 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 22540 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_247
timestamp 1604681595
transform 1 0 23828 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_241
timestamp 1604681595
transform 1 0 23276 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23644 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_255
timestamp 1604681595
transform 1 0 24564 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_258
timestamp 1604681595
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_254
timestamp 1604681595
transform 1 0 24472 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24656 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_267
timestamp 1604681595
transform 1 0 25668 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_266
timestamp 1604681595
transform 1 0 25576 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 25300 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 25208 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_270
timestamp 1604681595
transform 1 0 25944 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 25760 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_276
timestamp 1604681595
transform 1 0 26496 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1604681595
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604681595
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1604681595
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1604681595
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_19
timestamp 1604681595
transform 1 0 2852 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1604681595
transform 1 0 4140 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1604681595
transform 1 0 3036 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1604681595
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_23
timestamp 1604681595
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_31
timestamp 1604681595
transform 1 0 3956 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_35
timestamp 1604681595
transform 1 0 4324 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_43
timestamp 1604681595
transform 1 0 5060 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1604681595
transform 1 0 5244 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_47
timestamp 1604681595
transform 1 0 5428 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_52
timestamp 1604681595
transform 1 0 5888 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 5704 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604681595
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8464 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6900 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8280 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_72
timestamp 1604681595
transform 1 0 7728 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_76
timestamp 1604681595
transform 1 0 8096 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 10028 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9476 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10488 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604681595
transform 1 0 9844 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_89
timestamp 1604681595
transform 1 0 9292 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_93
timestamp 1604681595
transform 1 0 9660 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_100
timestamp 1604681595
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_104
timestamp 1604681595
transform 1 0 10672 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10856 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1604681595
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12972 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14352 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_138
timestamp 1604681595
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_142
timestamp 1604681595
transform 1 0 14168 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604681595
transform 1 0 14628 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15732 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15180 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_146
timestamp 1604681595
transform 1 0 14536 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_151
timestamp 1604681595
transform 1 0 14996 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_155
timestamp 1604681595
transform 1 0 15364 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_176
timestamp 1604681595
transform 1 0 17296 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_172
timestamp 1604681595
transform 1 0 16928 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_168
timestamp 1604681595
transform 1 0 16560 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16744 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_179
timestamp 1604681595
transform 1 0 17572 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18124 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19964 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19780 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_194
timestamp 1604681595
transform 1 0 18952 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_198
timestamp 1604681595
transform 1 0 19320 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_202
timestamp 1604681595
transform 1 0 19688 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22172 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20976 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21988 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_214
timestamp 1604681595
transform 1 0 20792 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_218
timestamp 1604681595
transform 1 0 21160 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_222
timestamp 1604681595
transform 1 0 21528 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_226
timestamp 1604681595
transform 1 0 21896 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22908 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_235
timestamp 1604681595
transform 1 0 22724 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1604681595
transform 1 0 23092 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1604681595
transform 1 0 23460 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 24564 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_259
timestamp 1604681595
transform 1 0 24932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_263
timestamp 1604681595
transform 1 0 25300 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_275
timestamp 1604681595
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_7
timestamp 1604681595
transform 1 0 1748 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_19
timestamp 1604681595
transform 1 0 2852 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_36
timestamp 1604681595
transform 1 0 4416 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 5704 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_48
timestamp 1604681595
transform 1 0 5520 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_54
timestamp 1604681595
transform 1 0 6072 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_58
timestamp 1604681595
transform 1 0 6440 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 7452 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 8556 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7084 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_67
timestamp 1604681595
transform 1 0 7268 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_73
timestamp 1604681595
transform 1 0 7820 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_77
timestamp 1604681595
transform 1 0 8188 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 10304 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9936 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1604681595
transform 1 0 8924 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_89
timestamp 1604681595
transform 1 0 9292 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_98
timestamp 1604681595
transform 1 0 10120 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_104
timestamp 1604681595
transform 1 0 10672 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 11408 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_116
timestamp 1604681595
transform 1 0 11776 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_120
timestamp 1604681595
transform 1 0 12144 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 14260 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 13616 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13984 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_134
timestamp 1604681595
transform 1 0 13432 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1604681595
transform 1 0 13800 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_142
timestamp 1604681595
transform 1 0 14168 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15640 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_147
timestamp 1604681595
transform 1 0 14628 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_151
timestamp 1604681595
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_167
timestamp 1604681595
transform 1 0 16468 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16652 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_171
timestamp 1604681595
transform 1 0 16836 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17020 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_178
timestamp 1604681595
transform 1 0 17480 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 17204 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_182
timestamp 1604681595
transform 1 0 17848 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 20056 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18492 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 19504 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_198
timestamp 1604681595
transform 1 0 19320 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_202
timestamp 1604681595
transform 1 0 19688 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_209
timestamp 1604681595
transform 1 0 20332 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_224
timestamp 1604681595
transform 1 0 21712 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22448 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_238
timestamp 1604681595
transform 1 0 23000 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_246
timestamp 1604681595
transform 1 0 23736 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 24564 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_259
timestamp 1604681595
transform 1 0 24932 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_271
timestamp 1604681595
transform 1 0 26036 0 -1 25568
box -38 -48 590 592
<< labels >>
rlabel metal2 s 19522 0 19578 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 294 27520 350 28000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 25134 0 25190 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 27618 27520 27674 28000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 8298 0 8354 480 6 ccff_head
port 4 nsew default input
rlabel metal2 s 13910 0 13966 480 6 ccff_tail
port 5 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 6 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[10]
port 7 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[11]
port 8 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[12]
port 9 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[13]
port 10 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chanx_left_in[14]
port 11 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[15]
port 12 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[16]
port 13 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[17]
port 14 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[18]
port 15 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[19]
port 16 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[1]
port 17 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[2]
port 18 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[3]
port 19 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[4]
port 20 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[5]
port 21 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[6]
port 22 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[7]
port 23 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[8]
port 24 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[9]
port 25 nsew default input
rlabel metal3 s 0 16056 480 16176 6 chanx_left_out[0]
port 26 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chanx_left_out[10]
port 27 nsew default tristate
rlabel metal3 s 0 22720 480 22840 6 chanx_left_out[11]
port 28 nsew default tristate
rlabel metal3 s 0 23400 480 23520 6 chanx_left_out[12]
port 29 nsew default tristate
rlabel metal3 s 0 23944 480 24064 6 chanx_left_out[13]
port 30 nsew default tristate
rlabel metal3 s 0 24624 480 24744 6 chanx_left_out[14]
port 31 nsew default tristate
rlabel metal3 s 0 25168 480 25288 6 chanx_left_out[15]
port 32 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[16]
port 33 nsew default tristate
rlabel metal3 s 0 26392 480 26512 6 chanx_left_out[17]
port 34 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[18]
port 35 nsew default tristate
rlabel metal3 s 0 27616 480 27736 6 chanx_left_out[19]
port 36 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[1]
port 37 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[2]
port 38 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[4]
port 40 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[5]
port 41 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[6]
port 42 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[7]
port 43 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 chanx_left_out[8]
port 44 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[9]
port 45 nsew default tristate
rlabel metal3 s 27520 3816 28000 3936 6 chanx_right_in[0]
port 46 nsew default input
rlabel metal3 s 27520 9936 28000 10056 6 chanx_right_in[10]
port 47 nsew default input
rlabel metal3 s 27520 10616 28000 10736 6 chanx_right_in[11]
port 48 nsew default input
rlabel metal3 s 27520 11160 28000 11280 6 chanx_right_in[12]
port 49 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_in[13]
port 50 nsew default input
rlabel metal3 s 27520 12384 28000 12504 6 chanx_right_in[14]
port 51 nsew default input
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_in[15]
port 52 nsew default input
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_in[16]
port 53 nsew default input
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_in[17]
port 54 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[18]
port 55 nsew default input
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_in[19]
port 56 nsew default input
rlabel metal3 s 27520 4496 28000 4616 6 chanx_right_in[1]
port 57 nsew default input
rlabel metal3 s 27520 5040 28000 5160 6 chanx_right_in[2]
port 58 nsew default input
rlabel metal3 s 27520 5720 28000 5840 6 chanx_right_in[3]
port 59 nsew default input
rlabel metal3 s 27520 6264 28000 6384 6 chanx_right_in[4]
port 60 nsew default input
rlabel metal3 s 27520 6944 28000 7064 6 chanx_right_in[5]
port 61 nsew default input
rlabel metal3 s 27520 7488 28000 7608 6 chanx_right_in[6]
port 62 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_in[7]
port 63 nsew default input
rlabel metal3 s 27520 8712 28000 8832 6 chanx_right_in[8]
port 64 nsew default input
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_in[9]
port 65 nsew default input
rlabel metal3 s 27520 16056 28000 16176 6 chanx_right_out[0]
port 66 nsew default tristate
rlabel metal3 s 27520 22176 28000 22296 6 chanx_right_out[10]
port 67 nsew default tristate
rlabel metal3 s 27520 22720 28000 22840 6 chanx_right_out[11]
port 68 nsew default tristate
rlabel metal3 s 27520 23400 28000 23520 6 chanx_right_out[12]
port 69 nsew default tristate
rlabel metal3 s 27520 23944 28000 24064 6 chanx_right_out[13]
port 70 nsew default tristate
rlabel metal3 s 27520 24624 28000 24744 6 chanx_right_out[14]
port 71 nsew default tristate
rlabel metal3 s 27520 25168 28000 25288 6 chanx_right_out[15]
port 72 nsew default tristate
rlabel metal3 s 27520 25848 28000 25968 6 chanx_right_out[16]
port 73 nsew default tristate
rlabel metal3 s 27520 26392 28000 26512 6 chanx_right_out[17]
port 74 nsew default tristate
rlabel metal3 s 27520 27072 28000 27192 6 chanx_right_out[18]
port 75 nsew default tristate
rlabel metal3 s 27520 27616 28000 27736 6 chanx_right_out[19]
port 76 nsew default tristate
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_out[1]
port 77 nsew default tristate
rlabel metal3 s 27520 17280 28000 17400 6 chanx_right_out[2]
port 78 nsew default tristate
rlabel metal3 s 27520 17824 28000 17944 6 chanx_right_out[3]
port 79 nsew default tristate
rlabel metal3 s 27520 18504 28000 18624 6 chanx_right_out[4]
port 80 nsew default tristate
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[5]
port 81 nsew default tristate
rlabel metal3 s 27520 19728 28000 19848 6 chanx_right_out[6]
port 82 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_out[7]
port 83 nsew default tristate
rlabel metal3 s 27520 20952 28000 21072 6 chanx_right_out[8]
port 84 nsew default tristate
rlabel metal3 s 27520 21496 28000 21616 6 chanx_right_out[9]
port 85 nsew default tristate
rlabel metal2 s 5262 27520 5318 28000 6 chany_top_in[0]
port 86 nsew default input
rlabel metal2 s 10874 27520 10930 28000 6 chany_top_in[10]
port 87 nsew default input
rlabel metal2 s 11426 27520 11482 28000 6 chany_top_in[11]
port 88 nsew default input
rlabel metal2 s 11978 27520 12034 28000 6 chany_top_in[12]
port 89 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[13]
port 90 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 chany_top_in[14]
port 91 nsew default input
rlabel metal2 s 13634 27520 13690 28000 6 chany_top_in[15]
port 92 nsew default input
rlabel metal2 s 14278 27520 14334 28000 6 chany_top_in[16]
port 93 nsew default input
rlabel metal2 s 14830 27520 14886 28000 6 chany_top_in[17]
port 94 nsew default input
rlabel metal2 s 15382 27520 15438 28000 6 chany_top_in[18]
port 95 nsew default input
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_in[19]
port 96 nsew default input
rlabel metal2 s 5814 27520 5870 28000 6 chany_top_in[1]
port 97 nsew default input
rlabel metal2 s 6366 27520 6422 28000 6 chany_top_in[2]
port 98 nsew default input
rlabel metal2 s 6918 27520 6974 28000 6 chany_top_in[3]
port 99 nsew default input
rlabel metal2 s 7562 27520 7618 28000 6 chany_top_in[4]
port 100 nsew default input
rlabel metal2 s 8114 27520 8170 28000 6 chany_top_in[5]
port 101 nsew default input
rlabel metal2 s 8666 27520 8722 28000 6 chany_top_in[6]
port 102 nsew default input
rlabel metal2 s 9218 27520 9274 28000 6 chany_top_in[7]
port 103 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[8]
port 104 nsew default input
rlabel metal2 s 10322 27520 10378 28000 6 chany_top_in[9]
port 105 nsew default input
rlabel metal2 s 16486 27520 16542 28000 6 chany_top_out[0]
port 106 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[10]
port 107 nsew default tristate
rlabel metal2 s 22650 27520 22706 28000 6 chany_top_out[11]
port 108 nsew default tristate
rlabel metal2 s 23202 27520 23258 28000 6 chany_top_out[12]
port 109 nsew default tristate
rlabel metal2 s 23754 27520 23810 28000 6 chany_top_out[13]
port 110 nsew default tristate
rlabel metal2 s 24306 27520 24362 28000 6 chany_top_out[14]
port 111 nsew default tristate
rlabel metal2 s 24858 27520 24914 28000 6 chany_top_out[15]
port 112 nsew default tristate
rlabel metal2 s 25410 27520 25466 28000 6 chany_top_out[16]
port 113 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[17]
port 114 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[18]
port 115 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[19]
port 116 nsew default tristate
rlabel metal2 s 17038 27520 17094 28000 6 chany_top_out[1]
port 117 nsew default tristate
rlabel metal2 s 17590 27520 17646 28000 6 chany_top_out[2]
port 118 nsew default tristate
rlabel metal2 s 18142 27520 18198 28000 6 chany_top_out[3]
port 119 nsew default tristate
rlabel metal2 s 18694 27520 18750 28000 6 chany_top_out[4]
port 120 nsew default tristate
rlabel metal2 s 19246 27520 19302 28000 6 chany_top_out[5]
port 121 nsew default tristate
rlabel metal2 s 19798 27520 19854 28000 6 chany_top_out[6]
port 122 nsew default tristate
rlabel metal2 s 20350 27520 20406 28000 6 chany_top_out[7]
port 123 nsew default tristate
rlabel metal2 s 20902 27520 20958 28000 6 chany_top_out[8]
port 124 nsew default tristate
rlabel metal2 s 21546 27520 21602 28000 6 chany_top_out[9]
port 125 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 left_bottom_grid_pin_11_
port 126 nsew default input
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_1_
port 127 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_3_
port 128 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_5_
port 129 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_7_
port 130 nsew default input
rlabel metal3 s 0 2592 480 2712 6 left_bottom_grid_pin_9_
port 131 nsew default input
rlabel metal2 s 2778 0 2834 480 6 prog_clk
port 132 nsew default input
rlabel metal3 s 27520 3272 28000 3392 6 right_bottom_grid_pin_11_
port 133 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_1_
port 134 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_bottom_grid_pin_3_
port 135 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_5_
port 136 nsew default input
rlabel metal3 s 27520 2048 28000 2168 6 right_bottom_grid_pin_7_
port 137 nsew default input
rlabel metal3 s 27520 2592 28000 2712 6 right_bottom_grid_pin_9_
port 138 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_42_
port 139 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_43_
port 140 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_44_
port 141 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_45_
port 142 nsew default input
rlabel metal2 s 3054 27520 3110 28000 6 top_left_grid_pin_46_
port 143 nsew default input
rlabel metal2 s 3606 27520 3662 28000 6 top_left_grid_pin_47_
port 144 nsew default input
rlabel metal2 s 4158 27520 4214 28000 6 top_left_grid_pin_48_
port 145 nsew default input
rlabel metal2 s 4710 27520 4766 28000 6 top_left_grid_pin_49_
port 146 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 147 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 148 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
