magic
tech EFS8A
magscale 1 2
timestamp 1604399188
<< viali >>
rect 1857 23137 1891 23171
rect 2041 23001 2075 23035
rect 2501 22525 2535 22559
rect 3053 22525 3087 22559
rect 1857 22389 1891 22423
rect 2685 22389 2719 22423
rect 3789 22049 3823 22083
rect 3973 21913 4007 21947
rect 4065 21641 4099 21675
rect 4433 21505 4467 21539
rect 3881 21437 3915 21471
rect 3789 21301 3823 21335
rect 5445 20009 5479 20043
rect 5261 19873 5295 19907
rect 6549 19261 6583 19295
rect 7101 19261 7135 19295
rect 5261 19125 5295 19159
rect 6733 19125 6767 19159
rect 6825 18921 6859 18955
rect 6641 18785 6675 18819
rect 6733 18037 6767 18071
rect 10689 17833 10723 17867
rect 7285 17697 7319 17731
rect 10505 17697 10539 17731
rect 7469 17561 7503 17595
rect 7929 17085 7963 17119
rect 7285 16949 7319 16983
rect 8113 16949 8147 16983
rect 8481 16949 8515 16983
rect 10505 16949 10539 16983
rect 9585 16745 9619 16779
rect 9401 16609 9435 16643
rect 9493 16201 9527 16235
rect 13633 16201 13667 16235
rect 9309 15997 9343 16031
rect 13449 15997 13483 16031
rect 9217 15861 9251 15895
rect 9861 15861 9895 15895
rect 14001 15861 14035 15895
rect 10873 15113 10907 15147
rect 17957 15113 17991 15147
rect 19429 15113 19463 15147
rect 16301 15045 16335 15079
rect 10689 14909 10723 14943
rect 16117 14909 16151 14943
rect 17773 14909 17807 14943
rect 18325 14909 18359 14943
rect 19245 14909 19279 14943
rect 19797 14909 19831 14943
rect 16577 14841 16611 14875
rect 11241 14773 11275 14807
rect 11241 14569 11275 14603
rect 15657 14569 15691 14603
rect 17773 14569 17807 14603
rect 19521 14569 19555 14603
rect 24489 14569 24523 14603
rect 12704 14501 12738 14535
rect 11057 14433 11091 14467
rect 16025 14433 16059 14467
rect 18141 14433 18175 14467
rect 19337 14433 19371 14467
rect 24305 14433 24339 14467
rect 12437 14365 12471 14399
rect 16117 14365 16151 14399
rect 16209 14365 16243 14399
rect 17681 14365 17715 14399
rect 18233 14365 18267 14399
rect 18417 14365 18451 14399
rect 13817 14229 13851 14263
rect 18785 14229 18819 14263
rect 12529 14025 12563 14059
rect 17589 14025 17623 14059
rect 16577 13889 16611 13923
rect 18233 13889 18267 13923
rect 18417 13889 18451 13923
rect 11057 13821 11091 13855
rect 14093 13821 14127 13855
rect 14277 13821 14311 13855
rect 16301 13821 16335 13855
rect 17221 13821 17255 13855
rect 12805 13753 12839 13787
rect 13817 13753 13851 13787
rect 14544 13753 14578 13787
rect 18662 13753 18696 13787
rect 15657 13685 15691 13719
rect 19797 13685 19831 13719
rect 24305 13685 24339 13719
rect 13817 13481 13851 13515
rect 14829 13481 14863 13515
rect 16117 13481 16151 13515
rect 18785 13481 18819 13515
rect 19337 13481 19371 13515
rect 23385 13481 23419 13515
rect 12437 13345 12471 13379
rect 12704 13345 12738 13379
rect 15381 13345 15415 13379
rect 17672 13345 17706 13379
rect 23201 13345 23235 13379
rect 14461 13277 14495 13311
rect 15473 13277 15507 13311
rect 15657 13277 15691 13311
rect 17405 13277 17439 13311
rect 20625 13277 20659 13311
rect 15013 13209 15047 13243
rect 13081 12937 13115 12971
rect 13633 12937 13667 12971
rect 14737 12937 14771 12971
rect 16577 12937 16611 12971
rect 18325 12937 18359 12971
rect 19061 12937 19095 12971
rect 15013 12869 15047 12903
rect 14185 12801 14219 12835
rect 15197 12801 15231 12835
rect 17865 12801 17899 12835
rect 19245 12801 19279 12835
rect 12161 12733 12195 12767
rect 12713 12733 12747 12767
rect 17405 12733 17439 12767
rect 19512 12733 19546 12767
rect 23569 12733 23603 12767
rect 13541 12665 13575 12699
rect 14001 12665 14035 12699
rect 15464 12665 15498 12699
rect 18785 12665 18819 12699
rect 12345 12597 12379 12631
rect 14093 12597 14127 12631
rect 20625 12597 20659 12631
rect 12529 12393 12563 12427
rect 14093 12393 14127 12427
rect 14369 12393 14403 12427
rect 15381 12393 15415 12427
rect 15749 12393 15783 12427
rect 17681 12393 17715 12427
rect 18877 12393 18911 12427
rect 19337 12393 19371 12427
rect 20993 12393 21027 12427
rect 14829 12325 14863 12359
rect 21085 12325 21119 12359
rect 13909 12257 13943 12291
rect 15197 12257 15231 12291
rect 16301 12257 16335 12291
rect 16568 12257 16602 12291
rect 19245 12257 19279 12291
rect 19521 12189 19555 12223
rect 21177 12189 21211 12223
rect 20625 12121 20659 12155
rect 13725 12053 13759 12087
rect 14277 11849 14311 11883
rect 15749 11849 15783 11883
rect 17129 11849 17163 11883
rect 17773 11849 17807 11883
rect 21361 11849 21395 11883
rect 22097 11849 22131 11883
rect 14737 11781 14771 11815
rect 16853 11781 16887 11815
rect 21729 11781 21763 11815
rect 13725 11713 13759 11747
rect 15381 11713 15415 11747
rect 16301 11713 16335 11747
rect 18325 11713 18359 11747
rect 18233 11645 18267 11679
rect 19429 11645 19463 11679
rect 24305 11645 24339 11679
rect 24857 11645 24891 11679
rect 15105 11577 15139 11611
rect 18141 11577 18175 11611
rect 19696 11577 19730 11611
rect 14553 11509 14587 11543
rect 15197 11509 15231 11543
rect 17497 11509 17531 11543
rect 18877 11509 18911 11543
rect 19337 11509 19371 11543
rect 20809 11509 20843 11543
rect 24489 11509 24523 11543
rect 18233 11305 18267 11339
rect 18877 11305 18911 11339
rect 19429 11305 19463 11339
rect 19797 11305 19831 11339
rect 14829 11237 14863 11271
rect 17865 11237 17899 11271
rect 20441 11237 20475 11271
rect 20892 11237 20926 11271
rect 18969 11101 19003 11135
rect 20625 11101 20659 11135
rect 22005 10965 22039 10999
rect 21085 10625 21119 10659
rect 22189 10625 22223 10659
rect 14645 10557 14679 10591
rect 19061 10557 19095 10591
rect 19328 10557 19362 10591
rect 21361 10557 21395 10591
rect 21913 10557 21947 10591
rect 22005 10557 22039 10591
rect 15289 10489 15323 10523
rect 18601 10489 18635 10523
rect 14829 10421 14863 10455
rect 18877 10421 18911 10455
rect 20441 10421 20475 10455
rect 21545 10421 21579 10455
rect 21085 10217 21119 10251
rect 21729 10217 21763 10251
rect 18417 10149 18451 10183
rect 19337 10149 19371 10183
rect 19245 10081 19279 10115
rect 20993 10081 21027 10115
rect 19521 10013 19555 10047
rect 21177 10013 21211 10047
rect 18785 9945 18819 9979
rect 18877 9877 18911 9911
rect 20349 9877 20383 9911
rect 20625 9877 20659 9911
rect 18049 9673 18083 9707
rect 21177 9673 21211 9707
rect 18417 9605 18451 9639
rect 14921 9537 14955 9571
rect 14369 9469 14403 9503
rect 18877 9469 18911 9503
rect 19122 9401 19156 9435
rect 14553 9333 14587 9367
rect 18785 9333 18819 9367
rect 20257 9333 20291 9367
rect 20901 9333 20935 9367
rect 18877 9129 18911 9163
rect 19521 9129 19555 9163
rect 20809 9129 20843 9163
rect 15933 8993 15967 9027
rect 18785 8993 18819 9027
rect 19061 8925 19095 8959
rect 16117 8789 16151 8823
rect 18417 8789 18451 8823
rect 14461 8585 14495 8619
rect 18693 8585 18727 8619
rect 14001 8517 14035 8551
rect 16025 8517 16059 8551
rect 18141 8449 18175 8483
rect 13817 8381 13851 8415
rect 19153 8381 19187 8415
rect 19420 8381 19454 8415
rect 18049 8313 18083 8347
rect 19061 8245 19095 8279
rect 20533 8245 20567 8279
rect 18509 8041 18543 8075
rect 16669 7905 16703 7939
rect 20993 7905 21027 7939
rect 19245 7837 19279 7871
rect 21085 7837 21119 7871
rect 21269 7837 21303 7871
rect 16853 7701 16887 7735
rect 20625 7701 20659 7735
rect 16393 7497 16427 7531
rect 16761 7497 16795 7531
rect 18417 7497 18451 7531
rect 22005 7497 22039 7531
rect 22281 7429 22315 7463
rect 19153 7361 19187 7395
rect 15749 7293 15783 7327
rect 17773 7293 17807 7327
rect 19613 7293 19647 7327
rect 19880 7293 19914 7327
rect 15933 7157 15967 7191
rect 17957 7157 17991 7191
rect 19521 7157 19555 7191
rect 20993 7157 21027 7191
rect 21545 7157 21579 7191
rect 19337 6953 19371 6987
rect 22281 6953 22315 6987
rect 17865 6817 17899 6851
rect 21168 6817 21202 6851
rect 19429 6749 19463 6783
rect 19521 6749 19555 6783
rect 20901 6749 20935 6783
rect 20165 6681 20199 6715
rect 18049 6613 18083 6647
rect 18969 6613 19003 6647
rect 17957 6409 17991 6443
rect 18509 6409 18543 6443
rect 19521 6409 19555 6443
rect 19981 6409 20015 6443
rect 19245 6273 19279 6307
rect 20165 6273 20199 6307
rect 18601 6205 18635 6239
rect 20432 6205 20466 6239
rect 18785 6069 18819 6103
rect 21545 6069 21579 6103
rect 22189 6069 22223 6103
rect 18233 5865 18267 5899
rect 19061 5865 19095 5899
rect 20165 5865 20199 5899
rect 16945 5729 16979 5763
rect 18049 5729 18083 5763
rect 19337 5729 19371 5763
rect 21361 5729 21395 5763
rect 21453 5661 21487 5695
rect 21637 5661 21671 5695
rect 17129 5525 17163 5559
rect 19521 5525 19555 5559
rect 20993 5525 21027 5559
rect 16945 5321 16979 5355
rect 18141 5321 18175 5355
rect 19429 5321 19463 5355
rect 22281 5321 22315 5355
rect 21729 5185 21763 5219
rect 21913 5185 21947 5219
rect 20257 5049 20291 5083
rect 21637 5049 21671 5083
rect 20165 4981 20199 5015
rect 20993 4981 21027 5015
rect 21269 4981 21303 5015
rect 21637 4777 21671 4811
rect 22005 4777 22039 4811
rect 21361 4709 21395 4743
rect 20717 4641 20751 4675
rect 24305 4641 24339 4675
rect 20901 4505 20935 4539
rect 24489 4437 24523 4471
rect 20625 4233 20659 4267
rect 24213 4233 24247 4267
rect 21361 4097 21395 4131
rect 20717 4029 20751 4063
rect 21821 4029 21855 4063
rect 22373 4029 22407 4063
rect 24305 4029 24339 4063
rect 24857 4029 24891 4063
rect 20901 3893 20935 3927
rect 22005 3893 22039 3927
rect 24489 3893 24523 3927
rect 24305 3553 24339 3587
rect 23661 3349 23695 3383
rect 24489 3349 24523 3383
rect 24397 3145 24431 3179
rect 23661 2941 23695 2975
rect 24765 2941 24799 2975
rect 23845 2805 23879 2839
rect 24949 2805 24983 2839
rect 25317 2805 25351 2839
rect 21545 2601 21579 2635
rect 22741 2601 22775 2635
rect 24857 2601 24891 2635
rect 20901 2465 20935 2499
rect 22557 2465 22591 2499
rect 24305 2465 24339 2499
rect 23201 2397 23235 2431
rect 21085 2261 21119 2295
rect 24489 2261 24523 2295
<< metal1 >>
rect 19230 26324 19236 26376
rect 19288 26364 19294 26376
rect 23830 26364 23836 26376
rect 19288 26336 23836 26364
rect 19288 26324 19294 26336
rect 23830 26324 23836 26336
rect 23888 26324 23894 26376
rect 13710 26256 13716 26308
rect 13768 26296 13774 26308
rect 24474 26296 24480 26308
rect 13768 26268 24480 26296
rect 13768 26256 13774 26268
rect 24474 26256 24480 26268
rect 24532 26256 24538 26308
rect 816 25594 26576 25616
rect 816 25542 10027 25594
rect 10079 25542 10091 25594
rect 10143 25542 10155 25594
rect 10207 25542 10219 25594
rect 10271 25542 19360 25594
rect 19412 25542 19424 25594
rect 19476 25542 19488 25594
rect 19540 25542 19552 25594
rect 19604 25542 26576 25594
rect 816 25520 26576 25542
rect 816 25050 26576 25072
rect 816 24998 5360 25050
rect 5412 24998 5424 25050
rect 5476 24998 5488 25050
rect 5540 24998 5552 25050
rect 5604 24998 14694 25050
rect 14746 24998 14758 25050
rect 14810 24998 14822 25050
rect 14874 24998 14886 25050
rect 14938 24998 24027 25050
rect 24079 24998 24091 25050
rect 24143 24998 24155 25050
rect 24207 24998 24219 25050
rect 24271 24998 26576 25050
rect 816 24976 26576 24998
rect 11226 24896 11232 24948
rect 11284 24936 11290 24948
rect 23830 24936 23836 24948
rect 11284 24908 23836 24936
rect 11284 24896 11290 24908
rect 23830 24896 23836 24908
rect 23888 24896 23894 24948
rect 10674 24828 10680 24880
rect 10732 24868 10738 24880
rect 24474 24868 24480 24880
rect 10732 24840 24480 24868
rect 10732 24828 10738 24840
rect 24474 24828 24480 24840
rect 24532 24828 24538 24880
rect 816 24506 26576 24528
rect 816 24454 10027 24506
rect 10079 24454 10091 24506
rect 10143 24454 10155 24506
rect 10207 24454 10219 24506
rect 10271 24454 19360 24506
rect 19412 24454 19424 24506
rect 19476 24454 19488 24506
rect 19540 24454 19552 24506
rect 19604 24454 26576 24506
rect 816 24432 26576 24454
rect 816 23962 26576 23984
rect 816 23910 5360 23962
rect 5412 23910 5424 23962
rect 5476 23910 5488 23962
rect 5540 23910 5552 23962
rect 5604 23910 14694 23962
rect 14746 23910 14758 23962
rect 14810 23910 14822 23962
rect 14874 23910 14886 23962
rect 14938 23910 24027 23962
rect 24079 23910 24091 23962
rect 24143 23910 24155 23962
rect 24207 23910 24219 23962
rect 24271 23910 26576 23962
rect 816 23888 26576 23910
rect 816 23418 26576 23440
rect 816 23366 10027 23418
rect 10079 23366 10091 23418
rect 10143 23366 10155 23418
rect 10207 23366 10219 23418
rect 10271 23366 19360 23418
rect 19412 23366 19424 23418
rect 19476 23366 19488 23418
rect 19540 23366 19552 23418
rect 19604 23366 26576 23418
rect 816 23344 26576 23366
rect 1842 23168 1848 23180
rect 1803 23140 1848 23168
rect 1842 23128 1848 23140
rect 1900 23128 1906 23180
rect 2026 23032 2032 23044
rect 1987 23004 2032 23032
rect 2026 22992 2032 23004
rect 2084 22992 2090 23044
rect 14446 22924 14452 22976
rect 14504 22964 14510 22976
rect 15090 22964 15096 22976
rect 14504 22936 15096 22964
rect 14504 22924 14510 22936
rect 15090 22924 15096 22936
rect 15148 22924 15154 22976
rect 816 22874 26576 22896
rect 816 22822 5360 22874
rect 5412 22822 5424 22874
rect 5476 22822 5488 22874
rect 5540 22822 5552 22874
rect 5604 22822 14694 22874
rect 14746 22822 14758 22874
rect 14810 22822 14822 22874
rect 14874 22822 14886 22874
rect 14938 22822 24027 22874
rect 24079 22822 24091 22874
rect 24143 22822 24155 22874
rect 24207 22822 24219 22874
rect 24271 22822 26576 22874
rect 816 22800 26576 22822
rect 2486 22516 2492 22568
rect 2544 22556 2550 22568
rect 3041 22559 3099 22565
rect 3041 22556 3053 22559
rect 2544 22528 3053 22556
rect 2544 22516 2550 22528
rect 3041 22525 3053 22528
rect 3087 22525 3099 22559
rect 3041 22519 3099 22525
rect 1842 22420 1848 22432
rect 1803 22392 1848 22420
rect 1842 22380 1848 22392
rect 1900 22380 1906 22432
rect 2670 22420 2676 22432
rect 2631 22392 2676 22420
rect 2670 22380 2676 22392
rect 2728 22380 2734 22432
rect 816 22330 26576 22352
rect 816 22278 10027 22330
rect 10079 22278 10091 22330
rect 10143 22278 10155 22330
rect 10207 22278 10219 22330
rect 10271 22278 19360 22330
rect 19412 22278 19424 22330
rect 19476 22278 19488 22330
rect 19540 22278 19552 22330
rect 19604 22278 26576 22330
rect 816 22256 26576 22278
rect 3774 22080 3780 22092
rect 3735 22052 3780 22080
rect 3774 22040 3780 22052
rect 3832 22040 3838 22092
rect 3958 21944 3964 21956
rect 3919 21916 3964 21944
rect 3958 21904 3964 21916
rect 4016 21904 4022 21956
rect 816 21786 26576 21808
rect 816 21734 5360 21786
rect 5412 21734 5424 21786
rect 5476 21734 5488 21786
rect 5540 21734 5552 21786
rect 5604 21734 14694 21786
rect 14746 21734 14758 21786
rect 14810 21734 14822 21786
rect 14874 21734 14886 21786
rect 14938 21734 24027 21786
rect 24079 21734 24091 21786
rect 24143 21734 24155 21786
rect 24207 21734 24219 21786
rect 24271 21734 26576 21786
rect 816 21712 26576 21734
rect 4050 21672 4056 21684
rect 4011 21644 4056 21672
rect 4050 21632 4056 21644
rect 4108 21632 4114 21684
rect 3774 21496 3780 21548
rect 3832 21536 3838 21548
rect 4421 21539 4479 21545
rect 4421 21536 4433 21539
rect 3832 21508 4433 21536
rect 3832 21496 3838 21508
rect 4421 21505 4433 21508
rect 4467 21505 4479 21539
rect 4421 21499 4479 21505
rect 3869 21471 3927 21477
rect 3869 21437 3881 21471
rect 3915 21437 3927 21471
rect 3869 21431 3927 21437
rect 3884 21344 3912 21431
rect 3777 21335 3835 21341
rect 3777 21301 3789 21335
rect 3823 21332 3835 21335
rect 3866 21332 3872 21344
rect 3823 21304 3872 21332
rect 3823 21301 3835 21304
rect 3777 21295 3835 21301
rect 3866 21292 3872 21304
rect 3924 21292 3930 21344
rect 816 21242 26576 21264
rect 816 21190 10027 21242
rect 10079 21190 10091 21242
rect 10143 21190 10155 21242
rect 10207 21190 10219 21242
rect 10271 21190 19360 21242
rect 19412 21190 19424 21242
rect 19476 21190 19488 21242
rect 19540 21190 19552 21242
rect 19604 21190 26576 21242
rect 816 21168 26576 21190
rect 816 20698 26576 20720
rect 816 20646 5360 20698
rect 5412 20646 5424 20698
rect 5476 20646 5488 20698
rect 5540 20646 5552 20698
rect 5604 20646 14694 20698
rect 14746 20646 14758 20698
rect 14810 20646 14822 20698
rect 14874 20646 14886 20698
rect 14938 20646 24027 20698
rect 24079 20646 24091 20698
rect 24143 20646 24155 20698
rect 24207 20646 24219 20698
rect 24271 20646 26576 20698
rect 816 20624 26576 20646
rect 816 20154 26576 20176
rect 816 20102 10027 20154
rect 10079 20102 10091 20154
rect 10143 20102 10155 20154
rect 10207 20102 10219 20154
rect 10271 20102 19360 20154
rect 19412 20102 19424 20154
rect 19476 20102 19488 20154
rect 19540 20102 19552 20154
rect 19604 20102 26576 20154
rect 816 20080 26576 20102
rect 5433 20043 5491 20049
rect 5433 20009 5445 20043
rect 5479 20040 5491 20043
rect 5706 20040 5712 20052
rect 5479 20012 5712 20040
rect 5479 20009 5491 20012
rect 5433 20003 5491 20009
rect 5706 20000 5712 20012
rect 5764 20000 5770 20052
rect 5246 19904 5252 19916
rect 5207 19876 5252 19904
rect 5246 19864 5252 19876
rect 5304 19864 5310 19916
rect 816 19610 26576 19632
rect 816 19558 5360 19610
rect 5412 19558 5424 19610
rect 5476 19558 5488 19610
rect 5540 19558 5552 19610
rect 5604 19558 14694 19610
rect 14746 19558 14758 19610
rect 14810 19558 14822 19610
rect 14874 19558 14886 19610
rect 14938 19558 24027 19610
rect 24079 19558 24091 19610
rect 24143 19558 24155 19610
rect 24207 19558 24219 19610
rect 24271 19558 26576 19610
rect 816 19536 26576 19558
rect 6534 19292 6540 19304
rect 6495 19264 6540 19292
rect 6534 19252 6540 19264
rect 6592 19292 6598 19304
rect 7089 19295 7147 19301
rect 7089 19292 7101 19295
rect 6592 19264 7101 19292
rect 6592 19252 6598 19264
rect 7089 19261 7101 19264
rect 7135 19261 7147 19295
rect 7089 19255 7147 19261
rect 21990 19252 21996 19304
rect 22048 19292 22054 19304
rect 22174 19292 22180 19304
rect 22048 19264 22180 19292
rect 22048 19252 22054 19264
rect 22174 19252 22180 19264
rect 22232 19252 22238 19304
rect 5246 19156 5252 19168
rect 5207 19128 5252 19156
rect 5246 19116 5252 19128
rect 5304 19116 5310 19168
rect 6718 19156 6724 19168
rect 6679 19128 6724 19156
rect 6718 19116 6724 19128
rect 6776 19116 6782 19168
rect 816 19066 26576 19088
rect 816 19014 10027 19066
rect 10079 19014 10091 19066
rect 10143 19014 10155 19066
rect 10207 19014 10219 19066
rect 10271 19014 19360 19066
rect 19412 19014 19424 19066
rect 19476 19014 19488 19066
rect 19540 19014 19552 19066
rect 19604 19014 26576 19066
rect 816 18992 26576 19014
rect 6810 18952 6816 18964
rect 6771 18924 6816 18952
rect 6810 18912 6816 18924
rect 6868 18912 6874 18964
rect 6629 18819 6687 18825
rect 6629 18785 6641 18819
rect 6675 18816 6687 18819
rect 6718 18816 6724 18828
rect 6675 18788 6724 18816
rect 6675 18785 6687 18788
rect 6629 18779 6687 18785
rect 6718 18776 6724 18788
rect 6776 18776 6782 18828
rect 816 18522 26576 18544
rect 816 18470 5360 18522
rect 5412 18470 5424 18522
rect 5476 18470 5488 18522
rect 5540 18470 5552 18522
rect 5604 18470 14694 18522
rect 14746 18470 14758 18522
rect 14810 18470 14822 18522
rect 14874 18470 14886 18522
rect 14938 18470 24027 18522
rect 24079 18470 24091 18522
rect 24143 18470 24155 18522
rect 24207 18470 24219 18522
rect 24271 18470 26576 18522
rect 816 18448 26576 18470
rect 6718 18068 6724 18080
rect 6679 18040 6724 18068
rect 6718 18028 6724 18040
rect 6776 18028 6782 18080
rect 816 17978 26576 18000
rect 816 17926 10027 17978
rect 10079 17926 10091 17978
rect 10143 17926 10155 17978
rect 10207 17926 10219 17978
rect 10271 17926 19360 17978
rect 19412 17926 19424 17978
rect 19476 17926 19488 17978
rect 19540 17926 19552 17978
rect 19604 17926 26576 17978
rect 816 17904 26576 17926
rect 10674 17864 10680 17876
rect 10635 17836 10680 17864
rect 10674 17824 10680 17836
rect 10732 17824 10738 17876
rect 7270 17728 7276 17740
rect 7231 17700 7276 17728
rect 7270 17688 7276 17700
rect 7328 17688 7334 17740
rect 10490 17728 10496 17740
rect 10451 17700 10496 17728
rect 10490 17688 10496 17700
rect 10548 17688 10554 17740
rect 7454 17592 7460 17604
rect 7415 17564 7460 17592
rect 7454 17552 7460 17564
rect 7512 17552 7518 17604
rect 816 17434 26576 17456
rect 816 17382 5360 17434
rect 5412 17382 5424 17434
rect 5476 17382 5488 17434
rect 5540 17382 5552 17434
rect 5604 17382 14694 17434
rect 14746 17382 14758 17434
rect 14810 17382 14822 17434
rect 14874 17382 14886 17434
rect 14938 17382 24027 17434
rect 24079 17382 24091 17434
rect 24143 17382 24155 17434
rect 24207 17382 24219 17434
rect 24271 17382 26576 17434
rect 816 17360 26576 17382
rect 7917 17119 7975 17125
rect 7917 17085 7929 17119
rect 7963 17116 7975 17119
rect 7963 17088 8512 17116
rect 7963 17085 7975 17088
rect 7917 17079 7975 17085
rect 8484 16992 8512 17088
rect 7270 16980 7276 16992
rect 7231 16952 7276 16980
rect 7270 16940 7276 16952
rect 7328 16940 7334 16992
rect 8098 16980 8104 16992
rect 8059 16952 8104 16980
rect 8098 16940 8104 16952
rect 8156 16940 8162 16992
rect 8466 16980 8472 16992
rect 8427 16952 8472 16980
rect 8466 16940 8472 16952
rect 8524 16940 8530 16992
rect 10490 16980 10496 16992
rect 10451 16952 10496 16980
rect 10490 16940 10496 16952
rect 10548 16940 10554 16992
rect 816 16890 26576 16912
rect 816 16838 10027 16890
rect 10079 16838 10091 16890
rect 10143 16838 10155 16890
rect 10207 16838 10219 16890
rect 10271 16838 19360 16890
rect 19412 16838 19424 16890
rect 19476 16838 19488 16890
rect 19540 16838 19552 16890
rect 19604 16838 26576 16890
rect 816 16816 26576 16838
rect 9570 16776 9576 16788
rect 9531 16748 9576 16776
rect 9570 16736 9576 16748
rect 9628 16736 9634 16788
rect 9389 16643 9447 16649
rect 9389 16609 9401 16643
rect 9435 16640 9447 16643
rect 9846 16640 9852 16652
rect 9435 16612 9852 16640
rect 9435 16609 9447 16612
rect 9389 16603 9447 16609
rect 9846 16600 9852 16612
rect 9904 16600 9910 16652
rect 816 16346 26576 16368
rect 816 16294 5360 16346
rect 5412 16294 5424 16346
rect 5476 16294 5488 16346
rect 5540 16294 5552 16346
rect 5604 16294 14694 16346
rect 14746 16294 14758 16346
rect 14810 16294 14822 16346
rect 14874 16294 14886 16346
rect 14938 16294 24027 16346
rect 24079 16294 24091 16346
rect 24143 16294 24155 16346
rect 24207 16294 24219 16346
rect 24271 16294 26576 16346
rect 816 16272 26576 16294
rect 9478 16232 9484 16244
rect 9439 16204 9484 16232
rect 9478 16192 9484 16204
rect 9536 16192 9542 16244
rect 13621 16235 13679 16241
rect 13621 16201 13633 16235
rect 13667 16232 13679 16235
rect 13710 16232 13716 16244
rect 13667 16204 13716 16232
rect 13667 16201 13679 16204
rect 13621 16195 13679 16201
rect 13710 16192 13716 16204
rect 13768 16192 13774 16244
rect 9297 16031 9355 16037
rect 9297 15997 9309 16031
rect 9343 15997 9355 16031
rect 9297 15991 9355 15997
rect 13437 16031 13495 16037
rect 13437 15997 13449 16031
rect 13483 16028 13495 16031
rect 13483 16000 13848 16028
rect 13483 15997 13495 16000
rect 13437 15991 13495 15997
rect 9312 15904 9340 15991
rect 13820 15904 13848 16000
rect 9205 15895 9263 15901
rect 9205 15861 9217 15895
rect 9251 15892 9263 15895
rect 9294 15892 9300 15904
rect 9251 15864 9300 15892
rect 9251 15861 9263 15864
rect 9205 15855 9263 15861
rect 9294 15852 9300 15864
rect 9352 15852 9358 15904
rect 9846 15892 9852 15904
rect 9807 15864 9852 15892
rect 9846 15852 9852 15864
rect 9904 15852 9910 15904
rect 13802 15852 13808 15904
rect 13860 15892 13866 15904
rect 13989 15895 14047 15901
rect 13989 15892 14001 15895
rect 13860 15864 14001 15892
rect 13860 15852 13866 15864
rect 13989 15861 14001 15864
rect 14035 15861 14047 15895
rect 13989 15855 14047 15861
rect 816 15802 26576 15824
rect 816 15750 10027 15802
rect 10079 15750 10091 15802
rect 10143 15750 10155 15802
rect 10207 15750 10219 15802
rect 10271 15750 19360 15802
rect 19412 15750 19424 15802
rect 19476 15750 19488 15802
rect 19540 15750 19552 15802
rect 19604 15750 26576 15802
rect 816 15728 26576 15750
rect 816 15258 26576 15280
rect 816 15206 5360 15258
rect 5412 15206 5424 15258
rect 5476 15206 5488 15258
rect 5540 15206 5552 15258
rect 5604 15206 14694 15258
rect 14746 15206 14758 15258
rect 14810 15206 14822 15258
rect 14874 15206 14886 15258
rect 14938 15206 24027 15258
rect 24079 15206 24091 15258
rect 24143 15206 24155 15258
rect 24207 15206 24219 15258
rect 24271 15206 26576 15258
rect 816 15184 26576 15206
rect 10858 15144 10864 15156
rect 10819 15116 10864 15144
rect 10858 15104 10864 15116
rect 10916 15104 10922 15156
rect 17942 15144 17948 15156
rect 17903 15116 17948 15144
rect 17942 15104 17948 15116
rect 18000 15104 18006 15156
rect 19417 15147 19475 15153
rect 19417 15113 19429 15147
rect 19463 15144 19475 15147
rect 19690 15144 19696 15156
rect 19463 15116 19696 15144
rect 19463 15113 19475 15116
rect 19417 15107 19475 15113
rect 19690 15104 19696 15116
rect 19748 15104 19754 15156
rect 16289 15079 16347 15085
rect 16289 15045 16301 15079
rect 16335 15045 16347 15079
rect 16289 15039 16347 15045
rect 10677 14943 10735 14949
rect 10677 14909 10689 14943
rect 10723 14940 10735 14943
rect 16105 14943 16163 14949
rect 10723 14912 11180 14940
rect 10723 14909 10735 14912
rect 10677 14903 10735 14909
rect 11152 14816 11180 14912
rect 16105 14909 16117 14943
rect 16151 14909 16163 14943
rect 16304 14940 16332 15039
rect 17761 14943 17819 14949
rect 17761 14940 17773 14943
rect 16304 14912 17773 14940
rect 16105 14903 16163 14909
rect 17761 14909 17773 14912
rect 17807 14940 17819 14943
rect 18313 14943 18371 14949
rect 18313 14940 18325 14943
rect 17807 14912 18325 14940
rect 17807 14909 17819 14912
rect 17761 14903 17819 14909
rect 18313 14909 18325 14912
rect 18359 14909 18371 14943
rect 18313 14903 18371 14909
rect 19233 14943 19291 14949
rect 19233 14909 19245 14943
rect 19279 14940 19291 14943
rect 19690 14940 19696 14952
rect 19279 14912 19696 14940
rect 19279 14909 19291 14912
rect 19233 14903 19291 14909
rect 15642 14832 15648 14884
rect 15700 14872 15706 14884
rect 16120 14872 16148 14903
rect 19690 14900 19696 14912
rect 19748 14940 19754 14952
rect 19785 14943 19843 14949
rect 19785 14940 19797 14943
rect 19748 14912 19797 14940
rect 19748 14900 19754 14912
rect 19785 14909 19797 14912
rect 19831 14909 19843 14943
rect 19785 14903 19843 14909
rect 16565 14875 16623 14881
rect 16565 14872 16577 14875
rect 15700 14844 16577 14872
rect 15700 14832 15706 14844
rect 16565 14841 16577 14844
rect 16611 14841 16623 14875
rect 16565 14835 16623 14841
rect 11134 14764 11140 14816
rect 11192 14804 11198 14816
rect 11229 14807 11287 14813
rect 11229 14804 11241 14807
rect 11192 14776 11241 14804
rect 11192 14764 11198 14776
rect 11229 14773 11241 14776
rect 11275 14773 11287 14807
rect 11229 14767 11287 14773
rect 816 14714 26576 14736
rect 816 14662 10027 14714
rect 10079 14662 10091 14714
rect 10143 14662 10155 14714
rect 10207 14662 10219 14714
rect 10271 14662 19360 14714
rect 19412 14662 19424 14714
rect 19476 14662 19488 14714
rect 19540 14662 19552 14714
rect 19604 14662 26576 14714
rect 816 14640 26576 14662
rect 11226 14600 11232 14612
rect 11187 14572 11232 14600
rect 11226 14560 11232 14572
rect 11284 14560 11290 14612
rect 15642 14600 15648 14612
rect 15603 14572 15648 14600
rect 15642 14560 15648 14572
rect 15700 14560 15706 14612
rect 17761 14603 17819 14609
rect 17761 14569 17773 14603
rect 17807 14569 17819 14603
rect 17761 14563 17819 14569
rect 19509 14603 19567 14609
rect 19509 14569 19521 14603
rect 19555 14600 19567 14603
rect 19690 14600 19696 14612
rect 19555 14572 19696 14600
rect 19555 14569 19567 14572
rect 19509 14563 19567 14569
rect 12514 14492 12520 14544
rect 12572 14532 12578 14544
rect 12692 14535 12750 14541
rect 12692 14532 12704 14535
rect 12572 14504 12704 14532
rect 12572 14492 12578 14504
rect 12692 14501 12704 14504
rect 12738 14532 12750 14535
rect 13342 14532 13348 14544
rect 12738 14504 13348 14532
rect 12738 14501 12750 14504
rect 12692 14495 12750 14501
rect 13342 14492 13348 14504
rect 13400 14492 13406 14544
rect 17776 14532 17804 14563
rect 19690 14560 19696 14572
rect 19748 14560 19754 14612
rect 24474 14600 24480 14612
rect 24435 14572 24480 14600
rect 24474 14560 24480 14572
rect 24532 14560 24538 14612
rect 19230 14532 19236 14544
rect 17776 14504 19236 14532
rect 19230 14492 19236 14504
rect 19288 14532 19294 14544
rect 19288 14504 19368 14532
rect 19288 14492 19294 14504
rect 11042 14464 11048 14476
rect 11003 14436 11048 14464
rect 11042 14424 11048 14436
rect 11100 14424 11106 14476
rect 16013 14467 16071 14473
rect 16013 14433 16025 14467
rect 16059 14464 16071 14467
rect 16286 14464 16292 14476
rect 16059 14436 16292 14464
rect 16059 14433 16071 14436
rect 16013 14427 16071 14433
rect 16286 14424 16292 14436
rect 16344 14424 16350 14476
rect 18126 14464 18132 14476
rect 18087 14436 18132 14464
rect 18126 14424 18132 14436
rect 18184 14424 18190 14476
rect 19340 14473 19368 14504
rect 19325 14467 19383 14473
rect 19325 14433 19337 14467
rect 19371 14433 19383 14467
rect 19325 14427 19383 14433
rect 24293 14467 24351 14473
rect 24293 14433 24305 14467
rect 24339 14464 24351 14467
rect 24382 14464 24388 14476
rect 24339 14436 24388 14464
rect 24339 14433 24351 14436
rect 24293 14427 24351 14433
rect 24382 14424 24388 14436
rect 24440 14424 24446 14476
rect 12422 14396 12428 14408
rect 12383 14368 12428 14396
rect 12422 14356 12428 14368
rect 12480 14356 12486 14408
rect 16102 14396 16108 14408
rect 16063 14368 16108 14396
rect 16102 14356 16108 14368
rect 16160 14356 16166 14408
rect 16194 14356 16200 14408
rect 16252 14396 16258 14408
rect 17669 14399 17727 14405
rect 16252 14368 16297 14396
rect 16252 14356 16258 14368
rect 17669 14365 17681 14399
rect 17715 14396 17727 14399
rect 17758 14396 17764 14408
rect 17715 14368 17764 14396
rect 17715 14365 17727 14368
rect 17669 14359 17727 14365
rect 17758 14356 17764 14368
rect 17816 14396 17822 14408
rect 18221 14399 18279 14405
rect 18221 14396 18233 14399
rect 17816 14368 18233 14396
rect 17816 14356 17822 14368
rect 18221 14365 18233 14368
rect 18267 14365 18279 14399
rect 18221 14359 18279 14365
rect 18405 14399 18463 14405
rect 18405 14365 18417 14399
rect 18451 14396 18463 14399
rect 18451 14368 18816 14396
rect 18451 14365 18463 14368
rect 18405 14359 18463 14365
rect 18788 14272 18816 14368
rect 13805 14263 13863 14269
rect 13805 14229 13817 14263
rect 13851 14260 13863 14263
rect 14170 14260 14176 14272
rect 13851 14232 14176 14260
rect 13851 14229 13863 14232
rect 13805 14223 13863 14229
rect 14170 14220 14176 14232
rect 14228 14220 14234 14272
rect 18770 14260 18776 14272
rect 18731 14232 18776 14260
rect 18770 14220 18776 14232
rect 18828 14220 18834 14272
rect 816 14170 26576 14192
rect 816 14118 5360 14170
rect 5412 14118 5424 14170
rect 5476 14118 5488 14170
rect 5540 14118 5552 14170
rect 5604 14118 14694 14170
rect 14746 14118 14758 14170
rect 14810 14118 14822 14170
rect 14874 14118 14886 14170
rect 14938 14118 24027 14170
rect 24079 14118 24091 14170
rect 24143 14118 24155 14170
rect 24207 14118 24219 14170
rect 24271 14118 26576 14170
rect 816 14096 26576 14118
rect 12514 14056 12520 14068
rect 12475 14028 12520 14056
rect 12514 14016 12520 14028
rect 12572 14016 12578 14068
rect 17577 14059 17635 14065
rect 17577 14025 17589 14059
rect 17623 14056 17635 14059
rect 18126 14056 18132 14068
rect 17623 14028 18132 14056
rect 17623 14025 17635 14028
rect 17577 14019 17635 14025
rect 18126 14016 18132 14028
rect 18184 14016 18190 14068
rect 16102 13920 16108 13932
rect 15660 13892 16108 13920
rect 11042 13852 11048 13864
rect 11003 13824 11048 13852
rect 11042 13812 11048 13824
rect 11100 13812 11106 13864
rect 14081 13855 14139 13861
rect 14081 13852 14093 13855
rect 12808 13824 14093 13852
rect 12808 13796 12836 13824
rect 14081 13821 14093 13824
rect 14127 13852 14139 13855
rect 14262 13852 14268 13864
rect 14127 13824 14268 13852
rect 14127 13821 14139 13824
rect 14081 13815 14139 13821
rect 14262 13812 14268 13824
rect 14320 13812 14326 13864
rect 14354 13812 14360 13864
rect 14412 13852 14418 13864
rect 15660 13852 15688 13892
rect 16102 13880 16108 13892
rect 16160 13920 16166 13932
rect 16565 13923 16623 13929
rect 16565 13920 16577 13923
rect 16160 13892 16577 13920
rect 16160 13880 16166 13892
rect 16565 13889 16577 13892
rect 16611 13889 16623 13923
rect 16565 13883 16623 13889
rect 17666 13880 17672 13932
rect 17724 13920 17730 13932
rect 18221 13923 18279 13929
rect 18221 13920 18233 13923
rect 17724 13892 18233 13920
rect 17724 13880 17730 13892
rect 18221 13889 18233 13892
rect 18267 13920 18279 13923
rect 18405 13923 18463 13929
rect 18405 13920 18417 13923
rect 18267 13892 18417 13920
rect 18267 13889 18279 13892
rect 18221 13883 18279 13889
rect 18405 13889 18417 13892
rect 18451 13889 18463 13923
rect 18405 13883 18463 13889
rect 16286 13852 16292 13864
rect 14412 13824 15688 13852
rect 16247 13824 16292 13852
rect 14412 13812 14418 13824
rect 16286 13812 16292 13824
rect 16344 13812 16350 13864
rect 17209 13855 17267 13861
rect 17209 13821 17221 13855
rect 17255 13852 17267 13855
rect 18420 13852 18448 13883
rect 17255 13824 18356 13852
rect 18420 13824 19000 13852
rect 17255 13821 17267 13824
rect 17209 13815 17267 13821
rect 12790 13784 12796 13796
rect 12751 13756 12796 13784
rect 12790 13744 12796 13756
rect 12848 13744 12854 13796
rect 13805 13787 13863 13793
rect 13805 13753 13817 13787
rect 13851 13784 13863 13787
rect 13894 13784 13900 13796
rect 13851 13756 13900 13784
rect 13851 13753 13863 13756
rect 13805 13747 13863 13753
rect 13894 13744 13900 13756
rect 13952 13784 13958 13796
rect 14532 13787 14590 13793
rect 14532 13784 14544 13787
rect 13952 13756 14544 13784
rect 13952 13744 13958 13756
rect 14532 13753 14544 13756
rect 14578 13784 14590 13787
rect 15734 13784 15740 13796
rect 14578 13756 15740 13784
rect 14578 13753 14590 13756
rect 14532 13747 14590 13753
rect 15734 13744 15740 13756
rect 15792 13744 15798 13796
rect 18328 13784 18356 13824
rect 18650 13787 18708 13793
rect 18650 13784 18662 13787
rect 18328 13756 18662 13784
rect 18650 13753 18662 13756
rect 18696 13784 18708 13787
rect 18770 13784 18776 13796
rect 18696 13756 18776 13784
rect 18696 13753 18708 13756
rect 18650 13747 18708 13753
rect 18770 13744 18776 13756
rect 18828 13744 18834 13796
rect 18972 13784 19000 13824
rect 19046 13784 19052 13796
rect 18972 13756 19052 13784
rect 19046 13744 19052 13756
rect 19104 13744 19110 13796
rect 15642 13716 15648 13728
rect 15603 13688 15648 13716
rect 15642 13676 15648 13688
rect 15700 13676 15706 13728
rect 19782 13716 19788 13728
rect 19743 13688 19788 13716
rect 19782 13676 19788 13688
rect 19840 13676 19846 13728
rect 24290 13716 24296 13728
rect 24251 13688 24296 13716
rect 24290 13676 24296 13688
rect 24348 13676 24354 13728
rect 816 13626 26576 13648
rect 816 13574 10027 13626
rect 10079 13574 10091 13626
rect 10143 13574 10155 13626
rect 10207 13574 10219 13626
rect 10271 13574 19360 13626
rect 19412 13574 19424 13626
rect 19476 13574 19488 13626
rect 19540 13574 19552 13626
rect 19604 13574 26576 13626
rect 816 13552 26576 13574
rect 13805 13515 13863 13521
rect 13805 13481 13817 13515
rect 13851 13512 13863 13515
rect 13894 13512 13900 13524
rect 13851 13484 13900 13512
rect 13851 13481 13863 13484
rect 13805 13475 13863 13481
rect 13894 13472 13900 13484
rect 13952 13472 13958 13524
rect 14817 13515 14875 13521
rect 14817 13481 14829 13515
rect 14863 13512 14875 13515
rect 15642 13512 15648 13524
rect 14863 13484 15648 13512
rect 14863 13481 14875 13484
rect 14817 13475 14875 13481
rect 15642 13472 15648 13484
rect 15700 13472 15706 13524
rect 16105 13515 16163 13521
rect 16105 13481 16117 13515
rect 16151 13512 16163 13515
rect 16194 13512 16200 13524
rect 16151 13484 16200 13512
rect 16151 13481 16163 13484
rect 16105 13475 16163 13481
rect 16194 13472 16200 13484
rect 16252 13472 16258 13524
rect 18770 13512 18776 13524
rect 18731 13484 18776 13512
rect 18770 13472 18776 13484
rect 18828 13472 18834 13524
rect 19230 13472 19236 13524
rect 19288 13512 19294 13524
rect 19325 13515 19383 13521
rect 19325 13512 19337 13515
rect 19288 13484 19337 13512
rect 19288 13472 19294 13484
rect 19325 13481 19337 13484
rect 19371 13481 19383 13515
rect 19325 13475 19383 13481
rect 23373 13515 23431 13521
rect 23373 13481 23385 13515
rect 23419 13512 23431 13515
rect 24290 13512 24296 13524
rect 23419 13484 24296 13512
rect 23419 13481 23431 13484
rect 23373 13475 23431 13481
rect 24290 13472 24296 13484
rect 24348 13472 24354 13524
rect 12790 13444 12796 13456
rect 12440 13416 12796 13444
rect 12440 13385 12468 13416
rect 12790 13404 12796 13416
rect 12848 13404 12854 13456
rect 12425 13379 12483 13385
rect 12425 13345 12437 13379
rect 12471 13345 12483 13379
rect 12425 13339 12483 13345
rect 12514 13336 12520 13388
rect 12572 13376 12578 13388
rect 12692 13379 12750 13385
rect 12692 13376 12704 13379
rect 12572 13348 12704 13376
rect 12572 13336 12578 13348
rect 12692 13345 12704 13348
rect 12738 13376 12750 13379
rect 14170 13376 14176 13388
rect 12738 13348 14176 13376
rect 12738 13345 12750 13348
rect 12692 13339 12750 13345
rect 14170 13336 14176 13348
rect 14228 13336 14234 13388
rect 15366 13376 15372 13388
rect 15327 13348 15372 13376
rect 15366 13336 15372 13348
rect 15424 13336 15430 13388
rect 17660 13379 17718 13385
rect 17660 13345 17672 13379
rect 17706 13376 17718 13379
rect 18034 13376 18040 13388
rect 17706 13348 18040 13376
rect 17706 13345 17718 13348
rect 17660 13339 17718 13345
rect 18034 13336 18040 13348
rect 18092 13336 18098 13388
rect 23189 13379 23247 13385
rect 23189 13345 23201 13379
rect 23235 13376 23247 13379
rect 23554 13376 23560 13388
rect 23235 13348 23560 13376
rect 23235 13345 23247 13348
rect 23189 13339 23247 13345
rect 23554 13336 23560 13348
rect 23612 13336 23618 13388
rect 13618 13268 13624 13320
rect 13676 13308 13682 13320
rect 14449 13311 14507 13317
rect 14449 13308 14461 13311
rect 13676 13280 14461 13308
rect 13676 13268 13682 13280
rect 14449 13277 14461 13280
rect 14495 13308 14507 13311
rect 15461 13311 15519 13317
rect 15461 13308 15473 13311
rect 14495 13280 15473 13308
rect 14495 13277 14507 13280
rect 14449 13271 14507 13277
rect 15461 13277 15473 13280
rect 15507 13277 15519 13311
rect 15461 13271 15519 13277
rect 15645 13311 15703 13317
rect 15645 13277 15657 13311
rect 15691 13308 15703 13311
rect 15734 13308 15740 13320
rect 15691 13280 15740 13308
rect 15691 13277 15703 13280
rect 15645 13271 15703 13277
rect 15734 13268 15740 13280
rect 15792 13268 15798 13320
rect 17390 13308 17396 13320
rect 17351 13280 17396 13308
rect 17390 13268 17396 13280
rect 17448 13268 17454 13320
rect 20610 13308 20616 13320
rect 20571 13280 20616 13308
rect 20610 13268 20616 13280
rect 20668 13268 20674 13320
rect 14538 13200 14544 13252
rect 14596 13240 14602 13252
rect 15001 13243 15059 13249
rect 15001 13240 15013 13243
rect 14596 13212 15013 13240
rect 14596 13200 14602 13212
rect 15001 13209 15013 13212
rect 15047 13209 15059 13243
rect 15001 13203 15059 13209
rect 816 13082 26576 13104
rect 816 13030 5360 13082
rect 5412 13030 5424 13082
rect 5476 13030 5488 13082
rect 5540 13030 5552 13082
rect 5604 13030 14694 13082
rect 14746 13030 14758 13082
rect 14810 13030 14822 13082
rect 14874 13030 14886 13082
rect 14938 13030 24027 13082
rect 24079 13030 24091 13082
rect 24143 13030 24155 13082
rect 24207 13030 24219 13082
rect 24271 13030 26576 13082
rect 816 13008 26576 13030
rect 12790 12928 12796 12980
rect 12848 12968 12854 12980
rect 13069 12971 13127 12977
rect 13069 12968 13081 12971
rect 12848 12940 13081 12968
rect 12848 12928 12854 12940
rect 13069 12937 13081 12940
rect 13115 12937 13127 12971
rect 13618 12968 13624 12980
rect 13579 12940 13624 12968
rect 13069 12931 13127 12937
rect 13618 12928 13624 12940
rect 13676 12928 13682 12980
rect 14446 12928 14452 12980
rect 14504 12968 14510 12980
rect 14725 12971 14783 12977
rect 14725 12968 14737 12971
rect 14504 12940 14737 12968
rect 14504 12928 14510 12940
rect 14725 12937 14737 12940
rect 14771 12968 14783 12971
rect 15366 12968 15372 12980
rect 14771 12940 15372 12968
rect 14771 12937 14783 12940
rect 14725 12931 14783 12937
rect 15366 12928 15372 12940
rect 15424 12928 15430 12980
rect 16194 12928 16200 12980
rect 16252 12968 16258 12980
rect 16562 12968 16568 12980
rect 16252 12940 16568 12968
rect 16252 12928 16258 12940
rect 16562 12928 16568 12940
rect 16620 12928 16626 12980
rect 17666 12928 17672 12980
rect 17724 12968 17730 12980
rect 18034 12968 18040 12980
rect 17724 12940 18040 12968
rect 17724 12928 17730 12940
rect 18034 12928 18040 12940
rect 18092 12968 18098 12980
rect 18310 12968 18316 12980
rect 18092 12940 18316 12968
rect 18092 12928 18098 12940
rect 18310 12928 18316 12940
rect 18368 12928 18374 12980
rect 19046 12968 19052 12980
rect 19007 12940 19052 12968
rect 19046 12928 19052 12940
rect 19104 12968 19110 12980
rect 19230 12968 19236 12980
rect 19104 12940 19236 12968
rect 19104 12928 19110 12940
rect 19230 12928 19236 12940
rect 19288 12928 19294 12980
rect 14262 12860 14268 12912
rect 14320 12900 14326 12912
rect 15001 12903 15059 12909
rect 15001 12900 15013 12903
rect 14320 12872 15013 12900
rect 14320 12860 14326 12872
rect 15001 12869 15013 12872
rect 15047 12900 15059 12903
rect 15047 12872 15228 12900
rect 15047 12869 15059 12872
rect 15001 12863 15059 12869
rect 14170 12832 14176 12844
rect 14131 12804 14176 12832
rect 14170 12792 14176 12804
rect 14228 12792 14234 12844
rect 15200 12841 15228 12872
rect 15185 12835 15243 12841
rect 15185 12801 15197 12835
rect 15231 12801 15243 12835
rect 15185 12795 15243 12801
rect 17853 12835 17911 12841
rect 17853 12801 17865 12835
rect 17899 12832 17911 12835
rect 18126 12832 18132 12844
rect 17899 12804 18132 12832
rect 17899 12801 17911 12804
rect 17853 12795 17911 12801
rect 12149 12767 12207 12773
rect 12149 12733 12161 12767
rect 12195 12764 12207 12767
rect 12698 12764 12704 12776
rect 12195 12736 12704 12764
rect 12195 12733 12207 12736
rect 12149 12727 12207 12733
rect 12698 12724 12704 12736
rect 12756 12724 12762 12776
rect 15200 12764 15228 12795
rect 18126 12792 18132 12804
rect 18184 12792 18190 12844
rect 19230 12832 19236 12844
rect 19191 12804 19236 12832
rect 19230 12792 19236 12804
rect 19288 12792 19294 12844
rect 16378 12764 16384 12776
rect 15200 12736 16384 12764
rect 16378 12724 16384 12736
rect 16436 12764 16442 12776
rect 17390 12764 17396 12776
rect 16436 12736 17396 12764
rect 16436 12724 16442 12736
rect 17390 12724 17396 12736
rect 17448 12724 17454 12776
rect 19500 12767 19558 12773
rect 19500 12764 19512 12767
rect 19340 12736 19512 12764
rect 13526 12696 13532 12708
rect 13439 12668 13532 12696
rect 13526 12656 13532 12668
rect 13584 12696 13590 12708
rect 13989 12699 14047 12705
rect 13989 12696 14001 12699
rect 13584 12668 14001 12696
rect 13584 12656 13590 12668
rect 13989 12665 14001 12668
rect 14035 12665 14047 12699
rect 13989 12659 14047 12665
rect 15452 12699 15510 12705
rect 15452 12665 15464 12699
rect 15498 12696 15510 12699
rect 15642 12696 15648 12708
rect 15498 12668 15648 12696
rect 15498 12665 15510 12668
rect 15452 12659 15510 12665
rect 15642 12656 15648 12668
rect 15700 12656 15706 12708
rect 18773 12699 18831 12705
rect 18773 12665 18785 12699
rect 18819 12696 18831 12699
rect 18862 12696 18868 12708
rect 18819 12668 18868 12696
rect 18819 12665 18831 12668
rect 18773 12659 18831 12665
rect 18862 12656 18868 12668
rect 18920 12696 18926 12708
rect 19340 12696 19368 12736
rect 19500 12733 19512 12736
rect 19546 12764 19558 12767
rect 19782 12764 19788 12776
rect 19546 12736 19788 12764
rect 19546 12733 19558 12736
rect 19500 12727 19558 12733
rect 19782 12724 19788 12736
rect 19840 12724 19846 12776
rect 23554 12764 23560 12776
rect 23515 12736 23560 12764
rect 23554 12724 23560 12736
rect 23612 12724 23618 12776
rect 18920 12668 19368 12696
rect 18920 12656 18926 12668
rect 12330 12628 12336 12640
rect 12291 12600 12336 12628
rect 12330 12588 12336 12600
rect 12388 12588 12394 12640
rect 14078 12628 14084 12640
rect 14039 12600 14084 12628
rect 14078 12588 14084 12600
rect 14136 12588 14142 12640
rect 20613 12631 20671 12637
rect 20613 12597 20625 12631
rect 20659 12628 20671 12631
rect 21162 12628 21168 12640
rect 20659 12600 21168 12628
rect 20659 12597 20671 12600
rect 20613 12591 20671 12597
rect 21162 12588 21168 12600
rect 21220 12588 21226 12640
rect 816 12538 26576 12560
rect 816 12486 10027 12538
rect 10079 12486 10091 12538
rect 10143 12486 10155 12538
rect 10207 12486 10219 12538
rect 10271 12486 19360 12538
rect 19412 12486 19424 12538
rect 19476 12486 19488 12538
rect 19540 12486 19552 12538
rect 19604 12486 26576 12538
rect 816 12464 26576 12486
rect 12514 12424 12520 12436
rect 12475 12396 12520 12424
rect 12514 12384 12520 12396
rect 12572 12384 12578 12436
rect 14081 12427 14139 12433
rect 14081 12393 14093 12427
rect 14127 12393 14139 12427
rect 14081 12387 14139 12393
rect 13897 12291 13955 12297
rect 13897 12257 13909 12291
rect 13943 12257 13955 12291
rect 14096 12288 14124 12387
rect 14170 12384 14176 12436
rect 14228 12424 14234 12436
rect 14357 12427 14415 12433
rect 14357 12424 14369 12427
rect 14228 12396 14369 12424
rect 14228 12384 14234 12396
rect 14357 12393 14369 12396
rect 14403 12393 14415 12427
rect 15366 12424 15372 12436
rect 15327 12396 15372 12424
rect 14357 12387 14415 12393
rect 15366 12384 15372 12396
rect 15424 12384 15430 12436
rect 15734 12424 15740 12436
rect 15695 12396 15740 12424
rect 15734 12384 15740 12396
rect 15792 12384 15798 12436
rect 17666 12424 17672 12436
rect 17627 12396 17672 12424
rect 17666 12384 17672 12396
rect 17724 12384 17730 12436
rect 18865 12427 18923 12433
rect 18865 12393 18877 12427
rect 18911 12393 18923 12427
rect 18865 12387 18923 12393
rect 14817 12359 14875 12365
rect 14817 12325 14829 12359
rect 14863 12356 14875 12359
rect 15642 12356 15648 12368
rect 14863 12328 15648 12356
rect 14863 12325 14875 12328
rect 14817 12319 14875 12325
rect 15642 12316 15648 12328
rect 15700 12316 15706 12368
rect 18880 12356 18908 12387
rect 19138 12384 19144 12436
rect 19196 12424 19202 12436
rect 19325 12427 19383 12433
rect 19325 12424 19337 12427
rect 19196 12396 19337 12424
rect 19196 12384 19202 12396
rect 19325 12393 19337 12396
rect 19371 12393 19383 12427
rect 19325 12387 19383 12393
rect 20610 12384 20616 12436
rect 20668 12424 20674 12436
rect 20981 12427 21039 12433
rect 20981 12424 20993 12427
rect 20668 12396 20993 12424
rect 20668 12384 20674 12396
rect 20981 12393 20993 12396
rect 21027 12424 21039 12427
rect 21346 12424 21352 12436
rect 21027 12396 21352 12424
rect 21027 12393 21039 12396
rect 20981 12387 21039 12393
rect 21346 12384 21352 12396
rect 21404 12384 21410 12436
rect 21073 12359 21131 12365
rect 21073 12356 21085 12359
rect 18880 12328 21085 12356
rect 21073 12325 21085 12328
rect 21119 12356 21131 12359
rect 22082 12356 22088 12368
rect 21119 12328 22088 12356
rect 21119 12325 21131 12328
rect 21073 12319 21131 12325
rect 22082 12316 22088 12328
rect 22140 12316 22146 12368
rect 15185 12291 15243 12297
rect 15185 12288 15197 12291
rect 14096 12260 15197 12288
rect 13897 12251 13955 12257
rect 15185 12257 15197 12260
rect 15231 12288 15243 12291
rect 15734 12288 15740 12300
rect 15231 12260 15740 12288
rect 15231 12257 15243 12260
rect 15185 12251 15243 12257
rect 13912 12220 13940 12251
rect 15734 12248 15740 12260
rect 15792 12248 15798 12300
rect 16289 12291 16347 12297
rect 16289 12257 16301 12291
rect 16335 12288 16347 12291
rect 16378 12288 16384 12300
rect 16335 12260 16384 12288
rect 16335 12257 16347 12260
rect 16289 12251 16347 12257
rect 16378 12248 16384 12260
rect 16436 12248 16442 12300
rect 16562 12297 16568 12300
rect 16556 12288 16568 12297
rect 16475 12260 16568 12288
rect 16556 12251 16568 12260
rect 16620 12288 16626 12300
rect 17114 12288 17120 12300
rect 16620 12260 17120 12288
rect 16562 12248 16568 12251
rect 16620 12248 16626 12260
rect 17114 12248 17120 12260
rect 17172 12248 17178 12300
rect 18770 12248 18776 12300
rect 18828 12288 18834 12300
rect 19233 12291 19291 12297
rect 19233 12288 19245 12291
rect 18828 12260 19245 12288
rect 18828 12248 18834 12260
rect 19233 12257 19245 12260
rect 19279 12257 19291 12291
rect 19233 12251 19291 12257
rect 14538 12220 14544 12232
rect 13912 12192 14544 12220
rect 14538 12180 14544 12192
rect 14596 12180 14602 12232
rect 19509 12223 19567 12229
rect 19509 12189 19521 12223
rect 19555 12220 19567 12223
rect 19782 12220 19788 12232
rect 19555 12192 19788 12220
rect 19555 12189 19567 12192
rect 19509 12183 19567 12189
rect 19782 12180 19788 12192
rect 19840 12180 19846 12232
rect 21162 12180 21168 12232
rect 21220 12220 21226 12232
rect 21220 12192 21265 12220
rect 21220 12180 21226 12192
rect 20613 12155 20671 12161
rect 20613 12121 20625 12155
rect 20659 12152 20671 12155
rect 21714 12152 21720 12164
rect 20659 12124 21720 12152
rect 20659 12121 20671 12124
rect 20613 12115 20671 12121
rect 21714 12112 21720 12124
rect 21772 12112 21778 12164
rect 13713 12087 13771 12093
rect 13713 12053 13725 12087
rect 13759 12084 13771 12087
rect 14078 12084 14084 12096
rect 13759 12056 14084 12084
rect 13759 12053 13771 12056
rect 13713 12047 13771 12053
rect 14078 12044 14084 12056
rect 14136 12084 14142 12096
rect 15182 12084 15188 12096
rect 14136 12056 15188 12084
rect 14136 12044 14142 12056
rect 15182 12044 15188 12056
rect 15240 12044 15246 12096
rect 816 11994 26576 12016
rect 816 11942 5360 11994
rect 5412 11942 5424 11994
rect 5476 11942 5488 11994
rect 5540 11942 5552 11994
rect 5604 11942 14694 11994
rect 14746 11942 14758 11994
rect 14810 11942 14822 11994
rect 14874 11942 14886 11994
rect 14938 11942 24027 11994
rect 24079 11942 24091 11994
rect 24143 11942 24155 11994
rect 24207 11942 24219 11994
rect 24271 11942 26576 11994
rect 816 11920 26576 11942
rect 14265 11883 14323 11889
rect 14265 11849 14277 11883
rect 14311 11880 14323 11883
rect 14538 11880 14544 11892
rect 14311 11852 14544 11880
rect 14311 11849 14323 11852
rect 14265 11843 14323 11849
rect 14538 11840 14544 11852
rect 14596 11840 14602 11892
rect 15734 11880 15740 11892
rect 15695 11852 15740 11880
rect 15734 11840 15740 11852
rect 15792 11840 15798 11892
rect 17114 11880 17120 11892
rect 17075 11852 17120 11880
rect 17114 11840 17120 11852
rect 17172 11840 17178 11892
rect 17758 11880 17764 11892
rect 17719 11852 17764 11880
rect 17758 11840 17764 11852
rect 17816 11840 17822 11892
rect 21346 11880 21352 11892
rect 21307 11852 21352 11880
rect 21346 11840 21352 11852
rect 21404 11840 21410 11892
rect 22082 11880 22088 11892
rect 22043 11852 22088 11880
rect 22082 11840 22088 11852
rect 22140 11840 22146 11892
rect 14354 11772 14360 11824
rect 14412 11812 14418 11824
rect 14725 11815 14783 11821
rect 14725 11812 14737 11815
rect 14412 11784 14737 11812
rect 14412 11772 14418 11784
rect 14725 11781 14737 11784
rect 14771 11781 14783 11815
rect 14725 11775 14783 11781
rect 16841 11815 16899 11821
rect 16841 11781 16853 11815
rect 16887 11812 16899 11815
rect 17390 11812 17396 11824
rect 16887 11784 17396 11812
rect 16887 11781 16899 11784
rect 16841 11775 16899 11781
rect 17390 11772 17396 11784
rect 17448 11772 17454 11824
rect 21162 11772 21168 11824
rect 21220 11812 21226 11824
rect 21717 11815 21775 11821
rect 21717 11812 21729 11815
rect 21220 11784 21729 11812
rect 21220 11772 21226 11784
rect 21717 11781 21729 11784
rect 21763 11781 21775 11815
rect 21717 11775 21775 11781
rect 13713 11747 13771 11753
rect 13713 11713 13725 11747
rect 13759 11744 13771 11747
rect 14446 11744 14452 11756
rect 13759 11716 14452 11744
rect 13759 11713 13771 11716
rect 13713 11707 13771 11713
rect 14446 11704 14452 11716
rect 14504 11704 14510 11756
rect 15369 11747 15427 11753
rect 15369 11713 15381 11747
rect 15415 11744 15427 11747
rect 15642 11744 15648 11756
rect 15415 11716 15648 11744
rect 15415 11713 15427 11716
rect 15369 11707 15427 11713
rect 15642 11704 15648 11716
rect 15700 11704 15706 11756
rect 16286 11704 16292 11756
rect 16344 11744 16350 11756
rect 18310 11744 18316 11756
rect 16344 11716 16389 11744
rect 18271 11716 18316 11744
rect 16344 11704 16350 11716
rect 18310 11704 18316 11716
rect 18368 11704 18374 11756
rect 18221 11679 18279 11685
rect 18221 11645 18233 11679
rect 18267 11676 18279 11679
rect 19046 11676 19052 11688
rect 18267 11648 19052 11676
rect 18267 11645 18279 11648
rect 18221 11639 18279 11645
rect 19046 11636 19052 11648
rect 19104 11636 19110 11688
rect 19230 11636 19236 11688
rect 19288 11676 19294 11688
rect 19417 11679 19475 11685
rect 19417 11676 19429 11679
rect 19288 11648 19429 11676
rect 19288 11636 19294 11648
rect 19417 11645 19429 11648
rect 19463 11645 19475 11679
rect 19417 11639 19475 11645
rect 24293 11679 24351 11685
rect 24293 11645 24305 11679
rect 24339 11676 24351 11679
rect 24474 11676 24480 11688
rect 24339 11648 24480 11676
rect 24339 11645 24351 11648
rect 24293 11639 24351 11645
rect 15093 11611 15151 11617
rect 15093 11608 15105 11611
rect 14556 11580 15105 11608
rect 14556 11552 14584 11580
rect 15093 11577 15105 11580
rect 15139 11577 15151 11611
rect 18129 11611 18187 11617
rect 18129 11608 18141 11611
rect 15093 11571 15151 11577
rect 17500 11580 18141 11608
rect 17500 11552 17528 11580
rect 18129 11577 18141 11580
rect 18175 11577 18187 11611
rect 18129 11571 18187 11577
rect 14538 11540 14544 11552
rect 14499 11512 14544 11540
rect 14538 11500 14544 11512
rect 14596 11500 14602 11552
rect 15182 11540 15188 11552
rect 15143 11512 15188 11540
rect 15182 11500 15188 11512
rect 15240 11500 15246 11552
rect 17482 11540 17488 11552
rect 17443 11512 17488 11540
rect 17482 11500 17488 11512
rect 17540 11500 17546 11552
rect 18770 11500 18776 11552
rect 18828 11540 18834 11552
rect 18865 11543 18923 11549
rect 18865 11540 18877 11543
rect 18828 11512 18877 11540
rect 18828 11500 18834 11512
rect 18865 11509 18877 11512
rect 18911 11509 18923 11543
rect 18865 11503 18923 11509
rect 19325 11543 19383 11549
rect 19325 11509 19337 11543
rect 19371 11540 19383 11543
rect 19432 11540 19460 11639
rect 24474 11636 24480 11648
rect 24532 11676 24538 11688
rect 24845 11679 24903 11685
rect 24845 11676 24857 11679
rect 24532 11648 24857 11676
rect 24532 11636 24538 11648
rect 24845 11645 24857 11648
rect 24891 11645 24903 11679
rect 24845 11639 24903 11645
rect 19684 11611 19742 11617
rect 19684 11577 19696 11611
rect 19730 11608 19742 11611
rect 19782 11608 19788 11620
rect 19730 11580 19788 11608
rect 19730 11577 19742 11580
rect 19684 11571 19742 11577
rect 19782 11568 19788 11580
rect 19840 11568 19846 11620
rect 20242 11540 20248 11552
rect 19371 11512 20248 11540
rect 19371 11509 19383 11512
rect 19325 11503 19383 11509
rect 20242 11500 20248 11512
rect 20300 11500 20306 11552
rect 20426 11500 20432 11552
rect 20484 11540 20490 11552
rect 20797 11543 20855 11549
rect 20797 11540 20809 11543
rect 20484 11512 20809 11540
rect 20484 11500 20490 11512
rect 20797 11509 20809 11512
rect 20843 11509 20855 11543
rect 24474 11540 24480 11552
rect 24435 11512 24480 11540
rect 20797 11503 20855 11509
rect 24474 11500 24480 11512
rect 24532 11500 24538 11552
rect 816 11450 26576 11472
rect 816 11398 10027 11450
rect 10079 11398 10091 11450
rect 10143 11398 10155 11450
rect 10207 11398 10219 11450
rect 10271 11398 19360 11450
rect 19412 11398 19424 11450
rect 19476 11398 19488 11450
rect 19540 11398 19552 11450
rect 19604 11398 26576 11450
rect 816 11376 26576 11398
rect 18221 11339 18279 11345
rect 18221 11305 18233 11339
rect 18267 11336 18279 11339
rect 18310 11336 18316 11348
rect 18267 11308 18316 11336
rect 18267 11305 18279 11308
rect 18221 11299 18279 11305
rect 18310 11296 18316 11308
rect 18368 11296 18374 11348
rect 18862 11336 18868 11348
rect 18823 11308 18868 11336
rect 18862 11296 18868 11308
rect 18920 11296 18926 11348
rect 19046 11296 19052 11348
rect 19104 11336 19110 11348
rect 19417 11339 19475 11345
rect 19417 11336 19429 11339
rect 19104 11308 19429 11336
rect 19104 11296 19110 11308
rect 19417 11305 19429 11308
rect 19463 11305 19475 11339
rect 19782 11336 19788 11348
rect 19743 11308 19788 11336
rect 19417 11299 19475 11305
rect 19782 11296 19788 11308
rect 19840 11296 19846 11348
rect 14817 11271 14875 11277
rect 14817 11237 14829 11271
rect 14863 11268 14875 11271
rect 15182 11268 15188 11280
rect 14863 11240 15188 11268
rect 14863 11237 14875 11240
rect 14817 11231 14875 11237
rect 15182 11228 15188 11240
rect 15240 11268 15246 11280
rect 17853 11271 17911 11277
rect 17853 11268 17865 11271
rect 15240 11240 17865 11268
rect 15240 11228 15246 11240
rect 17853 11237 17865 11240
rect 17899 11268 17911 11271
rect 19064 11268 19092 11296
rect 17899 11240 19092 11268
rect 20429 11271 20487 11277
rect 17899 11237 17911 11240
rect 17853 11231 17911 11237
rect 20429 11237 20441 11271
rect 20475 11268 20487 11271
rect 20880 11271 20938 11277
rect 20880 11268 20892 11271
rect 20475 11240 20892 11268
rect 20475 11237 20487 11240
rect 20429 11231 20487 11237
rect 20880 11237 20892 11240
rect 20926 11268 20938 11271
rect 21162 11268 21168 11280
rect 20926 11240 21168 11268
rect 20926 11237 20938 11240
rect 20880 11231 20938 11237
rect 21162 11228 21168 11240
rect 21220 11228 21226 11280
rect 18957 11135 19015 11141
rect 18957 11101 18969 11135
rect 19003 11101 19015 11135
rect 18957 11095 19015 11101
rect 18972 10996 19000 11095
rect 20242 11092 20248 11144
rect 20300 11132 20306 11144
rect 20613 11135 20671 11141
rect 20613 11132 20625 11135
rect 20300 11104 20625 11132
rect 20300 11092 20306 11104
rect 20613 11101 20625 11104
rect 20659 11101 20671 11135
rect 20613 11095 20671 11101
rect 19782 11024 19788 11076
rect 19840 11064 19846 11076
rect 19840 11036 20380 11064
rect 19840 11024 19846 11036
rect 19230 10996 19236 11008
rect 18972 10968 19236 10996
rect 19230 10956 19236 10968
rect 19288 10956 19294 11008
rect 20352 10996 20380 11036
rect 21993 10999 22051 11005
rect 21993 10996 22005 10999
rect 20352 10968 22005 10996
rect 21993 10965 22005 10968
rect 22039 10996 22051 10999
rect 22358 10996 22364 11008
rect 22039 10968 22364 10996
rect 22039 10965 22051 10968
rect 21993 10959 22051 10965
rect 22358 10956 22364 10968
rect 22416 10956 22422 11008
rect 816 10906 26576 10928
rect 816 10854 5360 10906
rect 5412 10854 5424 10906
rect 5476 10854 5488 10906
rect 5540 10854 5552 10906
rect 5604 10854 14694 10906
rect 14746 10854 14758 10906
rect 14810 10854 14822 10906
rect 14874 10854 14886 10906
rect 14938 10854 24027 10906
rect 24079 10854 24091 10906
rect 24143 10854 24155 10906
rect 24207 10854 24219 10906
rect 24271 10854 26576 10906
rect 816 10832 26576 10854
rect 21073 10659 21131 10665
rect 21073 10625 21085 10659
rect 21119 10656 21131 10659
rect 22177 10659 22235 10665
rect 21119 10628 22036 10656
rect 21119 10625 21131 10628
rect 21073 10619 21131 10625
rect 14633 10591 14691 10597
rect 14633 10557 14645 10591
rect 14679 10557 14691 10591
rect 14633 10551 14691 10557
rect 14648 10520 14676 10551
rect 18678 10548 18684 10600
rect 18736 10588 18742 10600
rect 19049 10591 19107 10597
rect 19049 10588 19061 10591
rect 18736 10560 19061 10588
rect 18736 10548 18742 10560
rect 19049 10557 19061 10560
rect 19095 10557 19107 10591
rect 19316 10591 19374 10597
rect 19316 10588 19328 10591
rect 19049 10551 19107 10557
rect 19248 10560 19328 10588
rect 15274 10520 15280 10532
rect 14648 10492 15280 10520
rect 15274 10480 15280 10492
rect 15332 10480 15338 10532
rect 18034 10480 18040 10532
rect 18092 10520 18098 10532
rect 18589 10523 18647 10529
rect 18589 10520 18601 10523
rect 18092 10492 18601 10520
rect 18092 10480 18098 10492
rect 18589 10489 18601 10492
rect 18635 10520 18647 10523
rect 19248 10520 19276 10560
rect 19316 10557 19328 10560
rect 19362 10588 19374 10591
rect 19690 10588 19696 10600
rect 19362 10560 19696 10588
rect 19362 10557 19374 10560
rect 19316 10551 19374 10557
rect 19690 10548 19696 10560
rect 19748 10588 19754 10600
rect 20334 10588 20340 10600
rect 19748 10560 20340 10588
rect 19748 10548 19754 10560
rect 20334 10548 20340 10560
rect 20392 10548 20398 10600
rect 20978 10548 20984 10600
rect 21036 10588 21042 10600
rect 22008 10597 22036 10628
rect 22177 10625 22189 10659
rect 22223 10656 22235 10659
rect 22358 10656 22364 10668
rect 22223 10628 22364 10656
rect 22223 10625 22235 10628
rect 22177 10619 22235 10625
rect 22358 10616 22364 10628
rect 22416 10616 22422 10668
rect 21349 10591 21407 10597
rect 21349 10588 21361 10591
rect 21036 10560 21361 10588
rect 21036 10548 21042 10560
rect 21349 10557 21361 10560
rect 21395 10588 21407 10591
rect 21901 10591 21959 10597
rect 21901 10588 21913 10591
rect 21395 10560 21913 10588
rect 21395 10557 21407 10560
rect 21349 10551 21407 10557
rect 21901 10557 21913 10560
rect 21947 10557 21959 10591
rect 21901 10551 21959 10557
rect 21993 10591 22051 10597
rect 21993 10557 22005 10591
rect 22039 10588 22051 10591
rect 23094 10588 23100 10600
rect 22039 10560 23100 10588
rect 22039 10557 22051 10560
rect 21993 10551 22051 10557
rect 23094 10548 23100 10560
rect 23152 10548 23158 10600
rect 18635 10492 19276 10520
rect 18635 10489 18647 10492
rect 18589 10483 18647 10489
rect 14538 10412 14544 10464
rect 14596 10452 14602 10464
rect 14817 10455 14875 10461
rect 14817 10452 14829 10455
rect 14596 10424 14829 10452
rect 14596 10412 14602 10424
rect 14817 10421 14829 10424
rect 14863 10421 14875 10455
rect 14817 10415 14875 10421
rect 18678 10412 18684 10464
rect 18736 10452 18742 10464
rect 18865 10455 18923 10461
rect 18865 10452 18877 10455
rect 18736 10424 18877 10452
rect 18736 10412 18742 10424
rect 18865 10421 18877 10424
rect 18911 10421 18923 10455
rect 20426 10452 20432 10464
rect 20387 10424 20432 10452
rect 18865 10415 18923 10421
rect 20426 10412 20432 10424
rect 20484 10412 20490 10464
rect 21530 10452 21536 10464
rect 21491 10424 21536 10452
rect 21530 10412 21536 10424
rect 21588 10412 21594 10464
rect 816 10362 26576 10384
rect 816 10310 10027 10362
rect 10079 10310 10091 10362
rect 10143 10310 10155 10362
rect 10207 10310 10219 10362
rect 10271 10310 19360 10362
rect 19412 10310 19424 10362
rect 19476 10310 19488 10362
rect 19540 10310 19552 10362
rect 19604 10310 26576 10362
rect 816 10288 26576 10310
rect 21070 10248 21076 10260
rect 21031 10220 21076 10248
rect 21070 10208 21076 10220
rect 21128 10208 21134 10260
rect 21717 10251 21775 10257
rect 21717 10217 21729 10251
rect 21763 10248 21775 10251
rect 22358 10248 22364 10260
rect 21763 10220 22364 10248
rect 21763 10217 21775 10220
rect 21717 10211 21775 10217
rect 22358 10208 22364 10220
rect 22416 10208 22422 10260
rect 18405 10183 18463 10189
rect 18405 10149 18417 10183
rect 18451 10180 18463 10183
rect 19325 10183 19383 10189
rect 19325 10180 19337 10183
rect 18451 10152 19337 10180
rect 18451 10149 18463 10152
rect 18405 10143 18463 10149
rect 19325 10149 19337 10152
rect 19371 10180 19383 10183
rect 21530 10180 21536 10192
rect 19371 10152 21536 10180
rect 19371 10149 19383 10152
rect 19325 10143 19383 10149
rect 21530 10140 21536 10152
rect 21588 10140 21594 10192
rect 19230 10112 19236 10124
rect 19191 10084 19236 10112
rect 19230 10072 19236 10084
rect 19288 10072 19294 10124
rect 20978 10112 20984 10124
rect 20939 10084 20984 10112
rect 20978 10072 20984 10084
rect 21036 10072 21042 10124
rect 19509 10047 19567 10053
rect 19509 10013 19521 10047
rect 19555 10044 19567 10047
rect 19690 10044 19696 10056
rect 19555 10016 19696 10044
rect 19555 10013 19567 10016
rect 19509 10007 19567 10013
rect 19690 10004 19696 10016
rect 19748 10004 19754 10056
rect 20426 10004 20432 10056
rect 20484 10044 20490 10056
rect 21165 10047 21223 10053
rect 21165 10044 21177 10047
rect 20484 10016 21177 10044
rect 20484 10004 20490 10016
rect 21165 10013 21177 10016
rect 21211 10013 21223 10047
rect 21165 10007 21223 10013
rect 18773 9979 18831 9985
rect 18773 9945 18785 9979
rect 18819 9976 18831 9979
rect 19046 9976 19052 9988
rect 18819 9948 19052 9976
rect 18819 9945 18831 9948
rect 18773 9939 18831 9945
rect 19046 9936 19052 9948
rect 19104 9936 19110 9988
rect 18862 9908 18868 9920
rect 18823 9880 18868 9908
rect 18862 9868 18868 9880
rect 18920 9868 18926 9920
rect 20334 9908 20340 9920
rect 20295 9880 20340 9908
rect 20334 9868 20340 9880
rect 20392 9868 20398 9920
rect 20610 9908 20616 9920
rect 20571 9880 20616 9908
rect 20610 9868 20616 9880
rect 20668 9868 20674 9920
rect 816 9818 26576 9840
rect 816 9766 5360 9818
rect 5412 9766 5424 9818
rect 5476 9766 5488 9818
rect 5540 9766 5552 9818
rect 5604 9766 14694 9818
rect 14746 9766 14758 9818
rect 14810 9766 14822 9818
rect 14874 9766 14886 9818
rect 14938 9766 24027 9818
rect 24079 9766 24091 9818
rect 24143 9766 24155 9818
rect 24207 9766 24219 9818
rect 24271 9766 26576 9818
rect 816 9744 26576 9766
rect 18034 9704 18040 9716
rect 17995 9676 18040 9704
rect 18034 9664 18040 9676
rect 18092 9664 18098 9716
rect 19230 9704 19236 9716
rect 18880 9676 19236 9704
rect 18405 9639 18463 9645
rect 18405 9605 18417 9639
rect 18451 9636 18463 9639
rect 18880 9636 18908 9676
rect 19230 9664 19236 9676
rect 19288 9664 19294 9716
rect 21070 9664 21076 9716
rect 21128 9704 21134 9716
rect 21165 9707 21223 9713
rect 21165 9704 21177 9707
rect 21128 9676 21177 9704
rect 21128 9664 21134 9676
rect 21165 9673 21177 9676
rect 21211 9673 21223 9707
rect 21165 9667 21223 9673
rect 21990 9664 21996 9716
rect 22048 9704 22054 9716
rect 22266 9704 22272 9716
rect 22048 9676 22272 9704
rect 22048 9664 22054 9676
rect 22266 9664 22272 9676
rect 22324 9664 22330 9716
rect 18451 9608 18908 9636
rect 18451 9605 18463 9608
rect 18405 9599 18463 9605
rect 14906 9568 14912 9580
rect 14372 9540 14912 9568
rect 14372 9509 14400 9540
rect 14906 9528 14912 9540
rect 14964 9528 14970 9580
rect 14357 9503 14415 9509
rect 14357 9469 14369 9503
rect 14403 9469 14415 9503
rect 14357 9463 14415 9469
rect 18678 9460 18684 9512
rect 18736 9500 18742 9512
rect 18865 9503 18923 9509
rect 18865 9500 18877 9503
rect 18736 9472 18877 9500
rect 18736 9460 18742 9472
rect 18865 9469 18877 9472
rect 18911 9500 18923 9503
rect 20334 9500 20340 9512
rect 18911 9472 20340 9500
rect 18911 9469 18923 9472
rect 18865 9463 18923 9469
rect 18880 9376 18908 9463
rect 20334 9460 20340 9472
rect 20392 9460 20398 9512
rect 19046 9392 19052 9444
rect 19104 9441 19110 9444
rect 19104 9435 19168 9441
rect 19104 9401 19122 9435
rect 19156 9432 19168 9435
rect 20426 9432 20432 9444
rect 19156 9404 20432 9432
rect 19156 9401 19168 9404
rect 19104 9395 19168 9401
rect 19104 9392 19110 9395
rect 20426 9392 20432 9404
rect 20484 9392 20490 9444
rect 14446 9324 14452 9376
rect 14504 9364 14510 9376
rect 14541 9367 14599 9373
rect 14541 9364 14553 9367
rect 14504 9336 14553 9364
rect 14504 9324 14510 9336
rect 14541 9333 14553 9336
rect 14587 9333 14599 9367
rect 14541 9327 14599 9333
rect 18773 9367 18831 9373
rect 18773 9333 18785 9367
rect 18819 9364 18831 9367
rect 18862 9364 18868 9376
rect 18819 9336 18868 9364
rect 18819 9333 18831 9336
rect 18773 9327 18831 9333
rect 18862 9324 18868 9336
rect 18920 9324 18926 9376
rect 20242 9364 20248 9376
rect 20203 9336 20248 9364
rect 20242 9324 20248 9336
rect 20300 9324 20306 9376
rect 20889 9367 20947 9373
rect 20889 9333 20901 9367
rect 20935 9364 20947 9367
rect 20978 9364 20984 9376
rect 20935 9336 20984 9364
rect 20935 9333 20947 9336
rect 20889 9327 20947 9333
rect 20978 9324 20984 9336
rect 21036 9364 21042 9376
rect 21346 9364 21352 9376
rect 21036 9336 21352 9364
rect 21036 9324 21042 9336
rect 21346 9324 21352 9336
rect 21404 9324 21410 9376
rect 816 9274 26576 9296
rect 816 9222 10027 9274
rect 10079 9222 10091 9274
rect 10143 9222 10155 9274
rect 10207 9222 10219 9274
rect 10271 9222 19360 9274
rect 19412 9222 19424 9274
rect 19476 9222 19488 9274
rect 19540 9222 19552 9274
rect 19604 9222 26576 9274
rect 816 9200 26576 9222
rect 18865 9163 18923 9169
rect 18865 9129 18877 9163
rect 18911 9160 18923 9163
rect 18954 9160 18960 9172
rect 18911 9132 18960 9160
rect 18911 9129 18923 9132
rect 18865 9123 18923 9129
rect 18954 9120 18960 9132
rect 19012 9120 19018 9172
rect 19509 9163 19567 9169
rect 19509 9129 19521 9163
rect 19555 9160 19567 9163
rect 20242 9160 20248 9172
rect 19555 9132 20248 9160
rect 19555 9129 19567 9132
rect 19509 9123 19567 9129
rect 15921 9027 15979 9033
rect 15921 8993 15933 9027
rect 15967 9024 15979 9027
rect 16010 9024 16016 9036
rect 15967 8996 16016 9024
rect 15967 8993 15979 8996
rect 15921 8987 15979 8993
rect 16010 8984 16016 8996
rect 16068 8984 16074 9036
rect 18678 8984 18684 9036
rect 18736 9024 18742 9036
rect 18773 9027 18831 9033
rect 18773 9024 18785 9027
rect 18736 8996 18785 9024
rect 18736 8984 18742 8996
rect 18773 8993 18785 8996
rect 18819 8993 18831 9027
rect 18773 8987 18831 8993
rect 19049 8959 19107 8965
rect 19049 8925 19061 8959
rect 19095 8956 19107 8959
rect 19414 8956 19420 8968
rect 19095 8928 19420 8956
rect 19095 8925 19107 8928
rect 19049 8919 19107 8925
rect 19414 8916 19420 8928
rect 19472 8956 19478 8968
rect 19524 8956 19552 9123
rect 20242 9120 20248 9132
rect 20300 9120 20306 9172
rect 20426 9120 20432 9172
rect 20484 9160 20490 9172
rect 20797 9163 20855 9169
rect 20797 9160 20809 9163
rect 20484 9132 20809 9160
rect 20484 9120 20490 9132
rect 20797 9129 20809 9132
rect 20843 9129 20855 9163
rect 20797 9123 20855 9129
rect 19472 8928 19552 8956
rect 19472 8916 19478 8928
rect 16105 8823 16163 8829
rect 16105 8789 16117 8823
rect 16151 8820 16163 8823
rect 16194 8820 16200 8832
rect 16151 8792 16200 8820
rect 16151 8789 16163 8792
rect 16105 8783 16163 8789
rect 16194 8780 16200 8792
rect 16252 8780 16258 8832
rect 17574 8780 17580 8832
rect 17632 8820 17638 8832
rect 18405 8823 18463 8829
rect 18405 8820 18417 8823
rect 17632 8792 18417 8820
rect 17632 8780 17638 8792
rect 18405 8789 18417 8792
rect 18451 8789 18463 8823
rect 18405 8783 18463 8789
rect 816 8730 26576 8752
rect 816 8678 5360 8730
rect 5412 8678 5424 8730
rect 5476 8678 5488 8730
rect 5540 8678 5552 8730
rect 5604 8678 14694 8730
rect 14746 8678 14758 8730
rect 14810 8678 14822 8730
rect 14874 8678 14886 8730
rect 14938 8678 24027 8730
rect 24079 8678 24091 8730
rect 24143 8678 24155 8730
rect 24207 8678 24219 8730
rect 24271 8678 26576 8730
rect 816 8656 26576 8678
rect 14446 8616 14452 8628
rect 13820 8588 14452 8616
rect 13820 8421 13848 8588
rect 14446 8576 14452 8588
rect 14504 8576 14510 8628
rect 18678 8616 18684 8628
rect 18639 8588 18684 8616
rect 18678 8576 18684 8588
rect 18736 8576 18742 8628
rect 13989 8551 14047 8557
rect 13989 8517 14001 8551
rect 14035 8548 14047 8551
rect 14262 8548 14268 8560
rect 14035 8520 14268 8548
rect 14035 8517 14047 8520
rect 13989 8511 14047 8517
rect 14262 8508 14268 8520
rect 14320 8508 14326 8560
rect 16010 8548 16016 8560
rect 15971 8520 16016 8548
rect 16010 8508 16016 8520
rect 16068 8508 16074 8560
rect 18129 8483 18187 8489
rect 18129 8449 18141 8483
rect 18175 8480 18187 8483
rect 18696 8480 18724 8576
rect 18175 8452 18724 8480
rect 18175 8449 18187 8452
rect 18129 8443 18187 8449
rect 13805 8415 13863 8421
rect 13805 8381 13817 8415
rect 13851 8381 13863 8415
rect 13805 8375 13863 8381
rect 18862 8372 18868 8424
rect 18920 8412 18926 8424
rect 19046 8412 19052 8424
rect 18920 8384 19052 8412
rect 18920 8372 18926 8384
rect 19046 8372 19052 8384
rect 19104 8412 19110 8424
rect 19414 8421 19420 8424
rect 19141 8415 19199 8421
rect 19141 8412 19153 8415
rect 19104 8384 19153 8412
rect 19104 8372 19110 8384
rect 19141 8381 19153 8384
rect 19187 8381 19199 8415
rect 19408 8412 19420 8421
rect 19141 8375 19199 8381
rect 19248 8384 19420 8412
rect 18037 8347 18095 8353
rect 18037 8313 18049 8347
rect 18083 8344 18095 8347
rect 19248 8344 19276 8384
rect 19408 8375 19420 8384
rect 19414 8372 19420 8375
rect 19472 8372 19478 8424
rect 18083 8316 19276 8344
rect 18083 8313 18095 8316
rect 18037 8307 18095 8313
rect 19046 8276 19052 8288
rect 19007 8248 19052 8276
rect 19046 8236 19052 8248
rect 19104 8236 19110 8288
rect 20521 8279 20579 8285
rect 20521 8245 20533 8279
rect 20567 8276 20579 8279
rect 21254 8276 21260 8288
rect 20567 8248 21260 8276
rect 20567 8245 20579 8248
rect 20521 8239 20579 8245
rect 21254 8236 21260 8248
rect 21312 8236 21318 8288
rect 816 8186 26576 8208
rect 816 8134 10027 8186
rect 10079 8134 10091 8186
rect 10143 8134 10155 8186
rect 10207 8134 10219 8186
rect 10271 8134 19360 8186
rect 19412 8134 19424 8186
rect 19476 8134 19488 8186
rect 19540 8134 19552 8186
rect 19604 8134 26576 8186
rect 816 8112 26576 8134
rect 18497 8075 18555 8081
rect 18497 8041 18509 8075
rect 18543 8072 18555 8075
rect 18954 8072 18960 8084
rect 18543 8044 18960 8072
rect 18543 8041 18555 8044
rect 18497 8035 18555 8041
rect 18954 8032 18960 8044
rect 19012 8032 19018 8084
rect 16657 7939 16715 7945
rect 16657 7905 16669 7939
rect 16703 7936 16715 7939
rect 16746 7936 16752 7948
rect 16703 7908 16752 7936
rect 16703 7905 16715 7908
rect 16657 7899 16715 7905
rect 16746 7896 16752 7908
rect 16804 7936 16810 7948
rect 17574 7936 17580 7948
rect 16804 7908 17580 7936
rect 16804 7896 16810 7908
rect 17574 7896 17580 7908
rect 17632 7896 17638 7948
rect 20981 7939 21039 7945
rect 20981 7905 20993 7939
rect 21027 7936 21039 7939
rect 21346 7936 21352 7948
rect 21027 7908 21352 7936
rect 21027 7905 21039 7908
rect 20981 7899 21039 7905
rect 21346 7896 21352 7908
rect 21404 7896 21410 7948
rect 19230 7868 19236 7880
rect 19191 7840 19236 7868
rect 19230 7828 19236 7840
rect 19288 7828 19294 7880
rect 21070 7868 21076 7880
rect 21031 7840 21076 7868
rect 21070 7828 21076 7840
rect 21128 7828 21134 7880
rect 21254 7868 21260 7880
rect 21215 7840 21260 7868
rect 21254 7828 21260 7840
rect 21312 7828 21318 7880
rect 16378 7692 16384 7744
rect 16436 7732 16442 7744
rect 16841 7735 16899 7741
rect 16841 7732 16853 7735
rect 16436 7704 16853 7732
rect 16436 7692 16442 7704
rect 16841 7701 16853 7704
rect 16887 7701 16899 7735
rect 20610 7732 20616 7744
rect 20571 7704 20616 7732
rect 16841 7695 16899 7701
rect 20610 7692 20616 7704
rect 20668 7692 20674 7744
rect 816 7642 26576 7664
rect 816 7590 5360 7642
rect 5412 7590 5424 7642
rect 5476 7590 5488 7642
rect 5540 7590 5552 7642
rect 5604 7590 14694 7642
rect 14746 7590 14758 7642
rect 14810 7590 14822 7642
rect 14874 7590 14886 7642
rect 14938 7590 24027 7642
rect 24079 7590 24091 7642
rect 24143 7590 24155 7642
rect 24207 7590 24219 7642
rect 24271 7590 26576 7642
rect 816 7568 26576 7590
rect 16378 7528 16384 7540
rect 16339 7500 16384 7528
rect 16378 7488 16384 7500
rect 16436 7488 16442 7540
rect 16746 7528 16752 7540
rect 16707 7500 16752 7528
rect 16746 7488 16752 7500
rect 16804 7488 16810 7540
rect 18402 7528 18408 7540
rect 18363 7500 18408 7528
rect 18402 7488 18408 7500
rect 18460 7488 18466 7540
rect 21070 7488 21076 7540
rect 21128 7528 21134 7540
rect 21993 7531 22051 7537
rect 21993 7528 22005 7531
rect 21128 7500 22005 7528
rect 21128 7488 21134 7500
rect 21993 7497 22005 7500
rect 22039 7528 22051 7531
rect 23094 7528 23100 7540
rect 22039 7500 23100 7528
rect 22039 7497 22051 7500
rect 21993 7491 22051 7497
rect 23094 7488 23100 7500
rect 23152 7488 23158 7540
rect 21254 7420 21260 7472
rect 21312 7460 21318 7472
rect 22269 7463 22327 7469
rect 22269 7460 22281 7463
rect 21312 7432 22281 7460
rect 21312 7420 21318 7432
rect 22269 7429 22281 7432
rect 22315 7429 22327 7463
rect 22269 7423 22327 7429
rect 19141 7395 19199 7401
rect 19141 7361 19153 7395
rect 19187 7392 19199 7395
rect 19187 7364 19736 7392
rect 19187 7361 19199 7364
rect 19141 7355 19199 7361
rect 15737 7327 15795 7333
rect 15737 7293 15749 7327
rect 15783 7324 15795 7327
rect 16378 7324 16384 7336
rect 15783 7296 16384 7324
rect 15783 7293 15795 7296
rect 15737 7287 15795 7293
rect 16378 7284 16384 7296
rect 16436 7284 16442 7336
rect 17761 7327 17819 7333
rect 17761 7293 17773 7327
rect 17807 7324 17819 7327
rect 18402 7324 18408 7336
rect 17807 7296 18408 7324
rect 17807 7293 17819 7296
rect 17761 7287 17819 7293
rect 18402 7284 18408 7296
rect 18460 7284 18466 7336
rect 19046 7284 19052 7336
rect 19104 7324 19110 7336
rect 19601 7327 19659 7333
rect 19601 7324 19613 7327
rect 19104 7296 19613 7324
rect 19104 7284 19110 7296
rect 19601 7293 19613 7296
rect 19647 7293 19659 7327
rect 19708 7324 19736 7364
rect 19868 7327 19926 7333
rect 19868 7324 19880 7327
rect 19708 7296 19880 7324
rect 19601 7287 19659 7293
rect 19868 7293 19880 7296
rect 19914 7324 19926 7327
rect 21272 7324 21300 7420
rect 19914 7296 21300 7324
rect 19914 7293 19926 7296
rect 19868 7287 19926 7293
rect 15642 7148 15648 7200
rect 15700 7188 15706 7200
rect 15921 7191 15979 7197
rect 15921 7188 15933 7191
rect 15700 7160 15933 7188
rect 15700 7148 15706 7160
rect 15921 7157 15933 7160
rect 15967 7157 15979 7191
rect 15921 7151 15979 7157
rect 17666 7148 17672 7200
rect 17724 7188 17730 7200
rect 17945 7191 18003 7197
rect 17945 7188 17957 7191
rect 17724 7160 17957 7188
rect 17724 7148 17730 7160
rect 17945 7157 17957 7160
rect 17991 7157 18003 7191
rect 17945 7151 18003 7157
rect 19509 7191 19567 7197
rect 19509 7157 19521 7191
rect 19555 7188 19567 7191
rect 19616 7188 19644 7287
rect 19966 7188 19972 7200
rect 19555 7160 19972 7188
rect 19555 7157 19567 7160
rect 19509 7151 19567 7157
rect 19966 7148 19972 7160
rect 20024 7148 20030 7200
rect 20426 7148 20432 7200
rect 20484 7188 20490 7200
rect 20981 7191 21039 7197
rect 20981 7188 20993 7191
rect 20484 7160 20993 7188
rect 20484 7148 20490 7160
rect 20981 7157 20993 7160
rect 21027 7157 21039 7191
rect 20981 7151 21039 7157
rect 21346 7148 21352 7200
rect 21404 7188 21410 7200
rect 21533 7191 21591 7197
rect 21533 7188 21545 7191
rect 21404 7160 21545 7188
rect 21404 7148 21410 7160
rect 21533 7157 21545 7160
rect 21579 7157 21591 7191
rect 21533 7151 21591 7157
rect 816 7098 26576 7120
rect 816 7046 10027 7098
rect 10079 7046 10091 7098
rect 10143 7046 10155 7098
rect 10207 7046 10219 7098
rect 10271 7046 19360 7098
rect 19412 7046 19424 7098
rect 19476 7046 19488 7098
rect 19540 7046 19552 7098
rect 19604 7046 26576 7098
rect 816 7024 26576 7046
rect 19230 6944 19236 6996
rect 19288 6984 19294 6996
rect 19325 6987 19383 6993
rect 19325 6984 19337 6987
rect 19288 6956 19337 6984
rect 19288 6944 19294 6956
rect 19325 6953 19337 6956
rect 19371 6953 19383 6987
rect 22266 6984 22272 6996
rect 22227 6956 22272 6984
rect 19325 6947 19383 6953
rect 22266 6944 22272 6956
rect 22324 6944 22330 6996
rect 20610 6916 20616 6928
rect 20352 6888 20616 6916
rect 17850 6848 17856 6860
rect 17811 6820 17856 6848
rect 17850 6808 17856 6820
rect 17908 6808 17914 6860
rect 20352 6848 20380 6888
rect 20610 6876 20616 6888
rect 20668 6876 20674 6928
rect 19432 6820 20380 6848
rect 21156 6851 21214 6857
rect 19138 6740 19144 6792
rect 19196 6780 19202 6792
rect 19432 6789 19460 6820
rect 21156 6817 21168 6851
rect 21202 6848 21214 6851
rect 21530 6848 21536 6860
rect 21202 6820 21536 6848
rect 21202 6817 21214 6820
rect 21156 6811 21214 6817
rect 21530 6808 21536 6820
rect 21588 6808 21594 6860
rect 19417 6783 19475 6789
rect 19417 6780 19429 6783
rect 19196 6752 19429 6780
rect 19196 6740 19202 6752
rect 19417 6749 19429 6752
rect 19463 6749 19475 6783
rect 19417 6743 19475 6749
rect 19509 6783 19567 6789
rect 19509 6749 19521 6783
rect 19555 6749 19567 6783
rect 19509 6743 19567 6749
rect 19046 6672 19052 6724
rect 19104 6712 19110 6724
rect 19524 6712 19552 6743
rect 19966 6740 19972 6792
rect 20024 6780 20030 6792
rect 20889 6783 20947 6789
rect 20889 6780 20901 6783
rect 20024 6752 20901 6780
rect 20024 6740 20030 6752
rect 20889 6749 20901 6752
rect 20935 6749 20947 6783
rect 20889 6743 20947 6749
rect 20153 6715 20211 6721
rect 20153 6712 20165 6715
rect 19104 6684 20165 6712
rect 19104 6672 19110 6684
rect 20153 6681 20165 6684
rect 20199 6712 20211 6715
rect 20426 6712 20432 6724
rect 20199 6684 20432 6712
rect 20199 6681 20211 6684
rect 20153 6675 20211 6681
rect 20426 6672 20432 6684
rect 20484 6672 20490 6724
rect 18037 6647 18095 6653
rect 18037 6613 18049 6647
rect 18083 6644 18095 6647
rect 18402 6644 18408 6656
rect 18083 6616 18408 6644
rect 18083 6613 18095 6616
rect 18037 6607 18095 6613
rect 18402 6604 18408 6616
rect 18460 6604 18466 6656
rect 18494 6604 18500 6656
rect 18552 6644 18558 6656
rect 18957 6647 19015 6653
rect 18957 6644 18969 6647
rect 18552 6616 18969 6644
rect 18552 6604 18558 6616
rect 18957 6613 18969 6616
rect 19003 6613 19015 6647
rect 18957 6607 19015 6613
rect 816 6554 26576 6576
rect 816 6502 5360 6554
rect 5412 6502 5424 6554
rect 5476 6502 5488 6554
rect 5540 6502 5552 6554
rect 5604 6502 14694 6554
rect 14746 6502 14758 6554
rect 14810 6502 14822 6554
rect 14874 6502 14886 6554
rect 14938 6502 24027 6554
rect 24079 6502 24091 6554
rect 24143 6502 24155 6554
rect 24207 6502 24219 6554
rect 24271 6502 26576 6554
rect 816 6480 26576 6502
rect 17850 6400 17856 6452
rect 17908 6440 17914 6452
rect 17945 6443 18003 6449
rect 17945 6440 17957 6443
rect 17908 6412 17957 6440
rect 17908 6400 17914 6412
rect 17945 6409 17957 6412
rect 17991 6409 18003 6443
rect 17945 6403 18003 6409
rect 18497 6443 18555 6449
rect 18497 6409 18509 6443
rect 18543 6440 18555 6443
rect 19138 6440 19144 6452
rect 18543 6412 19144 6440
rect 18543 6409 18555 6412
rect 18497 6403 18555 6409
rect 19138 6400 19144 6412
rect 19196 6400 19202 6452
rect 19230 6400 19236 6452
rect 19288 6440 19294 6452
rect 19509 6443 19567 6449
rect 19509 6440 19521 6443
rect 19288 6412 19521 6440
rect 19288 6400 19294 6412
rect 19509 6409 19521 6412
rect 19555 6409 19567 6443
rect 19966 6440 19972 6452
rect 19927 6412 19972 6440
rect 19509 6403 19567 6409
rect 19966 6400 19972 6412
rect 20024 6400 20030 6452
rect 19230 6304 19236 6316
rect 19191 6276 19236 6304
rect 19230 6264 19236 6276
rect 19288 6264 19294 6316
rect 19984 6304 20012 6400
rect 20153 6307 20211 6313
rect 20153 6304 20165 6307
rect 19984 6276 20165 6304
rect 20153 6273 20165 6276
rect 20199 6273 20211 6307
rect 20153 6267 20211 6273
rect 18589 6239 18647 6245
rect 18589 6205 18601 6239
rect 18635 6236 18647 6239
rect 19248 6236 19276 6264
rect 20426 6245 20432 6248
rect 20420 6236 20432 6245
rect 18635 6208 19276 6236
rect 20387 6208 20432 6236
rect 18635 6205 18647 6208
rect 18589 6199 18647 6205
rect 20420 6199 20432 6208
rect 20426 6196 20432 6199
rect 20484 6196 20490 6248
rect 18773 6103 18831 6109
rect 18773 6069 18785 6103
rect 18819 6100 18831 6103
rect 18954 6100 18960 6112
rect 18819 6072 18960 6100
rect 18819 6069 18831 6072
rect 18773 6063 18831 6069
rect 18954 6060 18960 6072
rect 19012 6060 19018 6112
rect 21530 6100 21536 6112
rect 21443 6072 21536 6100
rect 21530 6060 21536 6072
rect 21588 6100 21594 6112
rect 22174 6100 22180 6112
rect 21588 6072 22180 6100
rect 21588 6060 21594 6072
rect 22174 6060 22180 6072
rect 22232 6060 22238 6112
rect 816 6010 26576 6032
rect 816 5958 10027 6010
rect 10079 5958 10091 6010
rect 10143 5958 10155 6010
rect 10207 5958 10219 6010
rect 10271 5958 19360 6010
rect 19412 5958 19424 6010
rect 19476 5958 19488 6010
rect 19540 5958 19552 6010
rect 19604 5958 26576 6010
rect 816 5936 26576 5958
rect 18221 5899 18279 5905
rect 18221 5865 18233 5899
rect 18267 5865 18279 5899
rect 19046 5896 19052 5908
rect 19007 5868 19052 5896
rect 18221 5859 18279 5865
rect 18236 5828 18264 5859
rect 19046 5856 19052 5868
rect 19104 5856 19110 5908
rect 19966 5856 19972 5908
rect 20024 5896 20030 5908
rect 20153 5899 20211 5905
rect 20153 5896 20165 5899
rect 20024 5868 20165 5896
rect 20024 5856 20030 5868
rect 20153 5865 20165 5868
rect 20199 5865 20211 5899
rect 20153 5859 20211 5865
rect 16948 5800 18264 5828
rect 16948 5772 16976 5800
rect 16930 5760 16936 5772
rect 16843 5732 16936 5760
rect 16930 5720 16936 5732
rect 16988 5720 16994 5772
rect 18037 5763 18095 5769
rect 18037 5729 18049 5763
rect 18083 5760 18095 5763
rect 18126 5760 18132 5772
rect 18083 5732 18132 5760
rect 18083 5729 18095 5732
rect 18037 5723 18095 5729
rect 18126 5720 18132 5732
rect 18184 5760 18190 5772
rect 18494 5760 18500 5772
rect 18184 5732 18500 5760
rect 18184 5720 18190 5732
rect 18494 5720 18500 5732
rect 18552 5720 18558 5772
rect 19325 5763 19383 5769
rect 19325 5729 19337 5763
rect 19371 5760 19383 5763
rect 19690 5760 19696 5772
rect 19371 5732 19696 5760
rect 19371 5729 19383 5732
rect 19325 5723 19383 5729
rect 19690 5720 19696 5732
rect 19748 5720 19754 5772
rect 20978 5720 20984 5772
rect 21036 5760 21042 5772
rect 21346 5760 21352 5772
rect 21036 5732 21352 5760
rect 21036 5720 21042 5732
rect 21346 5720 21352 5732
rect 21404 5720 21410 5772
rect 21438 5692 21444 5704
rect 21399 5664 21444 5692
rect 21438 5652 21444 5664
rect 21496 5652 21502 5704
rect 21625 5695 21683 5701
rect 21625 5661 21637 5695
rect 21671 5692 21683 5695
rect 22174 5692 22180 5704
rect 21671 5664 22180 5692
rect 21671 5661 21683 5664
rect 21625 5655 21683 5661
rect 22174 5652 22180 5664
rect 22232 5652 22238 5704
rect 17022 5516 17028 5568
rect 17080 5556 17086 5568
rect 17117 5559 17175 5565
rect 17117 5556 17129 5559
rect 17080 5528 17129 5556
rect 17080 5516 17086 5528
rect 17117 5525 17129 5528
rect 17163 5525 17175 5559
rect 17117 5519 17175 5525
rect 19509 5559 19567 5565
rect 19509 5525 19521 5559
rect 19555 5556 19567 5559
rect 19782 5556 19788 5568
rect 19555 5528 19788 5556
rect 19555 5525 19567 5528
rect 19509 5519 19567 5525
rect 19782 5516 19788 5528
rect 19840 5516 19846 5568
rect 20981 5559 21039 5565
rect 20981 5525 20993 5559
rect 21027 5556 21039 5559
rect 21714 5556 21720 5568
rect 21027 5528 21720 5556
rect 21027 5525 21039 5528
rect 20981 5519 21039 5525
rect 21714 5516 21720 5528
rect 21772 5516 21778 5568
rect 816 5466 26576 5488
rect 816 5414 5360 5466
rect 5412 5414 5424 5466
rect 5476 5414 5488 5466
rect 5540 5414 5552 5466
rect 5604 5414 14694 5466
rect 14746 5414 14758 5466
rect 14810 5414 14822 5466
rect 14874 5414 14886 5466
rect 14938 5414 24027 5466
rect 24079 5414 24091 5466
rect 24143 5414 24155 5466
rect 24207 5414 24219 5466
rect 24271 5414 26576 5466
rect 816 5392 26576 5414
rect 16930 5352 16936 5364
rect 16891 5324 16936 5352
rect 16930 5312 16936 5324
rect 16988 5312 16994 5364
rect 18126 5352 18132 5364
rect 18087 5324 18132 5352
rect 18126 5312 18132 5324
rect 18184 5312 18190 5364
rect 19417 5355 19475 5361
rect 19417 5321 19429 5355
rect 19463 5352 19475 5355
rect 19690 5352 19696 5364
rect 19463 5324 19696 5352
rect 19463 5321 19475 5324
rect 19417 5315 19475 5321
rect 19690 5312 19696 5324
rect 19748 5312 19754 5364
rect 22174 5312 22180 5364
rect 22232 5352 22238 5364
rect 22269 5355 22327 5361
rect 22269 5352 22281 5355
rect 22232 5324 22281 5352
rect 22232 5312 22238 5324
rect 22269 5321 22281 5324
rect 22315 5321 22327 5355
rect 22269 5315 22327 5321
rect 21714 5216 21720 5228
rect 21675 5188 21720 5216
rect 21714 5176 21720 5188
rect 21772 5176 21778 5228
rect 21806 5176 21812 5228
rect 21864 5216 21870 5228
rect 21901 5219 21959 5225
rect 21901 5216 21913 5219
rect 21864 5188 21913 5216
rect 21864 5176 21870 5188
rect 21901 5185 21913 5188
rect 21947 5216 21959 5219
rect 22266 5216 22272 5228
rect 21947 5188 22272 5216
rect 21947 5185 21959 5188
rect 21901 5179 21959 5185
rect 22266 5176 22272 5188
rect 22324 5176 22330 5228
rect 20245 5083 20303 5089
rect 20245 5049 20257 5083
rect 20291 5080 20303 5083
rect 21622 5080 21628 5092
rect 20291 5052 21628 5080
rect 20291 5049 20303 5052
rect 20245 5043 20303 5049
rect 21622 5040 21628 5052
rect 21680 5040 21686 5092
rect 20150 5012 20156 5024
rect 20111 4984 20156 5012
rect 20150 4972 20156 4984
rect 20208 4972 20214 5024
rect 20978 5012 20984 5024
rect 20939 4984 20984 5012
rect 20978 4972 20984 4984
rect 21036 4972 21042 5024
rect 21254 5012 21260 5024
rect 21215 4984 21260 5012
rect 21254 4972 21260 4984
rect 21312 4972 21318 5024
rect 816 4922 26576 4944
rect 816 4870 10027 4922
rect 10079 4870 10091 4922
rect 10143 4870 10155 4922
rect 10207 4870 10219 4922
rect 10271 4870 19360 4922
rect 19412 4870 19424 4922
rect 19476 4870 19488 4922
rect 19540 4870 19552 4922
rect 19604 4870 26576 4922
rect 816 4848 26576 4870
rect 21622 4808 21628 4820
rect 21583 4780 21628 4808
rect 21622 4768 21628 4780
rect 21680 4768 21686 4820
rect 21714 4768 21720 4820
rect 21772 4808 21778 4820
rect 21993 4811 22051 4817
rect 21993 4808 22005 4811
rect 21772 4780 22005 4808
rect 21772 4768 21778 4780
rect 21993 4777 22005 4780
rect 22039 4777 22051 4811
rect 21993 4771 22051 4777
rect 21349 4743 21407 4749
rect 21349 4709 21361 4743
rect 21395 4740 21407 4743
rect 21806 4740 21812 4752
rect 21395 4712 21812 4740
rect 21395 4709 21407 4712
rect 21349 4703 21407 4709
rect 21806 4700 21812 4712
rect 21864 4700 21870 4752
rect 20610 4632 20616 4684
rect 20668 4672 20674 4684
rect 20705 4675 20763 4681
rect 20705 4672 20717 4675
rect 20668 4644 20717 4672
rect 20668 4632 20674 4644
rect 20705 4641 20717 4644
rect 20751 4672 20763 4675
rect 21254 4672 21260 4684
rect 20751 4644 21260 4672
rect 20751 4641 20763 4644
rect 20705 4635 20763 4641
rect 21254 4632 21260 4644
rect 21312 4632 21318 4684
rect 24290 4672 24296 4684
rect 24251 4644 24296 4672
rect 24290 4632 24296 4644
rect 24348 4632 24354 4684
rect 20889 4539 20947 4545
rect 20889 4505 20901 4539
rect 20935 4536 20947 4539
rect 21806 4536 21812 4548
rect 20935 4508 21812 4536
rect 20935 4505 20947 4508
rect 20889 4499 20947 4505
rect 21806 4496 21812 4508
rect 21864 4496 21870 4548
rect 23186 4428 23192 4480
rect 23244 4468 23250 4480
rect 24477 4471 24535 4477
rect 24477 4468 24489 4471
rect 23244 4440 24489 4468
rect 23244 4428 23250 4440
rect 24477 4437 24489 4440
rect 24523 4437 24535 4471
rect 24477 4431 24535 4437
rect 816 4378 26576 4400
rect 816 4326 5360 4378
rect 5412 4326 5424 4378
rect 5476 4326 5488 4378
rect 5540 4326 5552 4378
rect 5604 4326 14694 4378
rect 14746 4326 14758 4378
rect 14810 4326 14822 4378
rect 14874 4326 14886 4378
rect 14938 4326 24027 4378
rect 24079 4326 24091 4378
rect 24143 4326 24155 4378
rect 24207 4326 24219 4378
rect 24271 4326 26576 4378
rect 816 4304 26576 4326
rect 20610 4264 20616 4276
rect 20571 4236 20616 4264
rect 20610 4224 20616 4236
rect 20668 4224 20674 4276
rect 24201 4267 24259 4273
rect 24201 4233 24213 4267
rect 24247 4264 24259 4267
rect 24382 4264 24388 4276
rect 24247 4236 24388 4264
rect 24247 4233 24259 4236
rect 24201 4227 24259 4233
rect 24382 4224 24388 4236
rect 24440 4224 24446 4276
rect 21349 4131 21407 4137
rect 21349 4128 21361 4131
rect 20720 4100 21361 4128
rect 20720 4069 20748 4100
rect 21349 4097 21361 4100
rect 21395 4128 21407 4131
rect 21530 4128 21536 4140
rect 21395 4100 21536 4128
rect 21395 4097 21407 4100
rect 21349 4091 21407 4097
rect 21530 4088 21536 4100
rect 21588 4088 21594 4140
rect 20705 4063 20763 4069
rect 20705 4029 20717 4063
rect 20751 4029 20763 4063
rect 20705 4023 20763 4029
rect 21806 4020 21812 4072
rect 21864 4060 21870 4072
rect 22361 4063 22419 4069
rect 22361 4060 22373 4063
rect 21864 4032 22373 4060
rect 21864 4020 21870 4032
rect 22361 4029 22373 4032
rect 22407 4029 22419 4063
rect 22361 4023 22419 4029
rect 23922 4020 23928 4072
rect 23980 4060 23986 4072
rect 24293 4063 24351 4069
rect 24293 4060 24305 4063
rect 23980 4032 24305 4060
rect 23980 4020 23986 4032
rect 24293 4029 24305 4032
rect 24339 4060 24351 4063
rect 24845 4063 24903 4069
rect 24845 4060 24857 4063
rect 24339 4032 24857 4060
rect 24339 4029 24351 4032
rect 24293 4023 24351 4029
rect 24845 4029 24857 4032
rect 24891 4029 24903 4063
rect 24845 4023 24903 4029
rect 22450 3992 22456 4004
rect 22008 3964 22456 3992
rect 20889 3927 20947 3933
rect 20889 3893 20901 3927
rect 20935 3924 20947 3927
rect 21070 3924 21076 3936
rect 20935 3896 21076 3924
rect 20935 3893 20947 3896
rect 20889 3887 20947 3893
rect 21070 3884 21076 3896
rect 21128 3884 21134 3936
rect 22008 3933 22036 3964
rect 22450 3952 22456 3964
rect 22508 3952 22514 4004
rect 21993 3927 22051 3933
rect 21993 3893 22005 3927
rect 22039 3893 22051 3927
rect 24474 3924 24480 3936
rect 24435 3896 24480 3924
rect 21993 3887 22051 3893
rect 24474 3884 24480 3896
rect 24532 3884 24538 3936
rect 816 3834 26576 3856
rect 816 3782 10027 3834
rect 10079 3782 10091 3834
rect 10143 3782 10155 3834
rect 10207 3782 10219 3834
rect 10271 3782 19360 3834
rect 19412 3782 19424 3834
rect 19476 3782 19488 3834
rect 19540 3782 19552 3834
rect 19604 3782 26576 3834
rect 816 3760 26576 3782
rect 24293 3587 24351 3593
rect 24293 3553 24305 3587
rect 24339 3584 24351 3587
rect 24382 3584 24388 3596
rect 24339 3556 24388 3584
rect 24339 3553 24351 3556
rect 24293 3547 24351 3553
rect 24382 3544 24388 3556
rect 24440 3544 24446 3596
rect 8006 3476 8012 3528
rect 8064 3516 8070 3528
rect 8834 3516 8840 3528
rect 8064 3488 8840 3516
rect 8064 3476 8070 3488
rect 8834 3476 8840 3488
rect 8892 3476 8898 3528
rect 10766 3476 10772 3528
rect 10824 3516 10830 3528
rect 11594 3516 11600 3528
rect 10824 3488 11600 3516
rect 10824 3476 10830 3488
rect 11594 3476 11600 3488
rect 11652 3476 11658 3528
rect 12238 3476 12244 3528
rect 12296 3516 12302 3528
rect 12698 3516 12704 3528
rect 12296 3488 12704 3516
rect 12296 3476 12302 3488
rect 12698 3476 12704 3488
rect 12756 3476 12762 3528
rect 12882 3476 12888 3528
rect 12940 3516 12946 3528
rect 13434 3516 13440 3528
rect 12940 3488 13440 3516
rect 12940 3476 12946 3488
rect 13434 3476 13440 3488
rect 13492 3476 13498 3528
rect 23646 3380 23652 3392
rect 23607 3352 23652 3380
rect 23646 3340 23652 3352
rect 23704 3340 23710 3392
rect 24477 3383 24535 3389
rect 24477 3349 24489 3383
rect 24523 3380 24535 3383
rect 25210 3380 25216 3392
rect 24523 3352 25216 3380
rect 24523 3349 24535 3352
rect 24477 3343 24535 3349
rect 25210 3340 25216 3352
rect 25268 3340 25274 3392
rect 816 3290 26576 3312
rect 816 3238 5360 3290
rect 5412 3238 5424 3290
rect 5476 3238 5488 3290
rect 5540 3238 5552 3290
rect 5604 3238 14694 3290
rect 14746 3238 14758 3290
rect 14810 3238 14822 3290
rect 14874 3238 14886 3290
rect 14938 3238 24027 3290
rect 24079 3238 24091 3290
rect 24143 3238 24155 3290
rect 24207 3238 24219 3290
rect 24271 3238 26576 3290
rect 816 3216 26576 3238
rect 21806 3136 21812 3188
rect 21864 3176 21870 3188
rect 23094 3176 23100 3188
rect 21864 3148 23100 3176
rect 21864 3136 21870 3148
rect 23094 3136 23100 3148
rect 23152 3136 23158 3188
rect 24382 3176 24388 3188
rect 24343 3148 24388 3176
rect 24382 3136 24388 3148
rect 24440 3136 24446 3188
rect 23646 2972 23652 2984
rect 23607 2944 23652 2972
rect 23646 2932 23652 2944
rect 23704 2932 23710 2984
rect 24753 2975 24811 2981
rect 24753 2941 24765 2975
rect 24799 2972 24811 2975
rect 24799 2944 25348 2972
rect 24799 2941 24811 2944
rect 24753 2935 24811 2941
rect 25320 2848 25348 2944
rect 23830 2836 23836 2848
rect 23791 2808 23836 2836
rect 23830 2796 23836 2808
rect 23888 2796 23894 2848
rect 24474 2796 24480 2848
rect 24532 2836 24538 2848
rect 24937 2839 24995 2845
rect 24937 2836 24949 2839
rect 24532 2808 24949 2836
rect 24532 2796 24538 2808
rect 24937 2805 24949 2808
rect 24983 2805 24995 2839
rect 25302 2836 25308 2848
rect 25263 2808 25308 2836
rect 24937 2799 24995 2805
rect 25302 2796 25308 2808
rect 25360 2796 25366 2848
rect 816 2746 26576 2768
rect 816 2694 10027 2746
rect 10079 2694 10091 2746
rect 10143 2694 10155 2746
rect 10207 2694 10219 2746
rect 10271 2694 19360 2746
rect 19412 2694 19424 2746
rect 19476 2694 19488 2746
rect 19540 2694 19552 2746
rect 19604 2694 26576 2746
rect 816 2672 26576 2694
rect 21533 2635 21591 2641
rect 21533 2601 21545 2635
rect 21579 2632 21591 2635
rect 21622 2632 21628 2644
rect 21579 2604 21628 2632
rect 21579 2601 21591 2604
rect 21533 2595 21591 2601
rect 20889 2499 20947 2505
rect 20889 2465 20901 2499
rect 20935 2496 20947 2499
rect 21548 2496 21576 2595
rect 21622 2592 21628 2604
rect 21680 2592 21686 2644
rect 22726 2632 22732 2644
rect 22687 2604 22732 2632
rect 22726 2592 22732 2604
rect 22784 2592 22790 2644
rect 24382 2592 24388 2644
rect 24440 2632 24446 2644
rect 24845 2635 24903 2641
rect 24845 2632 24857 2635
rect 24440 2604 24857 2632
rect 24440 2592 24446 2604
rect 24845 2601 24857 2604
rect 24891 2601 24903 2635
rect 24845 2595 24903 2601
rect 20935 2468 21576 2496
rect 22545 2499 22603 2505
rect 20935 2465 20947 2468
rect 20889 2459 20947 2465
rect 22545 2465 22557 2499
rect 22591 2465 22603 2499
rect 22545 2459 22603 2465
rect 24293 2499 24351 2505
rect 24293 2465 24305 2499
rect 24339 2496 24351 2499
rect 24400 2496 24428 2592
rect 24339 2468 24428 2496
rect 24339 2465 24351 2468
rect 24293 2459 24351 2465
rect 22560 2428 22588 2459
rect 23189 2431 23247 2437
rect 23189 2428 23201 2431
rect 22560 2400 23201 2428
rect 23189 2397 23201 2400
rect 23235 2428 23247 2431
rect 23278 2428 23284 2440
rect 23235 2400 23284 2428
rect 23235 2397 23247 2400
rect 23189 2391 23247 2397
rect 23278 2388 23284 2400
rect 23336 2388 23342 2440
rect 20426 2252 20432 2304
rect 20484 2292 20490 2304
rect 21073 2295 21131 2301
rect 21073 2292 21085 2295
rect 20484 2264 21085 2292
rect 20484 2252 20490 2264
rect 21073 2261 21085 2264
rect 21119 2261 21131 2295
rect 21073 2255 21131 2261
rect 23186 2252 23192 2304
rect 23244 2292 23250 2304
rect 24477 2295 24535 2301
rect 24477 2292 24489 2295
rect 23244 2264 24489 2292
rect 23244 2252 23250 2264
rect 24477 2261 24489 2264
rect 24523 2261 24535 2295
rect 24477 2255 24535 2261
rect 816 2202 26576 2224
rect 816 2150 5360 2202
rect 5412 2150 5424 2202
rect 5476 2150 5488 2202
rect 5540 2150 5552 2202
rect 5604 2150 14694 2202
rect 14746 2150 14758 2202
rect 14810 2150 14822 2202
rect 14874 2150 14886 2202
rect 14938 2150 24027 2202
rect 24079 2150 24091 2202
rect 24143 2150 24155 2202
rect 24207 2150 24219 2202
rect 24271 2150 26576 2202
rect 816 2128 26576 2150
rect 7270 552 7276 604
rect 7328 592 7334 604
rect 7454 592 7460 604
rect 7328 564 7460 592
rect 7328 552 7334 564
rect 7454 552 7460 564
rect 7512 552 7518 604
rect 8098 552 8104 604
rect 8156 592 8162 604
rect 8466 592 8472 604
rect 8156 564 8472 592
rect 8156 552 8162 564
rect 8466 552 8472 564
rect 8524 552 8530 604
rect 13618 552 13624 604
rect 13676 592 13682 604
rect 13802 592 13808 604
rect 13676 564 13808 592
rect 13676 552 13682 564
rect 13802 552 13808 564
rect 13860 552 13866 604
<< via1 >>
rect 19236 26324 19288 26376
rect 23836 26324 23888 26376
rect 13716 26256 13768 26308
rect 24480 26256 24532 26308
rect 10027 25542 10079 25594
rect 10091 25542 10143 25594
rect 10155 25542 10207 25594
rect 10219 25542 10271 25594
rect 19360 25542 19412 25594
rect 19424 25542 19476 25594
rect 19488 25542 19540 25594
rect 19552 25542 19604 25594
rect 5360 24998 5412 25050
rect 5424 24998 5476 25050
rect 5488 24998 5540 25050
rect 5552 24998 5604 25050
rect 14694 24998 14746 25050
rect 14758 24998 14810 25050
rect 14822 24998 14874 25050
rect 14886 24998 14938 25050
rect 24027 24998 24079 25050
rect 24091 24998 24143 25050
rect 24155 24998 24207 25050
rect 24219 24998 24271 25050
rect 11232 24896 11284 24948
rect 23836 24896 23888 24948
rect 10680 24828 10732 24880
rect 24480 24828 24532 24880
rect 10027 24454 10079 24506
rect 10091 24454 10143 24506
rect 10155 24454 10207 24506
rect 10219 24454 10271 24506
rect 19360 24454 19412 24506
rect 19424 24454 19476 24506
rect 19488 24454 19540 24506
rect 19552 24454 19604 24506
rect 5360 23910 5412 23962
rect 5424 23910 5476 23962
rect 5488 23910 5540 23962
rect 5552 23910 5604 23962
rect 14694 23910 14746 23962
rect 14758 23910 14810 23962
rect 14822 23910 14874 23962
rect 14886 23910 14938 23962
rect 24027 23910 24079 23962
rect 24091 23910 24143 23962
rect 24155 23910 24207 23962
rect 24219 23910 24271 23962
rect 10027 23366 10079 23418
rect 10091 23366 10143 23418
rect 10155 23366 10207 23418
rect 10219 23366 10271 23418
rect 19360 23366 19412 23418
rect 19424 23366 19476 23418
rect 19488 23366 19540 23418
rect 19552 23366 19604 23418
rect 1848 23171 1900 23180
rect 1848 23137 1857 23171
rect 1857 23137 1891 23171
rect 1891 23137 1900 23171
rect 1848 23128 1900 23137
rect 2032 23035 2084 23044
rect 2032 23001 2041 23035
rect 2041 23001 2075 23035
rect 2075 23001 2084 23035
rect 2032 22992 2084 23001
rect 14452 22924 14504 22976
rect 15096 22924 15148 22976
rect 5360 22822 5412 22874
rect 5424 22822 5476 22874
rect 5488 22822 5540 22874
rect 5552 22822 5604 22874
rect 14694 22822 14746 22874
rect 14758 22822 14810 22874
rect 14822 22822 14874 22874
rect 14886 22822 14938 22874
rect 24027 22822 24079 22874
rect 24091 22822 24143 22874
rect 24155 22822 24207 22874
rect 24219 22822 24271 22874
rect 2492 22559 2544 22568
rect 2492 22525 2501 22559
rect 2501 22525 2535 22559
rect 2535 22525 2544 22559
rect 2492 22516 2544 22525
rect 1848 22423 1900 22432
rect 1848 22389 1857 22423
rect 1857 22389 1891 22423
rect 1891 22389 1900 22423
rect 1848 22380 1900 22389
rect 2676 22423 2728 22432
rect 2676 22389 2685 22423
rect 2685 22389 2719 22423
rect 2719 22389 2728 22423
rect 2676 22380 2728 22389
rect 10027 22278 10079 22330
rect 10091 22278 10143 22330
rect 10155 22278 10207 22330
rect 10219 22278 10271 22330
rect 19360 22278 19412 22330
rect 19424 22278 19476 22330
rect 19488 22278 19540 22330
rect 19552 22278 19604 22330
rect 3780 22083 3832 22092
rect 3780 22049 3789 22083
rect 3789 22049 3823 22083
rect 3823 22049 3832 22083
rect 3780 22040 3832 22049
rect 3964 21947 4016 21956
rect 3964 21913 3973 21947
rect 3973 21913 4007 21947
rect 4007 21913 4016 21947
rect 3964 21904 4016 21913
rect 5360 21734 5412 21786
rect 5424 21734 5476 21786
rect 5488 21734 5540 21786
rect 5552 21734 5604 21786
rect 14694 21734 14746 21786
rect 14758 21734 14810 21786
rect 14822 21734 14874 21786
rect 14886 21734 14938 21786
rect 24027 21734 24079 21786
rect 24091 21734 24143 21786
rect 24155 21734 24207 21786
rect 24219 21734 24271 21786
rect 4056 21675 4108 21684
rect 4056 21641 4065 21675
rect 4065 21641 4099 21675
rect 4099 21641 4108 21675
rect 4056 21632 4108 21641
rect 3780 21496 3832 21548
rect 3872 21292 3924 21344
rect 10027 21190 10079 21242
rect 10091 21190 10143 21242
rect 10155 21190 10207 21242
rect 10219 21190 10271 21242
rect 19360 21190 19412 21242
rect 19424 21190 19476 21242
rect 19488 21190 19540 21242
rect 19552 21190 19604 21242
rect 5360 20646 5412 20698
rect 5424 20646 5476 20698
rect 5488 20646 5540 20698
rect 5552 20646 5604 20698
rect 14694 20646 14746 20698
rect 14758 20646 14810 20698
rect 14822 20646 14874 20698
rect 14886 20646 14938 20698
rect 24027 20646 24079 20698
rect 24091 20646 24143 20698
rect 24155 20646 24207 20698
rect 24219 20646 24271 20698
rect 10027 20102 10079 20154
rect 10091 20102 10143 20154
rect 10155 20102 10207 20154
rect 10219 20102 10271 20154
rect 19360 20102 19412 20154
rect 19424 20102 19476 20154
rect 19488 20102 19540 20154
rect 19552 20102 19604 20154
rect 5712 20000 5764 20052
rect 5252 19907 5304 19916
rect 5252 19873 5261 19907
rect 5261 19873 5295 19907
rect 5295 19873 5304 19907
rect 5252 19864 5304 19873
rect 5360 19558 5412 19610
rect 5424 19558 5476 19610
rect 5488 19558 5540 19610
rect 5552 19558 5604 19610
rect 14694 19558 14746 19610
rect 14758 19558 14810 19610
rect 14822 19558 14874 19610
rect 14886 19558 14938 19610
rect 24027 19558 24079 19610
rect 24091 19558 24143 19610
rect 24155 19558 24207 19610
rect 24219 19558 24271 19610
rect 6540 19295 6592 19304
rect 6540 19261 6549 19295
rect 6549 19261 6583 19295
rect 6583 19261 6592 19295
rect 6540 19252 6592 19261
rect 21996 19252 22048 19304
rect 22180 19252 22232 19304
rect 5252 19159 5304 19168
rect 5252 19125 5261 19159
rect 5261 19125 5295 19159
rect 5295 19125 5304 19159
rect 5252 19116 5304 19125
rect 6724 19159 6776 19168
rect 6724 19125 6733 19159
rect 6733 19125 6767 19159
rect 6767 19125 6776 19159
rect 6724 19116 6776 19125
rect 10027 19014 10079 19066
rect 10091 19014 10143 19066
rect 10155 19014 10207 19066
rect 10219 19014 10271 19066
rect 19360 19014 19412 19066
rect 19424 19014 19476 19066
rect 19488 19014 19540 19066
rect 19552 19014 19604 19066
rect 6816 18955 6868 18964
rect 6816 18921 6825 18955
rect 6825 18921 6859 18955
rect 6859 18921 6868 18955
rect 6816 18912 6868 18921
rect 6724 18776 6776 18828
rect 5360 18470 5412 18522
rect 5424 18470 5476 18522
rect 5488 18470 5540 18522
rect 5552 18470 5604 18522
rect 14694 18470 14746 18522
rect 14758 18470 14810 18522
rect 14822 18470 14874 18522
rect 14886 18470 14938 18522
rect 24027 18470 24079 18522
rect 24091 18470 24143 18522
rect 24155 18470 24207 18522
rect 24219 18470 24271 18522
rect 6724 18071 6776 18080
rect 6724 18037 6733 18071
rect 6733 18037 6767 18071
rect 6767 18037 6776 18071
rect 6724 18028 6776 18037
rect 10027 17926 10079 17978
rect 10091 17926 10143 17978
rect 10155 17926 10207 17978
rect 10219 17926 10271 17978
rect 19360 17926 19412 17978
rect 19424 17926 19476 17978
rect 19488 17926 19540 17978
rect 19552 17926 19604 17978
rect 10680 17867 10732 17876
rect 10680 17833 10689 17867
rect 10689 17833 10723 17867
rect 10723 17833 10732 17867
rect 10680 17824 10732 17833
rect 7276 17731 7328 17740
rect 7276 17697 7285 17731
rect 7285 17697 7319 17731
rect 7319 17697 7328 17731
rect 7276 17688 7328 17697
rect 10496 17731 10548 17740
rect 10496 17697 10505 17731
rect 10505 17697 10539 17731
rect 10539 17697 10548 17731
rect 10496 17688 10548 17697
rect 7460 17595 7512 17604
rect 7460 17561 7469 17595
rect 7469 17561 7503 17595
rect 7503 17561 7512 17595
rect 7460 17552 7512 17561
rect 5360 17382 5412 17434
rect 5424 17382 5476 17434
rect 5488 17382 5540 17434
rect 5552 17382 5604 17434
rect 14694 17382 14746 17434
rect 14758 17382 14810 17434
rect 14822 17382 14874 17434
rect 14886 17382 14938 17434
rect 24027 17382 24079 17434
rect 24091 17382 24143 17434
rect 24155 17382 24207 17434
rect 24219 17382 24271 17434
rect 7276 16983 7328 16992
rect 7276 16949 7285 16983
rect 7285 16949 7319 16983
rect 7319 16949 7328 16983
rect 7276 16940 7328 16949
rect 8104 16983 8156 16992
rect 8104 16949 8113 16983
rect 8113 16949 8147 16983
rect 8147 16949 8156 16983
rect 8104 16940 8156 16949
rect 8472 16983 8524 16992
rect 8472 16949 8481 16983
rect 8481 16949 8515 16983
rect 8515 16949 8524 16983
rect 8472 16940 8524 16949
rect 10496 16983 10548 16992
rect 10496 16949 10505 16983
rect 10505 16949 10539 16983
rect 10539 16949 10548 16983
rect 10496 16940 10548 16949
rect 10027 16838 10079 16890
rect 10091 16838 10143 16890
rect 10155 16838 10207 16890
rect 10219 16838 10271 16890
rect 19360 16838 19412 16890
rect 19424 16838 19476 16890
rect 19488 16838 19540 16890
rect 19552 16838 19604 16890
rect 9576 16779 9628 16788
rect 9576 16745 9585 16779
rect 9585 16745 9619 16779
rect 9619 16745 9628 16779
rect 9576 16736 9628 16745
rect 9852 16600 9904 16652
rect 5360 16294 5412 16346
rect 5424 16294 5476 16346
rect 5488 16294 5540 16346
rect 5552 16294 5604 16346
rect 14694 16294 14746 16346
rect 14758 16294 14810 16346
rect 14822 16294 14874 16346
rect 14886 16294 14938 16346
rect 24027 16294 24079 16346
rect 24091 16294 24143 16346
rect 24155 16294 24207 16346
rect 24219 16294 24271 16346
rect 9484 16235 9536 16244
rect 9484 16201 9493 16235
rect 9493 16201 9527 16235
rect 9527 16201 9536 16235
rect 9484 16192 9536 16201
rect 13716 16192 13768 16244
rect 9300 15852 9352 15904
rect 9852 15895 9904 15904
rect 9852 15861 9861 15895
rect 9861 15861 9895 15895
rect 9895 15861 9904 15895
rect 9852 15852 9904 15861
rect 13808 15852 13860 15904
rect 10027 15750 10079 15802
rect 10091 15750 10143 15802
rect 10155 15750 10207 15802
rect 10219 15750 10271 15802
rect 19360 15750 19412 15802
rect 19424 15750 19476 15802
rect 19488 15750 19540 15802
rect 19552 15750 19604 15802
rect 5360 15206 5412 15258
rect 5424 15206 5476 15258
rect 5488 15206 5540 15258
rect 5552 15206 5604 15258
rect 14694 15206 14746 15258
rect 14758 15206 14810 15258
rect 14822 15206 14874 15258
rect 14886 15206 14938 15258
rect 24027 15206 24079 15258
rect 24091 15206 24143 15258
rect 24155 15206 24207 15258
rect 24219 15206 24271 15258
rect 10864 15147 10916 15156
rect 10864 15113 10873 15147
rect 10873 15113 10907 15147
rect 10907 15113 10916 15147
rect 10864 15104 10916 15113
rect 17948 15147 18000 15156
rect 17948 15113 17957 15147
rect 17957 15113 17991 15147
rect 17991 15113 18000 15147
rect 17948 15104 18000 15113
rect 19696 15104 19748 15156
rect 15648 14832 15700 14884
rect 19696 14900 19748 14952
rect 11140 14764 11192 14816
rect 10027 14662 10079 14714
rect 10091 14662 10143 14714
rect 10155 14662 10207 14714
rect 10219 14662 10271 14714
rect 19360 14662 19412 14714
rect 19424 14662 19476 14714
rect 19488 14662 19540 14714
rect 19552 14662 19604 14714
rect 11232 14603 11284 14612
rect 11232 14569 11241 14603
rect 11241 14569 11275 14603
rect 11275 14569 11284 14603
rect 11232 14560 11284 14569
rect 15648 14603 15700 14612
rect 15648 14569 15657 14603
rect 15657 14569 15691 14603
rect 15691 14569 15700 14603
rect 15648 14560 15700 14569
rect 12520 14492 12572 14544
rect 13348 14492 13400 14544
rect 19696 14560 19748 14612
rect 24480 14603 24532 14612
rect 24480 14569 24489 14603
rect 24489 14569 24523 14603
rect 24523 14569 24532 14603
rect 24480 14560 24532 14569
rect 19236 14492 19288 14544
rect 11048 14467 11100 14476
rect 11048 14433 11057 14467
rect 11057 14433 11091 14467
rect 11091 14433 11100 14467
rect 11048 14424 11100 14433
rect 16292 14424 16344 14476
rect 18132 14467 18184 14476
rect 18132 14433 18141 14467
rect 18141 14433 18175 14467
rect 18175 14433 18184 14467
rect 18132 14424 18184 14433
rect 24388 14424 24440 14476
rect 12428 14399 12480 14408
rect 12428 14365 12437 14399
rect 12437 14365 12471 14399
rect 12471 14365 12480 14399
rect 12428 14356 12480 14365
rect 16108 14399 16160 14408
rect 16108 14365 16117 14399
rect 16117 14365 16151 14399
rect 16151 14365 16160 14399
rect 16108 14356 16160 14365
rect 16200 14399 16252 14408
rect 16200 14365 16209 14399
rect 16209 14365 16243 14399
rect 16243 14365 16252 14399
rect 16200 14356 16252 14365
rect 17764 14356 17816 14408
rect 14176 14220 14228 14272
rect 18776 14263 18828 14272
rect 18776 14229 18785 14263
rect 18785 14229 18819 14263
rect 18819 14229 18828 14263
rect 18776 14220 18828 14229
rect 5360 14118 5412 14170
rect 5424 14118 5476 14170
rect 5488 14118 5540 14170
rect 5552 14118 5604 14170
rect 14694 14118 14746 14170
rect 14758 14118 14810 14170
rect 14822 14118 14874 14170
rect 14886 14118 14938 14170
rect 24027 14118 24079 14170
rect 24091 14118 24143 14170
rect 24155 14118 24207 14170
rect 24219 14118 24271 14170
rect 12520 14059 12572 14068
rect 12520 14025 12529 14059
rect 12529 14025 12563 14059
rect 12563 14025 12572 14059
rect 12520 14016 12572 14025
rect 18132 14016 18184 14068
rect 11048 13855 11100 13864
rect 11048 13821 11057 13855
rect 11057 13821 11091 13855
rect 11091 13821 11100 13855
rect 11048 13812 11100 13821
rect 14268 13855 14320 13864
rect 14268 13821 14277 13855
rect 14277 13821 14311 13855
rect 14311 13821 14320 13855
rect 14268 13812 14320 13821
rect 14360 13812 14412 13864
rect 16108 13880 16160 13932
rect 17672 13880 17724 13932
rect 16292 13855 16344 13864
rect 16292 13821 16301 13855
rect 16301 13821 16335 13855
rect 16335 13821 16344 13855
rect 16292 13812 16344 13821
rect 12796 13787 12848 13796
rect 12796 13753 12805 13787
rect 12805 13753 12839 13787
rect 12839 13753 12848 13787
rect 12796 13744 12848 13753
rect 13900 13744 13952 13796
rect 15740 13744 15792 13796
rect 18776 13744 18828 13796
rect 19052 13744 19104 13796
rect 15648 13719 15700 13728
rect 15648 13685 15657 13719
rect 15657 13685 15691 13719
rect 15691 13685 15700 13719
rect 15648 13676 15700 13685
rect 19788 13719 19840 13728
rect 19788 13685 19797 13719
rect 19797 13685 19831 13719
rect 19831 13685 19840 13719
rect 19788 13676 19840 13685
rect 24296 13719 24348 13728
rect 24296 13685 24305 13719
rect 24305 13685 24339 13719
rect 24339 13685 24348 13719
rect 24296 13676 24348 13685
rect 10027 13574 10079 13626
rect 10091 13574 10143 13626
rect 10155 13574 10207 13626
rect 10219 13574 10271 13626
rect 19360 13574 19412 13626
rect 19424 13574 19476 13626
rect 19488 13574 19540 13626
rect 19552 13574 19604 13626
rect 13900 13472 13952 13524
rect 15648 13472 15700 13524
rect 16200 13472 16252 13524
rect 18776 13515 18828 13524
rect 18776 13481 18785 13515
rect 18785 13481 18819 13515
rect 18819 13481 18828 13515
rect 18776 13472 18828 13481
rect 19236 13472 19288 13524
rect 24296 13472 24348 13524
rect 12796 13404 12848 13456
rect 12520 13336 12572 13388
rect 14176 13336 14228 13388
rect 15372 13379 15424 13388
rect 15372 13345 15381 13379
rect 15381 13345 15415 13379
rect 15415 13345 15424 13379
rect 15372 13336 15424 13345
rect 18040 13336 18092 13388
rect 23560 13336 23612 13388
rect 13624 13268 13676 13320
rect 15740 13268 15792 13320
rect 17396 13311 17448 13320
rect 17396 13277 17405 13311
rect 17405 13277 17439 13311
rect 17439 13277 17448 13311
rect 17396 13268 17448 13277
rect 20616 13311 20668 13320
rect 20616 13277 20625 13311
rect 20625 13277 20659 13311
rect 20659 13277 20668 13311
rect 20616 13268 20668 13277
rect 14544 13200 14596 13252
rect 5360 13030 5412 13082
rect 5424 13030 5476 13082
rect 5488 13030 5540 13082
rect 5552 13030 5604 13082
rect 14694 13030 14746 13082
rect 14758 13030 14810 13082
rect 14822 13030 14874 13082
rect 14886 13030 14938 13082
rect 24027 13030 24079 13082
rect 24091 13030 24143 13082
rect 24155 13030 24207 13082
rect 24219 13030 24271 13082
rect 12796 12928 12848 12980
rect 13624 12971 13676 12980
rect 13624 12937 13633 12971
rect 13633 12937 13667 12971
rect 13667 12937 13676 12971
rect 13624 12928 13676 12937
rect 14452 12928 14504 12980
rect 15372 12928 15424 12980
rect 16200 12928 16252 12980
rect 16568 12971 16620 12980
rect 16568 12937 16577 12971
rect 16577 12937 16611 12971
rect 16611 12937 16620 12971
rect 16568 12928 16620 12937
rect 17672 12928 17724 12980
rect 18040 12928 18092 12980
rect 18316 12971 18368 12980
rect 18316 12937 18325 12971
rect 18325 12937 18359 12971
rect 18359 12937 18368 12971
rect 18316 12928 18368 12937
rect 19052 12971 19104 12980
rect 19052 12937 19061 12971
rect 19061 12937 19095 12971
rect 19095 12937 19104 12971
rect 19052 12928 19104 12937
rect 19236 12928 19288 12980
rect 14268 12860 14320 12912
rect 14176 12835 14228 12844
rect 14176 12801 14185 12835
rect 14185 12801 14219 12835
rect 14219 12801 14228 12835
rect 14176 12792 14228 12801
rect 12704 12767 12756 12776
rect 12704 12733 12713 12767
rect 12713 12733 12747 12767
rect 12747 12733 12756 12767
rect 12704 12724 12756 12733
rect 18132 12792 18184 12844
rect 19236 12835 19288 12844
rect 19236 12801 19245 12835
rect 19245 12801 19279 12835
rect 19279 12801 19288 12835
rect 19236 12792 19288 12801
rect 16384 12724 16436 12776
rect 17396 12767 17448 12776
rect 17396 12733 17405 12767
rect 17405 12733 17439 12767
rect 17439 12733 17448 12767
rect 17396 12724 17448 12733
rect 13532 12699 13584 12708
rect 13532 12665 13541 12699
rect 13541 12665 13575 12699
rect 13575 12665 13584 12699
rect 13532 12656 13584 12665
rect 15648 12656 15700 12708
rect 18868 12656 18920 12708
rect 19788 12724 19840 12776
rect 23560 12767 23612 12776
rect 23560 12733 23569 12767
rect 23569 12733 23603 12767
rect 23603 12733 23612 12767
rect 23560 12724 23612 12733
rect 12336 12631 12388 12640
rect 12336 12597 12345 12631
rect 12345 12597 12379 12631
rect 12379 12597 12388 12631
rect 12336 12588 12388 12597
rect 14084 12631 14136 12640
rect 14084 12597 14093 12631
rect 14093 12597 14127 12631
rect 14127 12597 14136 12631
rect 14084 12588 14136 12597
rect 21168 12588 21220 12640
rect 10027 12486 10079 12538
rect 10091 12486 10143 12538
rect 10155 12486 10207 12538
rect 10219 12486 10271 12538
rect 19360 12486 19412 12538
rect 19424 12486 19476 12538
rect 19488 12486 19540 12538
rect 19552 12486 19604 12538
rect 12520 12427 12572 12436
rect 12520 12393 12529 12427
rect 12529 12393 12563 12427
rect 12563 12393 12572 12427
rect 12520 12384 12572 12393
rect 14176 12384 14228 12436
rect 15372 12427 15424 12436
rect 15372 12393 15381 12427
rect 15381 12393 15415 12427
rect 15415 12393 15424 12427
rect 15372 12384 15424 12393
rect 15740 12427 15792 12436
rect 15740 12393 15749 12427
rect 15749 12393 15783 12427
rect 15783 12393 15792 12427
rect 15740 12384 15792 12393
rect 17672 12427 17724 12436
rect 17672 12393 17681 12427
rect 17681 12393 17715 12427
rect 17715 12393 17724 12427
rect 17672 12384 17724 12393
rect 15648 12316 15700 12368
rect 19144 12384 19196 12436
rect 20616 12384 20668 12436
rect 21352 12384 21404 12436
rect 22088 12316 22140 12368
rect 15740 12248 15792 12300
rect 16384 12248 16436 12300
rect 16568 12291 16620 12300
rect 16568 12257 16602 12291
rect 16602 12257 16620 12291
rect 16568 12248 16620 12257
rect 17120 12248 17172 12300
rect 18776 12248 18828 12300
rect 14544 12180 14596 12232
rect 19788 12180 19840 12232
rect 21168 12223 21220 12232
rect 21168 12189 21177 12223
rect 21177 12189 21211 12223
rect 21211 12189 21220 12223
rect 21168 12180 21220 12189
rect 21720 12112 21772 12164
rect 14084 12044 14136 12096
rect 15188 12044 15240 12096
rect 5360 11942 5412 11994
rect 5424 11942 5476 11994
rect 5488 11942 5540 11994
rect 5552 11942 5604 11994
rect 14694 11942 14746 11994
rect 14758 11942 14810 11994
rect 14822 11942 14874 11994
rect 14886 11942 14938 11994
rect 24027 11942 24079 11994
rect 24091 11942 24143 11994
rect 24155 11942 24207 11994
rect 24219 11942 24271 11994
rect 14544 11840 14596 11892
rect 15740 11883 15792 11892
rect 15740 11849 15749 11883
rect 15749 11849 15783 11883
rect 15783 11849 15792 11883
rect 15740 11840 15792 11849
rect 17120 11883 17172 11892
rect 17120 11849 17129 11883
rect 17129 11849 17163 11883
rect 17163 11849 17172 11883
rect 17120 11840 17172 11849
rect 17764 11883 17816 11892
rect 17764 11849 17773 11883
rect 17773 11849 17807 11883
rect 17807 11849 17816 11883
rect 17764 11840 17816 11849
rect 21352 11883 21404 11892
rect 21352 11849 21361 11883
rect 21361 11849 21395 11883
rect 21395 11849 21404 11883
rect 21352 11840 21404 11849
rect 22088 11883 22140 11892
rect 22088 11849 22097 11883
rect 22097 11849 22131 11883
rect 22131 11849 22140 11883
rect 22088 11840 22140 11849
rect 14360 11772 14412 11824
rect 17396 11772 17448 11824
rect 21168 11772 21220 11824
rect 14452 11704 14504 11756
rect 15648 11704 15700 11756
rect 16292 11747 16344 11756
rect 16292 11713 16301 11747
rect 16301 11713 16335 11747
rect 16335 11713 16344 11747
rect 18316 11747 18368 11756
rect 16292 11704 16344 11713
rect 18316 11713 18325 11747
rect 18325 11713 18359 11747
rect 18359 11713 18368 11747
rect 18316 11704 18368 11713
rect 19052 11636 19104 11688
rect 19236 11636 19288 11688
rect 14544 11543 14596 11552
rect 14544 11509 14553 11543
rect 14553 11509 14587 11543
rect 14587 11509 14596 11543
rect 14544 11500 14596 11509
rect 15188 11543 15240 11552
rect 15188 11509 15197 11543
rect 15197 11509 15231 11543
rect 15231 11509 15240 11543
rect 15188 11500 15240 11509
rect 17488 11543 17540 11552
rect 17488 11509 17497 11543
rect 17497 11509 17531 11543
rect 17531 11509 17540 11543
rect 17488 11500 17540 11509
rect 18776 11500 18828 11552
rect 24480 11636 24532 11688
rect 19788 11568 19840 11620
rect 20248 11500 20300 11552
rect 20432 11500 20484 11552
rect 24480 11543 24532 11552
rect 24480 11509 24489 11543
rect 24489 11509 24523 11543
rect 24523 11509 24532 11543
rect 24480 11500 24532 11509
rect 10027 11398 10079 11450
rect 10091 11398 10143 11450
rect 10155 11398 10207 11450
rect 10219 11398 10271 11450
rect 19360 11398 19412 11450
rect 19424 11398 19476 11450
rect 19488 11398 19540 11450
rect 19552 11398 19604 11450
rect 18316 11296 18368 11348
rect 18868 11339 18920 11348
rect 18868 11305 18877 11339
rect 18877 11305 18911 11339
rect 18911 11305 18920 11339
rect 18868 11296 18920 11305
rect 19052 11296 19104 11348
rect 19788 11339 19840 11348
rect 19788 11305 19797 11339
rect 19797 11305 19831 11339
rect 19831 11305 19840 11339
rect 19788 11296 19840 11305
rect 15188 11228 15240 11280
rect 21168 11228 21220 11280
rect 20248 11092 20300 11144
rect 19788 11024 19840 11076
rect 19236 10956 19288 11008
rect 22364 10956 22416 11008
rect 5360 10854 5412 10906
rect 5424 10854 5476 10906
rect 5488 10854 5540 10906
rect 5552 10854 5604 10906
rect 14694 10854 14746 10906
rect 14758 10854 14810 10906
rect 14822 10854 14874 10906
rect 14886 10854 14938 10906
rect 24027 10854 24079 10906
rect 24091 10854 24143 10906
rect 24155 10854 24207 10906
rect 24219 10854 24271 10906
rect 18684 10548 18736 10600
rect 15280 10523 15332 10532
rect 15280 10489 15289 10523
rect 15289 10489 15323 10523
rect 15323 10489 15332 10523
rect 15280 10480 15332 10489
rect 18040 10480 18092 10532
rect 19696 10548 19748 10600
rect 20340 10548 20392 10600
rect 20984 10548 21036 10600
rect 22364 10616 22416 10668
rect 23100 10548 23152 10600
rect 14544 10412 14596 10464
rect 18684 10412 18736 10464
rect 20432 10455 20484 10464
rect 20432 10421 20441 10455
rect 20441 10421 20475 10455
rect 20475 10421 20484 10455
rect 20432 10412 20484 10421
rect 21536 10455 21588 10464
rect 21536 10421 21545 10455
rect 21545 10421 21579 10455
rect 21579 10421 21588 10455
rect 21536 10412 21588 10421
rect 10027 10310 10079 10362
rect 10091 10310 10143 10362
rect 10155 10310 10207 10362
rect 10219 10310 10271 10362
rect 19360 10310 19412 10362
rect 19424 10310 19476 10362
rect 19488 10310 19540 10362
rect 19552 10310 19604 10362
rect 21076 10251 21128 10260
rect 21076 10217 21085 10251
rect 21085 10217 21119 10251
rect 21119 10217 21128 10251
rect 21076 10208 21128 10217
rect 22364 10208 22416 10260
rect 21536 10140 21588 10192
rect 19236 10115 19288 10124
rect 19236 10081 19245 10115
rect 19245 10081 19279 10115
rect 19279 10081 19288 10115
rect 19236 10072 19288 10081
rect 20984 10115 21036 10124
rect 20984 10081 20993 10115
rect 20993 10081 21027 10115
rect 21027 10081 21036 10115
rect 20984 10072 21036 10081
rect 19696 10004 19748 10056
rect 20432 10004 20484 10056
rect 19052 9936 19104 9988
rect 18868 9911 18920 9920
rect 18868 9877 18877 9911
rect 18877 9877 18911 9911
rect 18911 9877 18920 9911
rect 18868 9868 18920 9877
rect 20340 9911 20392 9920
rect 20340 9877 20349 9911
rect 20349 9877 20383 9911
rect 20383 9877 20392 9911
rect 20340 9868 20392 9877
rect 20616 9911 20668 9920
rect 20616 9877 20625 9911
rect 20625 9877 20659 9911
rect 20659 9877 20668 9911
rect 20616 9868 20668 9877
rect 5360 9766 5412 9818
rect 5424 9766 5476 9818
rect 5488 9766 5540 9818
rect 5552 9766 5604 9818
rect 14694 9766 14746 9818
rect 14758 9766 14810 9818
rect 14822 9766 14874 9818
rect 14886 9766 14938 9818
rect 24027 9766 24079 9818
rect 24091 9766 24143 9818
rect 24155 9766 24207 9818
rect 24219 9766 24271 9818
rect 18040 9707 18092 9716
rect 18040 9673 18049 9707
rect 18049 9673 18083 9707
rect 18083 9673 18092 9707
rect 18040 9664 18092 9673
rect 19236 9664 19288 9716
rect 21076 9664 21128 9716
rect 21996 9664 22048 9716
rect 22272 9664 22324 9716
rect 14912 9571 14964 9580
rect 14912 9537 14921 9571
rect 14921 9537 14955 9571
rect 14955 9537 14964 9571
rect 14912 9528 14964 9537
rect 18684 9460 18736 9512
rect 20340 9460 20392 9512
rect 19052 9392 19104 9444
rect 20432 9392 20484 9444
rect 14452 9324 14504 9376
rect 18868 9324 18920 9376
rect 20248 9367 20300 9376
rect 20248 9333 20257 9367
rect 20257 9333 20291 9367
rect 20291 9333 20300 9367
rect 20248 9324 20300 9333
rect 20984 9324 21036 9376
rect 21352 9324 21404 9376
rect 10027 9222 10079 9274
rect 10091 9222 10143 9274
rect 10155 9222 10207 9274
rect 10219 9222 10271 9274
rect 19360 9222 19412 9274
rect 19424 9222 19476 9274
rect 19488 9222 19540 9274
rect 19552 9222 19604 9274
rect 18960 9120 19012 9172
rect 16016 8984 16068 9036
rect 18684 8984 18736 9036
rect 19420 8916 19472 8968
rect 20248 9120 20300 9172
rect 20432 9120 20484 9172
rect 16200 8780 16252 8832
rect 17580 8780 17632 8832
rect 5360 8678 5412 8730
rect 5424 8678 5476 8730
rect 5488 8678 5540 8730
rect 5552 8678 5604 8730
rect 14694 8678 14746 8730
rect 14758 8678 14810 8730
rect 14822 8678 14874 8730
rect 14886 8678 14938 8730
rect 24027 8678 24079 8730
rect 24091 8678 24143 8730
rect 24155 8678 24207 8730
rect 24219 8678 24271 8730
rect 14452 8619 14504 8628
rect 14452 8585 14461 8619
rect 14461 8585 14495 8619
rect 14495 8585 14504 8619
rect 14452 8576 14504 8585
rect 18684 8619 18736 8628
rect 18684 8585 18693 8619
rect 18693 8585 18727 8619
rect 18727 8585 18736 8619
rect 18684 8576 18736 8585
rect 14268 8508 14320 8560
rect 16016 8551 16068 8560
rect 16016 8517 16025 8551
rect 16025 8517 16059 8551
rect 16059 8517 16068 8551
rect 16016 8508 16068 8517
rect 18868 8372 18920 8424
rect 19052 8372 19104 8424
rect 19420 8415 19472 8424
rect 19420 8381 19454 8415
rect 19454 8381 19472 8415
rect 19420 8372 19472 8381
rect 19052 8279 19104 8288
rect 19052 8245 19061 8279
rect 19061 8245 19095 8279
rect 19095 8245 19104 8279
rect 19052 8236 19104 8245
rect 21260 8236 21312 8288
rect 10027 8134 10079 8186
rect 10091 8134 10143 8186
rect 10155 8134 10207 8186
rect 10219 8134 10271 8186
rect 19360 8134 19412 8186
rect 19424 8134 19476 8186
rect 19488 8134 19540 8186
rect 19552 8134 19604 8186
rect 18960 8032 19012 8084
rect 16752 7896 16804 7948
rect 17580 7896 17632 7948
rect 21352 7896 21404 7948
rect 19236 7871 19288 7880
rect 19236 7837 19245 7871
rect 19245 7837 19279 7871
rect 19279 7837 19288 7871
rect 19236 7828 19288 7837
rect 21076 7871 21128 7880
rect 21076 7837 21085 7871
rect 21085 7837 21119 7871
rect 21119 7837 21128 7871
rect 21076 7828 21128 7837
rect 21260 7871 21312 7880
rect 21260 7837 21269 7871
rect 21269 7837 21303 7871
rect 21303 7837 21312 7871
rect 21260 7828 21312 7837
rect 16384 7692 16436 7744
rect 20616 7735 20668 7744
rect 20616 7701 20625 7735
rect 20625 7701 20659 7735
rect 20659 7701 20668 7735
rect 20616 7692 20668 7701
rect 5360 7590 5412 7642
rect 5424 7590 5476 7642
rect 5488 7590 5540 7642
rect 5552 7590 5604 7642
rect 14694 7590 14746 7642
rect 14758 7590 14810 7642
rect 14822 7590 14874 7642
rect 14886 7590 14938 7642
rect 24027 7590 24079 7642
rect 24091 7590 24143 7642
rect 24155 7590 24207 7642
rect 24219 7590 24271 7642
rect 16384 7531 16436 7540
rect 16384 7497 16393 7531
rect 16393 7497 16427 7531
rect 16427 7497 16436 7531
rect 16384 7488 16436 7497
rect 16752 7531 16804 7540
rect 16752 7497 16761 7531
rect 16761 7497 16795 7531
rect 16795 7497 16804 7531
rect 16752 7488 16804 7497
rect 18408 7531 18460 7540
rect 18408 7497 18417 7531
rect 18417 7497 18451 7531
rect 18451 7497 18460 7531
rect 18408 7488 18460 7497
rect 21076 7488 21128 7540
rect 23100 7488 23152 7540
rect 21260 7420 21312 7472
rect 16384 7284 16436 7336
rect 18408 7284 18460 7336
rect 19052 7284 19104 7336
rect 15648 7148 15700 7200
rect 17672 7148 17724 7200
rect 19972 7148 20024 7200
rect 20432 7148 20484 7200
rect 21352 7148 21404 7200
rect 10027 7046 10079 7098
rect 10091 7046 10143 7098
rect 10155 7046 10207 7098
rect 10219 7046 10271 7098
rect 19360 7046 19412 7098
rect 19424 7046 19476 7098
rect 19488 7046 19540 7098
rect 19552 7046 19604 7098
rect 19236 6944 19288 6996
rect 22272 6987 22324 6996
rect 22272 6953 22281 6987
rect 22281 6953 22315 6987
rect 22315 6953 22324 6987
rect 22272 6944 22324 6953
rect 17856 6851 17908 6860
rect 17856 6817 17865 6851
rect 17865 6817 17899 6851
rect 17899 6817 17908 6851
rect 17856 6808 17908 6817
rect 20616 6876 20668 6928
rect 19144 6740 19196 6792
rect 21536 6808 21588 6860
rect 19052 6672 19104 6724
rect 19972 6740 20024 6792
rect 20432 6672 20484 6724
rect 18408 6604 18460 6656
rect 18500 6604 18552 6656
rect 5360 6502 5412 6554
rect 5424 6502 5476 6554
rect 5488 6502 5540 6554
rect 5552 6502 5604 6554
rect 14694 6502 14746 6554
rect 14758 6502 14810 6554
rect 14822 6502 14874 6554
rect 14886 6502 14938 6554
rect 24027 6502 24079 6554
rect 24091 6502 24143 6554
rect 24155 6502 24207 6554
rect 24219 6502 24271 6554
rect 17856 6400 17908 6452
rect 19144 6400 19196 6452
rect 19236 6400 19288 6452
rect 19972 6443 20024 6452
rect 19972 6409 19981 6443
rect 19981 6409 20015 6443
rect 20015 6409 20024 6443
rect 19972 6400 20024 6409
rect 19236 6307 19288 6316
rect 19236 6273 19245 6307
rect 19245 6273 19279 6307
rect 19279 6273 19288 6307
rect 19236 6264 19288 6273
rect 20432 6239 20484 6248
rect 20432 6205 20466 6239
rect 20466 6205 20484 6239
rect 20432 6196 20484 6205
rect 18960 6060 19012 6112
rect 21536 6103 21588 6112
rect 21536 6069 21545 6103
rect 21545 6069 21579 6103
rect 21579 6069 21588 6103
rect 22180 6103 22232 6112
rect 21536 6060 21588 6069
rect 22180 6069 22189 6103
rect 22189 6069 22223 6103
rect 22223 6069 22232 6103
rect 22180 6060 22232 6069
rect 10027 5958 10079 6010
rect 10091 5958 10143 6010
rect 10155 5958 10207 6010
rect 10219 5958 10271 6010
rect 19360 5958 19412 6010
rect 19424 5958 19476 6010
rect 19488 5958 19540 6010
rect 19552 5958 19604 6010
rect 19052 5899 19104 5908
rect 19052 5865 19061 5899
rect 19061 5865 19095 5899
rect 19095 5865 19104 5899
rect 19052 5856 19104 5865
rect 19972 5856 20024 5908
rect 16936 5763 16988 5772
rect 16936 5729 16945 5763
rect 16945 5729 16979 5763
rect 16979 5729 16988 5763
rect 16936 5720 16988 5729
rect 18132 5720 18184 5772
rect 18500 5720 18552 5772
rect 19696 5720 19748 5772
rect 20984 5720 21036 5772
rect 21352 5763 21404 5772
rect 21352 5729 21361 5763
rect 21361 5729 21395 5763
rect 21395 5729 21404 5763
rect 21352 5720 21404 5729
rect 21444 5695 21496 5704
rect 21444 5661 21453 5695
rect 21453 5661 21487 5695
rect 21487 5661 21496 5695
rect 21444 5652 21496 5661
rect 22180 5652 22232 5704
rect 17028 5516 17080 5568
rect 19788 5516 19840 5568
rect 21720 5516 21772 5568
rect 5360 5414 5412 5466
rect 5424 5414 5476 5466
rect 5488 5414 5540 5466
rect 5552 5414 5604 5466
rect 14694 5414 14746 5466
rect 14758 5414 14810 5466
rect 14822 5414 14874 5466
rect 14886 5414 14938 5466
rect 24027 5414 24079 5466
rect 24091 5414 24143 5466
rect 24155 5414 24207 5466
rect 24219 5414 24271 5466
rect 16936 5355 16988 5364
rect 16936 5321 16945 5355
rect 16945 5321 16979 5355
rect 16979 5321 16988 5355
rect 16936 5312 16988 5321
rect 18132 5355 18184 5364
rect 18132 5321 18141 5355
rect 18141 5321 18175 5355
rect 18175 5321 18184 5355
rect 18132 5312 18184 5321
rect 19696 5312 19748 5364
rect 22180 5312 22232 5364
rect 21720 5219 21772 5228
rect 21720 5185 21729 5219
rect 21729 5185 21763 5219
rect 21763 5185 21772 5219
rect 21720 5176 21772 5185
rect 21812 5176 21864 5228
rect 22272 5176 22324 5228
rect 21628 5083 21680 5092
rect 21628 5049 21637 5083
rect 21637 5049 21671 5083
rect 21671 5049 21680 5083
rect 21628 5040 21680 5049
rect 20156 5015 20208 5024
rect 20156 4981 20165 5015
rect 20165 4981 20199 5015
rect 20199 4981 20208 5015
rect 20156 4972 20208 4981
rect 20984 5015 21036 5024
rect 20984 4981 20993 5015
rect 20993 4981 21027 5015
rect 21027 4981 21036 5015
rect 20984 4972 21036 4981
rect 21260 5015 21312 5024
rect 21260 4981 21269 5015
rect 21269 4981 21303 5015
rect 21303 4981 21312 5015
rect 21260 4972 21312 4981
rect 10027 4870 10079 4922
rect 10091 4870 10143 4922
rect 10155 4870 10207 4922
rect 10219 4870 10271 4922
rect 19360 4870 19412 4922
rect 19424 4870 19476 4922
rect 19488 4870 19540 4922
rect 19552 4870 19604 4922
rect 21628 4811 21680 4820
rect 21628 4777 21637 4811
rect 21637 4777 21671 4811
rect 21671 4777 21680 4811
rect 21628 4768 21680 4777
rect 21720 4768 21772 4820
rect 21812 4700 21864 4752
rect 20616 4632 20668 4684
rect 21260 4632 21312 4684
rect 24296 4675 24348 4684
rect 24296 4641 24305 4675
rect 24305 4641 24339 4675
rect 24339 4641 24348 4675
rect 24296 4632 24348 4641
rect 21812 4496 21864 4548
rect 23192 4428 23244 4480
rect 5360 4326 5412 4378
rect 5424 4326 5476 4378
rect 5488 4326 5540 4378
rect 5552 4326 5604 4378
rect 14694 4326 14746 4378
rect 14758 4326 14810 4378
rect 14822 4326 14874 4378
rect 14886 4326 14938 4378
rect 24027 4326 24079 4378
rect 24091 4326 24143 4378
rect 24155 4326 24207 4378
rect 24219 4326 24271 4378
rect 20616 4267 20668 4276
rect 20616 4233 20625 4267
rect 20625 4233 20659 4267
rect 20659 4233 20668 4267
rect 20616 4224 20668 4233
rect 24388 4224 24440 4276
rect 21536 4088 21588 4140
rect 21812 4063 21864 4072
rect 21812 4029 21821 4063
rect 21821 4029 21855 4063
rect 21855 4029 21864 4063
rect 21812 4020 21864 4029
rect 23928 4020 23980 4072
rect 21076 3884 21128 3936
rect 22456 3952 22508 4004
rect 24480 3927 24532 3936
rect 24480 3893 24489 3927
rect 24489 3893 24523 3927
rect 24523 3893 24532 3927
rect 24480 3884 24532 3893
rect 10027 3782 10079 3834
rect 10091 3782 10143 3834
rect 10155 3782 10207 3834
rect 10219 3782 10271 3834
rect 19360 3782 19412 3834
rect 19424 3782 19476 3834
rect 19488 3782 19540 3834
rect 19552 3782 19604 3834
rect 24388 3544 24440 3596
rect 8012 3476 8064 3528
rect 8840 3476 8892 3528
rect 10772 3476 10824 3528
rect 11600 3476 11652 3528
rect 12244 3476 12296 3528
rect 12704 3476 12756 3528
rect 12888 3476 12940 3528
rect 13440 3476 13492 3528
rect 23652 3383 23704 3392
rect 23652 3349 23661 3383
rect 23661 3349 23695 3383
rect 23695 3349 23704 3383
rect 23652 3340 23704 3349
rect 25216 3340 25268 3392
rect 5360 3238 5412 3290
rect 5424 3238 5476 3290
rect 5488 3238 5540 3290
rect 5552 3238 5604 3290
rect 14694 3238 14746 3290
rect 14758 3238 14810 3290
rect 14822 3238 14874 3290
rect 14886 3238 14938 3290
rect 24027 3238 24079 3290
rect 24091 3238 24143 3290
rect 24155 3238 24207 3290
rect 24219 3238 24271 3290
rect 21812 3136 21864 3188
rect 23100 3136 23152 3188
rect 24388 3179 24440 3188
rect 24388 3145 24397 3179
rect 24397 3145 24431 3179
rect 24431 3145 24440 3179
rect 24388 3136 24440 3145
rect 23652 2975 23704 2984
rect 23652 2941 23661 2975
rect 23661 2941 23695 2975
rect 23695 2941 23704 2975
rect 23652 2932 23704 2941
rect 23836 2839 23888 2848
rect 23836 2805 23845 2839
rect 23845 2805 23879 2839
rect 23879 2805 23888 2839
rect 23836 2796 23888 2805
rect 24480 2796 24532 2848
rect 25308 2839 25360 2848
rect 25308 2805 25317 2839
rect 25317 2805 25351 2839
rect 25351 2805 25360 2839
rect 25308 2796 25360 2805
rect 10027 2694 10079 2746
rect 10091 2694 10143 2746
rect 10155 2694 10207 2746
rect 10219 2694 10271 2746
rect 19360 2694 19412 2746
rect 19424 2694 19476 2746
rect 19488 2694 19540 2746
rect 19552 2694 19604 2746
rect 21628 2592 21680 2644
rect 22732 2635 22784 2644
rect 22732 2601 22741 2635
rect 22741 2601 22775 2635
rect 22775 2601 22784 2635
rect 22732 2592 22784 2601
rect 24388 2592 24440 2644
rect 23284 2388 23336 2440
rect 20432 2252 20484 2304
rect 23192 2252 23244 2304
rect 5360 2150 5412 2202
rect 5424 2150 5476 2202
rect 5488 2150 5540 2202
rect 5552 2150 5604 2202
rect 14694 2150 14746 2202
rect 14758 2150 14810 2202
rect 14822 2150 14874 2202
rect 14886 2150 14938 2202
rect 24027 2150 24079 2202
rect 24091 2150 24143 2202
rect 24155 2150 24207 2202
rect 24219 2150 24271 2202
rect 7276 552 7328 604
rect 7460 552 7512 604
rect 8104 552 8156 604
rect 8472 552 8524 604
rect 13624 552 13676 604
rect 13808 552 13860 604
<< metal2 >>
rect 4330 27520 4386 28000
rect 13622 27520 13678 28000
rect 22914 27520 22970 28000
rect 23834 27568 23890 27577
rect 1848 23180 1900 23186
rect 1848 23122 1900 23128
rect 1860 22438 1888 23122
rect 2030 23080 2086 23089
rect 2030 23015 2032 23024
rect 2084 23015 2086 23024
rect 2032 22986 2084 22992
rect 2492 22568 2544 22574
rect 2492 22510 2544 22516
rect 2674 22536 2730 22545
rect 1848 22432 1900 22438
rect 1848 22374 1900 22380
rect 650 4040 706 4049
rect 650 3975 706 3984
rect 6 3496 62 3505
rect 6 3431 62 3440
rect 20 480 48 3431
rect 664 480 692 3975
rect 1860 3346 1888 22374
rect 2504 3346 2532 22510
rect 2674 22471 2730 22480
rect 2688 22438 2716 22471
rect 2676 22432 2728 22438
rect 2676 22374 2728 22380
rect 4054 22400 4110 22409
rect 4054 22335 4110 22344
rect 3780 22092 3832 22098
rect 3780 22034 3832 22040
rect 3792 21554 3820 22034
rect 3962 21992 4018 22001
rect 3962 21927 3964 21936
rect 4016 21927 4018 21936
rect 3964 21898 4016 21904
rect 4068 21690 4096 22335
rect 4056 21684 4108 21690
rect 4056 21626 4108 21632
rect 3780 21548 3832 21554
rect 3780 21490 3832 21496
rect 3792 3482 3820 21490
rect 3872 21344 3924 21350
rect 3872 21286 3924 21292
rect 3424 3454 3820 3482
rect 1860 3318 2072 3346
rect 2504 3318 2716 3346
rect 1294 3088 1350 3097
rect 1294 3023 1350 3032
rect 1308 480 1336 3023
rect 2044 480 2072 3318
rect 2688 480 2716 3318
rect 3424 480 3452 3454
rect 3884 3346 3912 21286
rect 4344 13841 4372 27520
rect 10001 25596 10297 25616
rect 10057 25594 10081 25596
rect 10137 25594 10161 25596
rect 10217 25594 10241 25596
rect 10079 25542 10081 25594
rect 10143 25542 10155 25594
rect 10217 25542 10219 25594
rect 10057 25540 10081 25542
rect 10137 25540 10161 25542
rect 10217 25540 10241 25542
rect 10001 25520 10297 25540
rect 5334 25052 5630 25072
rect 5390 25050 5414 25052
rect 5470 25050 5494 25052
rect 5550 25050 5574 25052
rect 5412 24998 5414 25050
rect 5476 24998 5488 25050
rect 5550 24998 5552 25050
rect 5390 24996 5414 24998
rect 5470 24996 5494 24998
rect 5550 24996 5574 24998
rect 5334 24976 5630 24996
rect 11232 24948 11284 24954
rect 11232 24890 11284 24896
rect 10680 24880 10732 24886
rect 10680 24822 10732 24828
rect 10001 24508 10297 24528
rect 10057 24506 10081 24508
rect 10137 24506 10161 24508
rect 10217 24506 10241 24508
rect 10079 24454 10081 24506
rect 10143 24454 10155 24506
rect 10217 24454 10219 24506
rect 10057 24452 10081 24454
rect 10137 24452 10161 24454
rect 10217 24452 10241 24454
rect 10001 24432 10297 24452
rect 5334 23964 5630 23984
rect 5390 23962 5414 23964
rect 5470 23962 5494 23964
rect 5550 23962 5574 23964
rect 5412 23910 5414 23962
rect 5476 23910 5488 23962
rect 5550 23910 5552 23962
rect 5390 23908 5414 23910
rect 5470 23908 5494 23910
rect 5550 23908 5574 23910
rect 5334 23888 5630 23908
rect 10001 23420 10297 23440
rect 10057 23418 10081 23420
rect 10137 23418 10161 23420
rect 10217 23418 10241 23420
rect 10079 23366 10081 23418
rect 10143 23366 10155 23418
rect 10217 23366 10219 23418
rect 10057 23364 10081 23366
rect 10137 23364 10161 23366
rect 10217 23364 10241 23366
rect 10001 23344 10297 23364
rect 5710 22944 5766 22953
rect 5334 22876 5630 22896
rect 5710 22879 5766 22888
rect 5390 22874 5414 22876
rect 5470 22874 5494 22876
rect 5550 22874 5574 22876
rect 5412 22822 5414 22874
rect 5476 22822 5488 22874
rect 5550 22822 5552 22874
rect 5390 22820 5414 22822
rect 5470 22820 5494 22822
rect 5550 22820 5574 22822
rect 5334 22800 5630 22820
rect 5724 22409 5752 22879
rect 5710 22400 5766 22409
rect 5710 22335 5766 22344
rect 10001 22332 10297 22352
rect 10057 22330 10081 22332
rect 10137 22330 10161 22332
rect 10217 22330 10241 22332
rect 10079 22278 10081 22330
rect 10143 22278 10155 22330
rect 10217 22278 10219 22330
rect 10057 22276 10081 22278
rect 10137 22276 10161 22278
rect 10217 22276 10241 22278
rect 10001 22256 10297 22276
rect 5334 21788 5630 21808
rect 5390 21786 5414 21788
rect 5470 21786 5494 21788
rect 5550 21786 5574 21788
rect 5412 21734 5414 21786
rect 5476 21734 5488 21786
rect 5550 21734 5552 21786
rect 5390 21732 5414 21734
rect 5470 21732 5494 21734
rect 5550 21732 5574 21734
rect 5334 21712 5630 21732
rect 10001 21244 10297 21264
rect 10057 21242 10081 21244
rect 10137 21242 10161 21244
rect 10217 21242 10241 21244
rect 10079 21190 10081 21242
rect 10143 21190 10155 21242
rect 10217 21190 10219 21242
rect 10057 21188 10081 21190
rect 10137 21188 10161 21190
rect 10217 21188 10241 21190
rect 10001 21168 10297 21188
rect 5710 20904 5766 20913
rect 5710 20839 5766 20848
rect 5334 20700 5630 20720
rect 5390 20698 5414 20700
rect 5470 20698 5494 20700
rect 5550 20698 5574 20700
rect 5412 20646 5414 20698
rect 5476 20646 5488 20698
rect 5550 20646 5552 20698
rect 5390 20644 5414 20646
rect 5470 20644 5494 20646
rect 5550 20644 5574 20646
rect 5334 20624 5630 20644
rect 5724 20058 5752 20839
rect 10001 20156 10297 20176
rect 10057 20154 10081 20156
rect 10137 20154 10161 20156
rect 10217 20154 10241 20156
rect 10079 20102 10081 20154
rect 10143 20102 10155 20154
rect 10217 20102 10219 20154
rect 10057 20100 10081 20102
rect 10137 20100 10161 20102
rect 10217 20100 10241 20102
rect 10001 20080 10297 20100
rect 5712 20052 5764 20058
rect 5712 19994 5764 20000
rect 6722 19952 6778 19961
rect 5252 19916 5304 19922
rect 6722 19887 6778 19896
rect 5252 19858 5304 19864
rect 5264 19174 5292 19858
rect 5334 19612 5630 19632
rect 5390 19610 5414 19612
rect 5470 19610 5494 19612
rect 5550 19610 5574 19612
rect 5412 19558 5414 19610
rect 5476 19558 5488 19610
rect 5550 19558 5552 19610
rect 5390 19556 5414 19558
rect 5470 19556 5494 19558
rect 5550 19556 5574 19558
rect 5334 19536 5630 19556
rect 6540 19304 6592 19310
rect 6540 19246 6592 19252
rect 5252 19168 5304 19174
rect 5252 19110 5304 19116
rect 4330 13832 4386 13841
rect 4330 13767 4386 13776
rect 4698 3632 4754 3641
rect 4698 3567 4754 3576
rect 3884 3318 4096 3346
rect 4068 480 4096 3318
rect 4712 480 4740 3567
rect 5264 1986 5292 19110
rect 5334 18524 5630 18544
rect 5390 18522 5414 18524
rect 5470 18522 5494 18524
rect 5550 18522 5574 18524
rect 5412 18470 5414 18522
rect 5476 18470 5488 18522
rect 5550 18470 5552 18522
rect 5390 18468 5414 18470
rect 5470 18468 5494 18470
rect 5550 18468 5574 18470
rect 5334 18448 5630 18468
rect 5334 17436 5630 17456
rect 5390 17434 5414 17436
rect 5470 17434 5494 17436
rect 5550 17434 5574 17436
rect 5412 17382 5414 17434
rect 5476 17382 5488 17434
rect 5550 17382 5552 17434
rect 5390 17380 5414 17382
rect 5470 17380 5494 17382
rect 5550 17380 5574 17382
rect 5334 17360 5630 17380
rect 5334 16348 5630 16368
rect 5390 16346 5414 16348
rect 5470 16346 5494 16348
rect 5550 16346 5574 16348
rect 5412 16294 5414 16346
rect 5476 16294 5488 16346
rect 5550 16294 5552 16346
rect 5390 16292 5414 16294
rect 5470 16292 5494 16294
rect 5550 16292 5574 16294
rect 5334 16272 5630 16292
rect 5334 15260 5630 15280
rect 5390 15258 5414 15260
rect 5470 15258 5494 15260
rect 5550 15258 5574 15260
rect 5412 15206 5414 15258
rect 5476 15206 5488 15258
rect 5550 15206 5552 15258
rect 5390 15204 5414 15206
rect 5470 15204 5494 15206
rect 5550 15204 5574 15206
rect 5334 15184 5630 15204
rect 5334 14172 5630 14192
rect 5390 14170 5414 14172
rect 5470 14170 5494 14172
rect 5550 14170 5574 14172
rect 5412 14118 5414 14170
rect 5476 14118 5488 14170
rect 5550 14118 5552 14170
rect 5390 14116 5414 14118
rect 5470 14116 5494 14118
rect 5550 14116 5574 14118
rect 5334 14096 5630 14116
rect 5334 13084 5630 13104
rect 5390 13082 5414 13084
rect 5470 13082 5494 13084
rect 5550 13082 5574 13084
rect 5412 13030 5414 13082
rect 5476 13030 5488 13082
rect 5550 13030 5552 13082
rect 5390 13028 5414 13030
rect 5470 13028 5494 13030
rect 5550 13028 5574 13030
rect 5334 13008 5630 13028
rect 5334 11996 5630 12016
rect 5390 11994 5414 11996
rect 5470 11994 5494 11996
rect 5550 11994 5574 11996
rect 5412 11942 5414 11994
rect 5476 11942 5488 11994
rect 5550 11942 5552 11994
rect 5390 11940 5414 11942
rect 5470 11940 5494 11942
rect 5550 11940 5574 11942
rect 5334 11920 5630 11940
rect 5334 10908 5630 10928
rect 5390 10906 5414 10908
rect 5470 10906 5494 10908
rect 5550 10906 5574 10908
rect 5412 10854 5414 10906
rect 5476 10854 5488 10906
rect 5550 10854 5552 10906
rect 5390 10852 5414 10854
rect 5470 10852 5494 10854
rect 5550 10852 5574 10854
rect 5334 10832 5630 10852
rect 5334 9820 5630 9840
rect 5390 9818 5414 9820
rect 5470 9818 5494 9820
rect 5550 9818 5574 9820
rect 5412 9766 5414 9818
rect 5476 9766 5488 9818
rect 5550 9766 5552 9818
rect 5390 9764 5414 9766
rect 5470 9764 5494 9766
rect 5550 9764 5574 9766
rect 5334 9744 5630 9764
rect 5334 8732 5630 8752
rect 5390 8730 5414 8732
rect 5470 8730 5494 8732
rect 5550 8730 5574 8732
rect 5412 8678 5414 8730
rect 5476 8678 5488 8730
rect 5550 8678 5552 8730
rect 5390 8676 5414 8678
rect 5470 8676 5494 8678
rect 5550 8676 5574 8678
rect 5334 8656 5630 8676
rect 5334 7644 5630 7664
rect 5390 7642 5414 7644
rect 5470 7642 5494 7644
rect 5550 7642 5574 7644
rect 5412 7590 5414 7642
rect 5476 7590 5488 7642
rect 5550 7590 5552 7642
rect 5390 7588 5414 7590
rect 5470 7588 5494 7590
rect 5550 7588 5574 7590
rect 5334 7568 5630 7588
rect 5334 6556 5630 6576
rect 5390 6554 5414 6556
rect 5470 6554 5494 6556
rect 5550 6554 5574 6556
rect 5412 6502 5414 6554
rect 5476 6502 5488 6554
rect 5550 6502 5552 6554
rect 5390 6500 5414 6502
rect 5470 6500 5494 6502
rect 5550 6500 5574 6502
rect 5334 6480 5630 6500
rect 5334 5468 5630 5488
rect 5390 5466 5414 5468
rect 5470 5466 5494 5468
rect 5550 5466 5574 5468
rect 5412 5414 5414 5466
rect 5476 5414 5488 5466
rect 5550 5414 5552 5466
rect 5390 5412 5414 5414
rect 5470 5412 5494 5414
rect 5550 5412 5574 5414
rect 5334 5392 5630 5412
rect 5334 4380 5630 4400
rect 5390 4378 5414 4380
rect 5470 4378 5494 4380
rect 5550 4378 5574 4380
rect 5412 4326 5414 4378
rect 5476 4326 5488 4378
rect 5550 4326 5552 4378
rect 5390 4324 5414 4326
rect 5470 4324 5494 4326
rect 5550 4324 5574 4326
rect 5334 4304 5630 4324
rect 6552 3482 6580 19246
rect 6736 19174 6764 19887
rect 6814 19408 6870 19417
rect 6814 19343 6870 19352
rect 6724 19168 6776 19174
rect 6724 19110 6776 19116
rect 6828 18970 6856 19343
rect 10001 19068 10297 19088
rect 10057 19066 10081 19068
rect 10137 19066 10161 19068
rect 10217 19066 10241 19068
rect 10079 19014 10081 19066
rect 10143 19014 10155 19066
rect 10217 19014 10219 19066
rect 10057 19012 10081 19014
rect 10137 19012 10161 19014
rect 10217 19012 10241 19014
rect 10001 18992 10297 19012
rect 6816 18964 6868 18970
rect 6816 18906 6868 18912
rect 6724 18828 6776 18834
rect 6724 18770 6776 18776
rect 6736 18086 6764 18770
rect 6724 18080 6776 18086
rect 6724 18022 6776 18028
rect 6092 3454 6580 3482
rect 5334 3292 5630 3312
rect 5390 3290 5414 3292
rect 5470 3290 5494 3292
rect 5550 3290 5574 3292
rect 5412 3238 5414 3290
rect 5476 3238 5488 3290
rect 5550 3238 5552 3290
rect 5390 3236 5414 3238
rect 5470 3236 5494 3238
rect 5550 3236 5574 3238
rect 5334 3216 5630 3236
rect 5334 2204 5630 2224
rect 5390 2202 5414 2204
rect 5470 2202 5494 2204
rect 5550 2202 5574 2204
rect 5412 2150 5414 2202
rect 5476 2150 5488 2202
rect 5550 2150 5552 2202
rect 5390 2148 5414 2150
rect 5470 2148 5494 2150
rect 5550 2148 5574 2150
rect 5334 2128 5630 2148
rect 5264 1958 5476 1986
rect 5448 480 5476 1958
rect 6092 480 6120 3454
rect 6736 626 6764 18022
rect 10001 17980 10297 18000
rect 10057 17978 10081 17980
rect 10137 17978 10161 17980
rect 10217 17978 10241 17980
rect 10079 17926 10081 17978
rect 10143 17926 10155 17978
rect 10217 17926 10219 17978
rect 10057 17924 10081 17926
rect 10137 17924 10161 17926
rect 10217 17924 10241 17926
rect 10001 17904 10297 17924
rect 10692 17882 10720 24822
rect 10680 17876 10732 17882
rect 10680 17818 10732 17824
rect 7276 17740 7328 17746
rect 7276 17682 7328 17688
rect 10496 17740 10548 17746
rect 10496 17682 10548 17688
rect 7288 16998 7316 17682
rect 7458 17640 7514 17649
rect 7458 17575 7460 17584
rect 7512 17575 7514 17584
rect 7460 17546 7512 17552
rect 9574 17232 9630 17241
rect 9574 17167 9630 17176
rect 8102 17096 8158 17105
rect 8102 17031 8158 17040
rect 8116 16998 8144 17031
rect 7276 16992 7328 16998
rect 7276 16934 7328 16940
rect 8104 16992 8156 16998
rect 8104 16934 8156 16940
rect 8472 16992 8524 16998
rect 8472 16934 8524 16940
rect 6736 598 6856 626
rect 7288 610 7316 16934
rect 8010 15192 8066 15201
rect 8010 15127 8066 15136
rect 8024 3534 8052 15127
rect 8012 3528 8064 3534
rect 8012 3470 8064 3476
rect 8484 610 8512 16934
rect 9588 16794 9616 17167
rect 10508 16998 10536 17682
rect 10496 16992 10548 16998
rect 10496 16934 10548 16940
rect 10001 16892 10297 16912
rect 10057 16890 10081 16892
rect 10137 16890 10161 16892
rect 10217 16890 10241 16892
rect 10079 16838 10081 16890
rect 10143 16838 10155 16890
rect 10217 16838 10219 16890
rect 10057 16836 10081 16838
rect 10137 16836 10161 16838
rect 10217 16836 10241 16838
rect 10001 16816 10297 16836
rect 9576 16788 9628 16794
rect 9576 16730 9628 16736
rect 9482 16688 9538 16697
rect 9482 16623 9538 16632
rect 9852 16652 9904 16658
rect 9496 16250 9524 16623
rect 9852 16594 9904 16600
rect 9484 16244 9536 16250
rect 9484 16186 9536 16192
rect 9864 15910 9892 16594
rect 9300 15904 9352 15910
rect 9300 15846 9352 15852
rect 9852 15904 9904 15910
rect 9852 15846 9904 15852
rect 8840 3528 8892 3534
rect 8840 3470 8892 3476
rect 9312 3482 9340 15846
rect 9864 15201 9892 15846
rect 10001 15804 10297 15824
rect 10057 15802 10081 15804
rect 10137 15802 10161 15804
rect 10217 15802 10241 15804
rect 10079 15750 10081 15802
rect 10143 15750 10155 15802
rect 10217 15750 10219 15802
rect 10057 15748 10081 15750
rect 10137 15748 10161 15750
rect 10217 15748 10241 15750
rect 10001 15728 10297 15748
rect 9850 15192 9906 15201
rect 9850 15127 9906 15136
rect 10001 14716 10297 14736
rect 10057 14714 10081 14716
rect 10137 14714 10161 14716
rect 10217 14714 10241 14716
rect 10079 14662 10081 14714
rect 10143 14662 10155 14714
rect 10217 14662 10219 14714
rect 10057 14660 10081 14662
rect 10137 14660 10161 14662
rect 10217 14660 10241 14662
rect 10001 14640 10297 14660
rect 10001 13628 10297 13648
rect 10057 13626 10081 13628
rect 10137 13626 10161 13628
rect 10217 13626 10241 13628
rect 10079 13574 10081 13626
rect 10143 13574 10155 13626
rect 10217 13574 10219 13626
rect 10057 13572 10081 13574
rect 10137 13572 10161 13574
rect 10217 13572 10241 13574
rect 10001 13552 10297 13572
rect 10001 12540 10297 12560
rect 10057 12538 10081 12540
rect 10137 12538 10161 12540
rect 10217 12538 10241 12540
rect 10079 12486 10081 12538
rect 10143 12486 10155 12538
rect 10217 12486 10219 12538
rect 10057 12484 10081 12486
rect 10137 12484 10161 12486
rect 10217 12484 10241 12486
rect 10001 12464 10297 12484
rect 10001 11452 10297 11472
rect 10057 11450 10081 11452
rect 10137 11450 10161 11452
rect 10217 11450 10241 11452
rect 10079 11398 10081 11450
rect 10143 11398 10155 11450
rect 10217 11398 10219 11450
rect 10057 11396 10081 11398
rect 10137 11396 10161 11398
rect 10217 11396 10241 11398
rect 10001 11376 10297 11396
rect 9390 11248 9446 11257
rect 9390 11183 9446 11192
rect 9404 3618 9432 11183
rect 10001 10364 10297 10384
rect 10057 10362 10081 10364
rect 10137 10362 10161 10364
rect 10217 10362 10241 10364
rect 10079 10310 10081 10362
rect 10143 10310 10155 10362
rect 10217 10310 10219 10362
rect 10057 10308 10081 10310
rect 10137 10308 10161 10310
rect 10217 10308 10241 10310
rect 10001 10288 10297 10308
rect 10001 9276 10297 9296
rect 10057 9274 10081 9276
rect 10137 9274 10161 9276
rect 10217 9274 10241 9276
rect 10079 9222 10081 9274
rect 10143 9222 10155 9274
rect 10217 9222 10219 9274
rect 10057 9220 10081 9222
rect 10137 9220 10161 9222
rect 10217 9220 10241 9222
rect 10001 9200 10297 9220
rect 10001 8188 10297 8208
rect 10057 8186 10081 8188
rect 10137 8186 10161 8188
rect 10217 8186 10241 8188
rect 10079 8134 10081 8186
rect 10143 8134 10155 8186
rect 10217 8134 10219 8186
rect 10057 8132 10081 8134
rect 10137 8132 10161 8134
rect 10217 8132 10241 8134
rect 10001 8112 10297 8132
rect 10001 7100 10297 7120
rect 10057 7098 10081 7100
rect 10137 7098 10161 7100
rect 10217 7098 10241 7100
rect 10079 7046 10081 7098
rect 10143 7046 10155 7098
rect 10217 7046 10219 7098
rect 10057 7044 10081 7046
rect 10137 7044 10161 7046
rect 10217 7044 10241 7046
rect 10001 7024 10297 7044
rect 10001 6012 10297 6032
rect 10057 6010 10081 6012
rect 10137 6010 10161 6012
rect 10217 6010 10241 6012
rect 10079 5958 10081 6010
rect 10143 5958 10155 6010
rect 10217 5958 10219 6010
rect 10057 5956 10081 5958
rect 10137 5956 10161 5958
rect 10217 5956 10241 5958
rect 10001 5936 10297 5956
rect 10001 4924 10297 4944
rect 10057 4922 10081 4924
rect 10137 4922 10161 4924
rect 10217 4922 10241 4924
rect 10079 4870 10081 4922
rect 10143 4870 10155 4922
rect 10217 4870 10219 4922
rect 10057 4868 10081 4870
rect 10137 4868 10161 4870
rect 10217 4868 10241 4870
rect 10001 4848 10297 4868
rect 10001 3836 10297 3856
rect 10057 3834 10081 3836
rect 10137 3834 10161 3836
rect 10217 3834 10241 3836
rect 10079 3782 10081 3834
rect 10143 3782 10155 3834
rect 10217 3782 10219 3834
rect 10057 3780 10081 3782
rect 10137 3780 10161 3782
rect 10217 3780 10241 3782
rect 10001 3760 10297 3780
rect 9404 3590 9708 3618
rect 6828 480 6856 598
rect 7276 604 7328 610
rect 7276 546 7328 552
rect 7460 604 7512 610
rect 7460 546 7512 552
rect 8104 604 8156 610
rect 8104 546 8156 552
rect 8472 604 8524 610
rect 8472 546 8524 552
rect 7472 480 7500 546
rect 8116 480 8144 546
rect 8852 480 8880 3470
rect 9312 3454 9524 3482
rect 9496 480 9524 3454
rect 9680 2394 9708 3590
rect 10508 3097 10536 16934
rect 10862 15464 10918 15473
rect 10862 15399 10918 15408
rect 10876 15162 10904 15399
rect 10864 15156 10916 15162
rect 10864 15098 10916 15104
rect 11140 14816 11192 14822
rect 11140 14758 11192 14764
rect 11048 14476 11100 14482
rect 11048 14418 11100 14424
rect 11060 13870 11088 14418
rect 11048 13864 11100 13870
rect 11048 13806 11100 13812
rect 10770 11520 10826 11529
rect 10770 11455 10826 11464
rect 10784 3534 10812 11455
rect 11060 4049 11088 13806
rect 11046 4040 11102 4049
rect 11046 3975 11102 3984
rect 10772 3528 10824 3534
rect 11152 3482 11180 14758
rect 11244 14618 11272 24890
rect 13636 20754 13664 27520
rect 19236 26376 19288 26382
rect 19236 26318 19288 26324
rect 13716 26308 13768 26314
rect 13716 26250 13768 26256
rect 13360 20726 13664 20754
rect 11232 14612 11284 14618
rect 11232 14554 11284 14560
rect 13360 14550 13388 20726
rect 13728 16250 13756 26250
rect 14668 25052 14964 25072
rect 14724 25050 14748 25052
rect 14804 25050 14828 25052
rect 14884 25050 14908 25052
rect 14746 24998 14748 25050
rect 14810 24998 14822 25050
rect 14884 24998 14886 25050
rect 14724 24996 14748 24998
rect 14804 24996 14828 24998
rect 14884 24996 14908 24998
rect 14668 24976 14964 24996
rect 14668 23964 14964 23984
rect 14724 23962 14748 23964
rect 14804 23962 14828 23964
rect 14884 23962 14908 23964
rect 14746 23910 14748 23962
rect 14810 23910 14822 23962
rect 14884 23910 14886 23962
rect 14724 23908 14748 23910
rect 14804 23908 14828 23910
rect 14884 23908 14908 23910
rect 14668 23888 14964 23908
rect 14452 22976 14504 22982
rect 14450 22944 14452 22953
rect 15096 22976 15148 22982
rect 14504 22944 14506 22953
rect 15094 22944 15096 22953
rect 15148 22944 15150 22953
rect 14450 22879 14506 22888
rect 14668 22876 14964 22896
rect 15094 22879 15150 22888
rect 14724 22874 14748 22876
rect 14804 22874 14828 22876
rect 14884 22874 14908 22876
rect 14746 22822 14748 22874
rect 14810 22822 14822 22874
rect 14884 22822 14886 22874
rect 14724 22820 14748 22822
rect 14804 22820 14828 22822
rect 14884 22820 14908 22822
rect 14668 22800 14964 22820
rect 14668 21788 14964 21808
rect 14724 21786 14748 21788
rect 14804 21786 14828 21788
rect 14884 21786 14908 21788
rect 14746 21734 14748 21786
rect 14810 21734 14822 21786
rect 14884 21734 14886 21786
rect 14724 21732 14748 21734
rect 14804 21732 14828 21734
rect 14884 21732 14908 21734
rect 14668 21712 14964 21732
rect 14174 21040 14230 21049
rect 14174 20975 14230 20984
rect 14188 20641 14216 20975
rect 14668 20700 14964 20720
rect 14724 20698 14748 20700
rect 14804 20698 14828 20700
rect 14884 20698 14908 20700
rect 14746 20646 14748 20698
rect 14810 20646 14822 20698
rect 14884 20646 14886 20698
rect 14724 20644 14748 20646
rect 14804 20644 14828 20646
rect 14884 20644 14908 20646
rect 14174 20632 14230 20641
rect 14668 20624 14964 20644
rect 14174 20567 14230 20576
rect 14668 19612 14964 19632
rect 14724 19610 14748 19612
rect 14804 19610 14828 19612
rect 14884 19610 14908 19612
rect 14746 19558 14748 19610
rect 14810 19558 14822 19610
rect 14884 19558 14886 19610
rect 14724 19556 14748 19558
rect 14804 19556 14828 19558
rect 14884 19556 14908 19558
rect 14668 19536 14964 19556
rect 14668 18524 14964 18544
rect 14724 18522 14748 18524
rect 14804 18522 14828 18524
rect 14884 18522 14908 18524
rect 14746 18470 14748 18522
rect 14810 18470 14822 18522
rect 14884 18470 14886 18522
rect 14724 18468 14748 18470
rect 14804 18468 14828 18470
rect 14884 18468 14908 18470
rect 14668 18448 14964 18468
rect 14668 17436 14964 17456
rect 14724 17434 14748 17436
rect 14804 17434 14828 17436
rect 14884 17434 14908 17436
rect 14746 17382 14748 17434
rect 14810 17382 14822 17434
rect 14884 17382 14886 17434
rect 14724 17380 14748 17382
rect 14804 17380 14828 17382
rect 14884 17380 14908 17382
rect 14668 17360 14964 17380
rect 16750 17368 16806 17377
rect 16750 17303 16806 17312
rect 16764 17105 16792 17303
rect 19248 17218 19276 26318
rect 19334 25596 19630 25616
rect 19390 25594 19414 25596
rect 19470 25594 19494 25596
rect 19550 25594 19574 25596
rect 19412 25542 19414 25594
rect 19476 25542 19488 25594
rect 19550 25542 19552 25594
rect 19390 25540 19414 25542
rect 19470 25540 19494 25542
rect 19550 25540 19574 25542
rect 19334 25520 19630 25540
rect 22928 24834 22956 27520
rect 23834 27503 23890 27512
rect 23848 26382 23876 27503
rect 24478 26888 24534 26897
rect 24478 26823 24534 26832
rect 23836 26376 23888 26382
rect 23836 26318 23888 26324
rect 24492 26314 24520 26823
rect 24480 26308 24532 26314
rect 24480 26250 24532 26256
rect 23834 26208 23890 26217
rect 23834 26143 23890 26152
rect 23848 24954 23876 26143
rect 24478 25528 24534 25537
rect 24478 25463 24534 25472
rect 24001 25052 24297 25072
rect 24057 25050 24081 25052
rect 24137 25050 24161 25052
rect 24217 25050 24241 25052
rect 24079 24998 24081 25050
rect 24143 24998 24155 25050
rect 24217 24998 24219 25050
rect 24057 24996 24081 24998
rect 24137 24996 24161 24998
rect 24217 24996 24241 24998
rect 24001 24976 24297 24996
rect 23836 24948 23888 24954
rect 23836 24890 23888 24896
rect 24492 24886 24520 25463
rect 24480 24880 24532 24886
rect 22192 24806 22956 24834
rect 23834 24848 23890 24857
rect 19334 24508 19630 24528
rect 19390 24506 19414 24508
rect 19470 24506 19494 24508
rect 19550 24506 19574 24508
rect 19412 24454 19414 24506
rect 19476 24454 19488 24506
rect 19550 24454 19552 24506
rect 19390 24452 19414 24454
rect 19470 24452 19494 24454
rect 19550 24452 19574 24454
rect 19334 24432 19630 24452
rect 19334 23420 19630 23440
rect 19390 23418 19414 23420
rect 19470 23418 19494 23420
rect 19550 23418 19574 23420
rect 19412 23366 19414 23418
rect 19476 23366 19488 23418
rect 19550 23366 19552 23418
rect 19390 23364 19414 23366
rect 19470 23364 19494 23366
rect 19550 23364 19574 23366
rect 19334 23344 19630 23364
rect 19334 22332 19630 22352
rect 19390 22330 19414 22332
rect 19470 22330 19494 22332
rect 19550 22330 19574 22332
rect 19412 22278 19414 22330
rect 19476 22278 19488 22330
rect 19550 22278 19552 22330
rect 19390 22276 19414 22278
rect 19470 22276 19494 22278
rect 19550 22276 19574 22278
rect 19334 22256 19630 22276
rect 19334 21244 19630 21264
rect 19390 21242 19414 21244
rect 19470 21242 19494 21244
rect 19550 21242 19574 21244
rect 19412 21190 19414 21242
rect 19476 21190 19488 21242
rect 19550 21190 19552 21242
rect 19390 21188 19414 21190
rect 19470 21188 19494 21190
rect 19550 21188 19574 21190
rect 19334 21168 19630 21188
rect 19334 20156 19630 20176
rect 19390 20154 19414 20156
rect 19470 20154 19494 20156
rect 19550 20154 19574 20156
rect 19412 20102 19414 20154
rect 19476 20102 19488 20154
rect 19550 20102 19552 20154
rect 19390 20100 19414 20102
rect 19470 20100 19494 20102
rect 19550 20100 19574 20102
rect 19334 20080 19630 20100
rect 19786 20088 19842 20097
rect 19786 20023 19842 20032
rect 19800 19417 19828 20023
rect 19786 19408 19842 19417
rect 19786 19343 19842 19352
rect 22192 19310 22220 24806
rect 24480 24822 24532 24828
rect 23834 24783 23890 24792
rect 23374 23488 23430 23497
rect 23374 23423 23430 23432
rect 23388 22001 23416 23423
rect 23848 23089 23876 24783
rect 24478 24168 24534 24177
rect 24478 24103 24534 24112
rect 24001 23964 24297 23984
rect 24057 23962 24081 23964
rect 24137 23962 24161 23964
rect 24217 23962 24241 23964
rect 24079 23910 24081 23962
rect 24143 23910 24155 23962
rect 24217 23910 24219 23962
rect 24057 23908 24081 23910
rect 24137 23908 24161 23910
rect 24217 23908 24241 23910
rect 24001 23888 24297 23908
rect 23834 23080 23890 23089
rect 23834 23015 23890 23024
rect 24001 22876 24297 22896
rect 24057 22874 24081 22876
rect 24137 22874 24161 22876
rect 24217 22874 24241 22876
rect 24079 22822 24081 22874
rect 24143 22822 24155 22874
rect 24217 22822 24219 22874
rect 24057 22820 24081 22822
rect 24137 22820 24161 22822
rect 24217 22820 24241 22822
rect 24001 22800 24297 22820
rect 24492 22545 24520 24103
rect 24478 22536 24534 22545
rect 24478 22471 24534 22480
rect 24478 22128 24534 22137
rect 24478 22063 24534 22072
rect 23374 21992 23430 22001
rect 23374 21927 23430 21936
rect 24001 21788 24297 21808
rect 24057 21786 24081 21788
rect 24137 21786 24161 21788
rect 24217 21786 24241 21788
rect 24079 21734 24081 21786
rect 24143 21734 24155 21786
rect 24217 21734 24219 21786
rect 24057 21732 24081 21734
rect 24137 21732 24161 21734
rect 24217 21732 24241 21734
rect 24001 21712 24297 21732
rect 24386 20768 24442 20777
rect 24001 20700 24297 20720
rect 24386 20703 24442 20712
rect 24057 20698 24081 20700
rect 24137 20698 24161 20700
rect 24217 20698 24241 20700
rect 24079 20646 24081 20698
rect 24143 20646 24155 20698
rect 24217 20646 24219 20698
rect 24057 20644 24081 20646
rect 24137 20644 24161 20646
rect 24217 20644 24241 20646
rect 24001 20624 24297 20644
rect 24400 19961 24428 20703
rect 24386 19952 24442 19961
rect 24386 19887 24442 19896
rect 24001 19612 24297 19632
rect 24057 19610 24081 19612
rect 24137 19610 24161 19612
rect 24217 19610 24241 19612
rect 24079 19558 24081 19610
rect 24143 19558 24155 19610
rect 24217 19558 24219 19610
rect 24057 19556 24081 19558
rect 24137 19556 24161 19558
rect 24217 19556 24241 19558
rect 24001 19536 24297 19556
rect 24386 19408 24442 19417
rect 24386 19343 24442 19352
rect 21996 19304 22048 19310
rect 21996 19246 22048 19252
rect 22180 19304 22232 19310
rect 22180 19246 22232 19252
rect 19334 19068 19630 19088
rect 19390 19066 19414 19068
rect 19470 19066 19494 19068
rect 19550 19066 19574 19068
rect 19412 19014 19414 19066
rect 19476 19014 19488 19066
rect 19550 19014 19552 19066
rect 19390 19012 19414 19014
rect 19470 19012 19494 19014
rect 19550 19012 19574 19014
rect 19334 18992 19630 19012
rect 19334 17980 19630 18000
rect 19390 17978 19414 17980
rect 19470 17978 19494 17980
rect 19550 17978 19574 17980
rect 19412 17926 19414 17978
rect 19476 17926 19488 17978
rect 19550 17926 19552 17978
rect 19390 17924 19414 17926
rect 19470 17924 19494 17926
rect 19550 17924 19574 17926
rect 19334 17904 19630 17924
rect 19156 17190 19276 17218
rect 16750 17096 16806 17105
rect 16750 17031 16806 17040
rect 14668 16348 14964 16368
rect 14724 16346 14748 16348
rect 14804 16346 14828 16348
rect 14884 16346 14908 16348
rect 14746 16294 14748 16346
rect 14810 16294 14822 16346
rect 14884 16294 14886 16346
rect 14724 16292 14748 16294
rect 14804 16292 14828 16294
rect 14884 16292 14908 16294
rect 14668 16272 14964 16292
rect 13716 16244 13768 16250
rect 13716 16186 13768 16192
rect 13808 15904 13860 15910
rect 13808 15846 13860 15852
rect 12520 14544 12572 14550
rect 12520 14486 12572 14492
rect 13348 14544 13400 14550
rect 13348 14486 13400 14492
rect 12428 14408 12480 14414
rect 12428 14350 12480 14356
rect 12440 13841 12468 14350
rect 12532 14074 12560 14486
rect 12520 14068 12572 14074
rect 12520 14010 12572 14016
rect 12426 13832 12482 13841
rect 12426 13767 12482 13776
rect 12794 13832 12850 13841
rect 12794 13767 12796 13776
rect 12848 13767 12850 13776
rect 12796 13738 12848 13744
rect 12808 13462 12836 13738
rect 12796 13456 12848 13462
rect 12796 13398 12848 13404
rect 12520 13388 12572 13394
rect 12520 13330 12572 13336
rect 12334 12744 12390 12753
rect 12334 12679 12390 12688
rect 12348 12646 12376 12679
rect 12336 12640 12388 12646
rect 12336 12582 12388 12588
rect 12532 12442 12560 13330
rect 12808 12986 12836 13398
rect 13624 13320 13676 13326
rect 13624 13262 13676 13268
rect 13636 12986 13664 13262
rect 12796 12980 12848 12986
rect 12796 12922 12848 12928
rect 13624 12980 13676 12986
rect 13624 12922 13676 12928
rect 12704 12776 12756 12782
rect 12704 12718 12756 12724
rect 12520 12436 12572 12442
rect 12520 12378 12572 12384
rect 12716 3534 12744 12718
rect 13532 12708 13584 12714
rect 13532 12650 13584 12656
rect 13544 11098 13572 12650
rect 13452 11070 13572 11098
rect 13452 3534 13480 11070
rect 10772 3470 10824 3476
rect 10876 3454 11180 3482
rect 11600 3528 11652 3534
rect 11600 3470 11652 3476
rect 12244 3528 12296 3534
rect 12244 3470 12296 3476
rect 12704 3528 12756 3534
rect 12704 3470 12756 3476
rect 12888 3528 12940 3534
rect 12888 3470 12940 3476
rect 13440 3528 13492 3534
rect 13440 3470 13492 3476
rect 10494 3088 10550 3097
rect 10494 3023 10550 3032
rect 10001 2748 10297 2768
rect 10057 2746 10081 2748
rect 10137 2746 10161 2748
rect 10217 2746 10241 2748
rect 10079 2694 10081 2746
rect 10143 2694 10155 2746
rect 10217 2694 10219 2746
rect 10057 2692 10081 2694
rect 10137 2692 10161 2694
rect 10217 2692 10241 2694
rect 10001 2672 10297 2692
rect 9680 2366 10260 2394
rect 10232 480 10260 2366
rect 10876 480 10904 3454
rect 11612 480 11640 3470
rect 12256 480 12284 3470
rect 12900 480 12928 3470
rect 13820 610 13848 15846
rect 17946 15464 18002 15473
rect 17946 15399 18002 15408
rect 14668 15260 14964 15280
rect 14724 15258 14748 15260
rect 14804 15258 14828 15260
rect 14884 15258 14908 15260
rect 14746 15206 14748 15258
rect 14810 15206 14822 15258
rect 14884 15206 14886 15258
rect 14724 15204 14748 15206
rect 14804 15204 14828 15206
rect 14884 15204 14908 15206
rect 14668 15184 14964 15204
rect 17960 15162 17988 15399
rect 17948 15156 18000 15162
rect 17948 15098 18000 15104
rect 15648 14884 15700 14890
rect 15648 14826 15700 14832
rect 15660 14618 15688 14826
rect 15648 14612 15700 14618
rect 15648 14554 15700 14560
rect 16292 14476 16344 14482
rect 16292 14418 16344 14424
rect 18132 14476 18184 14482
rect 18132 14418 18184 14424
rect 16108 14408 16160 14414
rect 16108 14350 16160 14356
rect 16200 14408 16252 14414
rect 16200 14350 16252 14356
rect 14176 14272 14228 14278
rect 14176 14214 14228 14220
rect 13900 13796 13952 13802
rect 13900 13738 13952 13744
rect 13912 13530 13940 13738
rect 13900 13524 13952 13530
rect 13900 13466 13952 13472
rect 14188 13394 14216 14214
rect 14668 14172 14964 14192
rect 14724 14170 14748 14172
rect 14804 14170 14828 14172
rect 14884 14170 14908 14172
rect 14746 14118 14748 14170
rect 14810 14118 14822 14170
rect 14884 14118 14886 14170
rect 14724 14116 14748 14118
rect 14804 14116 14828 14118
rect 14884 14116 14908 14118
rect 14668 14096 14964 14116
rect 15462 13968 15518 13977
rect 16120 13938 16148 14350
rect 15462 13903 15518 13912
rect 16108 13932 16160 13938
rect 14268 13864 14320 13870
rect 14268 13806 14320 13812
rect 14360 13864 14412 13870
rect 14360 13806 14412 13812
rect 14176 13388 14228 13394
rect 14176 13330 14228 13336
rect 14188 12850 14216 13330
rect 14280 12918 14308 13806
rect 14268 12912 14320 12918
rect 14268 12854 14320 12860
rect 14176 12844 14228 12850
rect 14176 12786 14228 12792
rect 14084 12640 14136 12646
rect 14084 12582 14136 12588
rect 14096 12102 14124 12582
rect 14188 12442 14216 12786
rect 14176 12436 14228 12442
rect 14176 12378 14228 12384
rect 14084 12096 14136 12102
rect 14084 12038 14136 12044
rect 14372 11830 14400 13806
rect 15372 13388 15424 13394
rect 15372 13330 15424 13336
rect 14544 13252 14596 13258
rect 14544 13194 14596 13200
rect 14452 12980 14504 12986
rect 14452 12922 14504 12928
rect 14360 11824 14412 11830
rect 14360 11766 14412 11772
rect 14464 11762 14492 12922
rect 14556 12238 14584 13194
rect 14668 13084 14964 13104
rect 14724 13082 14748 13084
rect 14804 13082 14828 13084
rect 14884 13082 14908 13084
rect 14746 13030 14748 13082
rect 14810 13030 14822 13082
rect 14884 13030 14886 13082
rect 14724 13028 14748 13030
rect 14804 13028 14828 13030
rect 14884 13028 14908 13030
rect 14668 13008 14964 13028
rect 15384 12986 15412 13330
rect 15372 12980 15424 12986
rect 15372 12922 15424 12928
rect 15476 12866 15504 13903
rect 16108 13874 16160 13880
rect 15740 13796 15792 13802
rect 15740 13738 15792 13744
rect 15648 13728 15700 13734
rect 15648 13670 15700 13676
rect 15660 13530 15688 13670
rect 15648 13524 15700 13530
rect 15648 13466 15700 13472
rect 15384 12838 15504 12866
rect 15384 12442 15412 12838
rect 15660 12714 15688 13466
rect 15752 13326 15780 13738
rect 16212 13530 16240 14350
rect 16304 13870 16332 14418
rect 17764 14408 17816 14414
rect 17764 14350 17816 14356
rect 17672 13932 17724 13938
rect 17672 13874 17724 13880
rect 16292 13864 16344 13870
rect 16292 13806 16344 13812
rect 16200 13524 16252 13530
rect 16200 13466 16252 13472
rect 15740 13320 15792 13326
rect 15740 13262 15792 13268
rect 15648 12708 15700 12714
rect 15648 12650 15700 12656
rect 15372 12436 15424 12442
rect 15372 12378 15424 12384
rect 15660 12374 15688 12650
rect 15752 12442 15780 13262
rect 16212 12986 16240 13466
rect 16200 12980 16252 12986
rect 16200 12922 16252 12928
rect 15740 12436 15792 12442
rect 15740 12378 15792 12384
rect 15648 12368 15700 12374
rect 15648 12310 15700 12316
rect 14544 12232 14596 12238
rect 14544 12174 14596 12180
rect 14556 11898 14584 12174
rect 15188 12096 15240 12102
rect 15188 12038 15240 12044
rect 14668 11996 14964 12016
rect 14724 11994 14748 11996
rect 14804 11994 14828 11996
rect 14884 11994 14908 11996
rect 14746 11942 14748 11994
rect 14810 11942 14822 11994
rect 14884 11942 14886 11994
rect 14724 11940 14748 11942
rect 14804 11940 14828 11942
rect 14884 11940 14908 11942
rect 14668 11920 14964 11940
rect 14544 11892 14596 11898
rect 14544 11834 14596 11840
rect 14452 11756 14504 11762
rect 14452 11698 14504 11704
rect 15200 11558 15228 12038
rect 15660 11762 15688 12310
rect 15740 12300 15792 12306
rect 15740 12242 15792 12248
rect 15752 11898 15780 12242
rect 15740 11892 15792 11898
rect 15740 11834 15792 11840
rect 16304 11762 16332 13806
rect 17684 13682 17712 13874
rect 17408 13654 17712 13682
rect 17408 13326 17436 13654
rect 17396 13320 17448 13326
rect 17396 13262 17448 13268
rect 16568 12980 16620 12986
rect 16568 12922 16620 12928
rect 16384 12776 16436 12782
rect 16384 12718 16436 12724
rect 16396 12306 16424 12718
rect 16580 12306 16608 12922
rect 17408 12782 17436 13262
rect 17672 12980 17724 12986
rect 17672 12922 17724 12928
rect 17396 12776 17448 12782
rect 17396 12718 17448 12724
rect 16384 12300 16436 12306
rect 16384 12242 16436 12248
rect 16568 12300 16620 12306
rect 16568 12242 16620 12248
rect 17120 12300 17172 12306
rect 17120 12242 17172 12248
rect 17132 11898 17160 12242
rect 17120 11892 17172 11898
rect 17120 11834 17172 11840
rect 17408 11830 17436 12718
rect 17684 12442 17712 12922
rect 17672 12436 17724 12442
rect 17672 12378 17724 12384
rect 17776 11898 17804 14350
rect 18144 14074 18172 14418
rect 18776 14272 18828 14278
rect 18776 14214 18828 14220
rect 18132 14068 18184 14074
rect 18132 14010 18184 14016
rect 18040 13388 18092 13394
rect 18040 13330 18092 13336
rect 18052 12986 18080 13330
rect 18040 12980 18092 12986
rect 18040 12922 18092 12928
rect 18144 12850 18172 14010
rect 18788 13802 18816 14214
rect 18776 13796 18828 13802
rect 18776 13738 18828 13744
rect 19052 13796 19104 13802
rect 19052 13738 19104 13744
rect 18788 13530 18816 13738
rect 18776 13524 18828 13530
rect 18776 13466 18828 13472
rect 19064 12986 19092 13738
rect 18316 12980 18368 12986
rect 18316 12922 18368 12928
rect 19052 12980 19104 12986
rect 19052 12922 19104 12928
rect 18132 12844 18184 12850
rect 18132 12786 18184 12792
rect 17764 11892 17816 11898
rect 17764 11834 17816 11840
rect 17396 11824 17448 11830
rect 17396 11766 17448 11772
rect 18328 11762 18356 12922
rect 18868 12708 18920 12714
rect 18868 12650 18920 12656
rect 18776 12300 18828 12306
rect 18776 12242 18828 12248
rect 15648 11756 15700 11762
rect 15648 11698 15700 11704
rect 16292 11756 16344 11762
rect 16292 11698 16344 11704
rect 18316 11756 18368 11762
rect 18316 11698 18368 11704
rect 14544 11552 14596 11558
rect 14542 11520 14544 11529
rect 15188 11552 15240 11558
rect 14596 11520 14598 11529
rect 15188 11494 15240 11500
rect 17488 11552 17540 11558
rect 17488 11494 17540 11500
rect 14542 11455 14598 11464
rect 15200 11286 15228 11494
rect 15188 11280 15240 11286
rect 17500 11257 17528 11494
rect 18328 11354 18356 11698
rect 18788 11558 18816 12242
rect 18776 11552 18828 11558
rect 18776 11494 18828 11500
rect 18316 11348 18368 11354
rect 18316 11290 18368 11296
rect 15188 11222 15240 11228
rect 17486 11248 17542 11257
rect 17486 11183 17542 11192
rect 14668 10908 14964 10928
rect 14724 10906 14748 10908
rect 14804 10906 14828 10908
rect 14884 10906 14908 10908
rect 14746 10854 14748 10906
rect 14810 10854 14822 10906
rect 14884 10854 14886 10906
rect 14724 10852 14748 10854
rect 14804 10852 14828 10854
rect 14884 10852 14908 10854
rect 14668 10832 14964 10852
rect 18684 10600 18736 10606
rect 15278 10568 15334 10577
rect 18684 10542 18736 10548
rect 15278 10503 15280 10512
rect 15332 10503 15334 10512
rect 18040 10532 18092 10538
rect 15280 10474 15332 10480
rect 18040 10474 18092 10480
rect 14544 10464 14596 10470
rect 14544 10406 14596 10412
rect 14452 9376 14504 9382
rect 14452 9318 14504 9324
rect 14464 8634 14492 9318
rect 14452 8628 14504 8634
rect 14452 8570 14504 8576
rect 14268 8560 14320 8566
rect 14268 8502 14320 8508
rect 13624 604 13676 610
rect 13624 546 13676 552
rect 13808 604 13860 610
rect 13808 546 13860 552
rect 13636 480 13664 546
rect 14280 480 14308 8502
rect 14556 4162 14584 10406
rect 14668 9820 14964 9840
rect 14724 9818 14748 9820
rect 14804 9818 14828 9820
rect 14884 9818 14908 9820
rect 14746 9766 14748 9818
rect 14810 9766 14822 9818
rect 14884 9766 14886 9818
rect 14724 9764 14748 9766
rect 14804 9764 14828 9766
rect 14884 9764 14908 9766
rect 14668 9744 14964 9764
rect 18052 9722 18080 10474
rect 18696 10470 18724 10542
rect 18684 10464 18736 10470
rect 18684 10406 18736 10412
rect 18040 9716 18092 9722
rect 18040 9658 18092 9664
rect 14910 9616 14966 9625
rect 14910 9551 14912 9560
rect 14964 9551 14966 9560
rect 14912 9522 14964 9528
rect 18696 9518 18724 10406
rect 18684 9512 18736 9518
rect 18684 9454 18736 9460
rect 18406 9072 18462 9081
rect 16016 9036 16068 9042
rect 18406 9007 18462 9016
rect 18684 9036 18736 9042
rect 16016 8978 16068 8984
rect 14668 8732 14964 8752
rect 14724 8730 14748 8732
rect 14804 8730 14828 8732
rect 14884 8730 14908 8732
rect 14746 8678 14748 8730
rect 14810 8678 14822 8730
rect 14884 8678 14886 8730
rect 14724 8676 14748 8678
rect 14804 8676 14828 8678
rect 14884 8676 14908 8678
rect 14668 8656 14964 8676
rect 16028 8566 16056 8978
rect 16200 8832 16252 8838
rect 16200 8774 16252 8780
rect 17580 8832 17632 8838
rect 17580 8774 17632 8780
rect 16016 8560 16068 8566
rect 16014 8528 16016 8537
rect 16068 8528 16070 8537
rect 16014 8463 16070 8472
rect 14668 7644 14964 7664
rect 14724 7642 14748 7644
rect 14804 7642 14828 7644
rect 14884 7642 14908 7644
rect 14746 7590 14748 7642
rect 14810 7590 14822 7642
rect 14884 7590 14886 7642
rect 14724 7588 14748 7590
rect 14804 7588 14828 7590
rect 14884 7588 14908 7590
rect 14668 7568 14964 7588
rect 15648 7200 15700 7206
rect 15648 7142 15700 7148
rect 14668 6556 14964 6576
rect 14724 6554 14748 6556
rect 14804 6554 14828 6556
rect 14884 6554 14908 6556
rect 14746 6502 14748 6554
rect 14810 6502 14822 6554
rect 14884 6502 14886 6554
rect 14724 6500 14748 6502
rect 14804 6500 14828 6502
rect 14884 6500 14908 6502
rect 14668 6480 14964 6500
rect 14668 5468 14964 5488
rect 14724 5466 14748 5468
rect 14804 5466 14828 5468
rect 14884 5466 14908 5468
rect 14746 5414 14748 5466
rect 14810 5414 14822 5466
rect 14884 5414 14886 5466
rect 14724 5412 14748 5414
rect 14804 5412 14828 5414
rect 14884 5412 14908 5414
rect 14668 5392 14964 5412
rect 14668 4380 14964 4400
rect 14724 4378 14748 4380
rect 14804 4378 14828 4380
rect 14884 4378 14908 4380
rect 14746 4326 14748 4378
rect 14810 4326 14822 4378
rect 14884 4326 14886 4378
rect 14724 4324 14748 4326
rect 14804 4324 14828 4326
rect 14884 4324 14908 4326
rect 14668 4304 14964 4324
rect 14556 4134 15044 4162
rect 14668 3292 14964 3312
rect 14724 3290 14748 3292
rect 14804 3290 14828 3292
rect 14884 3290 14908 3292
rect 14746 3238 14748 3290
rect 14810 3238 14822 3290
rect 14884 3238 14886 3290
rect 14724 3236 14748 3238
rect 14804 3236 14828 3238
rect 14884 3236 14908 3238
rect 14668 3216 14964 3236
rect 14668 2204 14964 2224
rect 14724 2202 14748 2204
rect 14804 2202 14828 2204
rect 14884 2202 14908 2204
rect 14746 2150 14748 2202
rect 14810 2150 14822 2202
rect 14884 2150 14886 2202
rect 14724 2148 14748 2150
rect 14804 2148 14828 2150
rect 14884 2148 14908 2150
rect 14668 2128 14964 2148
rect 15016 480 15044 4134
rect 15660 480 15688 7142
rect 16212 4026 16240 8774
rect 17592 7954 17620 8774
rect 17854 7984 17910 7993
rect 16752 7948 16804 7954
rect 16752 7890 16804 7896
rect 17580 7948 17632 7954
rect 17854 7919 17910 7928
rect 17580 7890 17632 7896
rect 16384 7744 16436 7750
rect 16384 7686 16436 7692
rect 16396 7546 16424 7686
rect 16764 7546 16792 7890
rect 16384 7540 16436 7546
rect 16384 7482 16436 7488
rect 16752 7540 16804 7546
rect 16752 7482 16804 7488
rect 16396 7342 16424 7482
rect 16384 7336 16436 7342
rect 16384 7278 16436 7284
rect 17672 7200 17724 7206
rect 17672 7142 17724 7148
rect 16936 5772 16988 5778
rect 16936 5714 16988 5720
rect 16948 5370 16976 5714
rect 17028 5568 17080 5574
rect 17028 5510 17080 5516
rect 16936 5364 16988 5370
rect 16936 5306 16988 5312
rect 16212 3998 16332 4026
rect 16304 480 16332 3998
rect 17040 480 17068 5510
rect 17684 480 17712 7142
rect 17868 6866 17896 7919
rect 18420 7546 18448 9007
rect 18684 8978 18736 8984
rect 18696 8634 18724 8978
rect 18684 8628 18736 8634
rect 18684 8570 18736 8576
rect 18408 7540 18460 7546
rect 18408 7482 18460 7488
rect 18420 7342 18448 7482
rect 18408 7336 18460 7342
rect 18408 7278 18460 7284
rect 17856 6860 17908 6866
rect 17856 6802 17908 6808
rect 17868 6458 17896 6802
rect 18408 6656 18460 6662
rect 18408 6598 18460 6604
rect 18500 6656 18552 6662
rect 18500 6598 18552 6604
rect 17856 6452 17908 6458
rect 17856 6394 17908 6400
rect 18132 5772 18184 5778
rect 18132 5714 18184 5720
rect 18144 5370 18172 5714
rect 18132 5364 18184 5370
rect 18132 5306 18184 5312
rect 18420 480 18448 6598
rect 18512 5778 18540 6598
rect 18500 5772 18552 5778
rect 18500 5714 18552 5720
rect 18788 3641 18816 11494
rect 18880 11354 18908 12650
rect 19156 12442 19184 17190
rect 19334 16892 19630 16912
rect 19390 16890 19414 16892
rect 19470 16890 19494 16892
rect 19550 16890 19574 16892
rect 19412 16838 19414 16890
rect 19476 16838 19488 16890
rect 19550 16838 19552 16890
rect 19390 16836 19414 16838
rect 19470 16836 19494 16838
rect 19550 16836 19574 16838
rect 19334 16816 19630 16836
rect 19694 16688 19750 16697
rect 19694 16623 19750 16632
rect 19334 15804 19630 15824
rect 19390 15802 19414 15804
rect 19470 15802 19494 15804
rect 19550 15802 19574 15804
rect 19412 15750 19414 15802
rect 19476 15750 19488 15802
rect 19550 15750 19552 15802
rect 19390 15748 19414 15750
rect 19470 15748 19494 15750
rect 19550 15748 19574 15750
rect 19334 15728 19630 15748
rect 19708 15162 19736 16623
rect 21718 15600 21774 15609
rect 21718 15535 21774 15544
rect 21732 15337 21760 15535
rect 21718 15328 21774 15337
rect 21718 15263 21774 15272
rect 19696 15156 19748 15162
rect 19696 15098 19748 15104
rect 19696 14952 19748 14958
rect 19696 14894 19748 14900
rect 19334 14716 19630 14736
rect 19390 14714 19414 14716
rect 19470 14714 19494 14716
rect 19550 14714 19574 14716
rect 19412 14662 19414 14714
rect 19476 14662 19488 14714
rect 19550 14662 19552 14714
rect 19390 14660 19414 14662
rect 19470 14660 19494 14662
rect 19550 14660 19574 14662
rect 19334 14640 19630 14660
rect 19708 14618 19736 14894
rect 19696 14612 19748 14618
rect 19696 14554 19748 14560
rect 19236 14544 19288 14550
rect 19236 14486 19288 14492
rect 19248 13530 19276 14486
rect 19788 13728 19840 13734
rect 19788 13670 19840 13676
rect 19334 13628 19630 13648
rect 19390 13626 19414 13628
rect 19470 13626 19494 13628
rect 19550 13626 19574 13628
rect 19412 13574 19414 13626
rect 19476 13574 19488 13626
rect 19550 13574 19552 13626
rect 19390 13572 19414 13574
rect 19470 13572 19494 13574
rect 19550 13572 19574 13574
rect 19334 13552 19630 13572
rect 19236 13524 19288 13530
rect 19236 13466 19288 13472
rect 19236 12980 19288 12986
rect 19236 12922 19288 12928
rect 19248 12850 19276 12922
rect 19236 12844 19288 12850
rect 19236 12786 19288 12792
rect 19144 12436 19196 12442
rect 19144 12378 19196 12384
rect 19156 11778 19184 12378
rect 19064 11750 19184 11778
rect 19064 11694 19092 11750
rect 19248 11694 19276 12786
rect 19800 12782 19828 13670
rect 20616 13320 20668 13326
rect 20616 13262 20668 13268
rect 19788 12776 19840 12782
rect 19788 12718 19840 12724
rect 19334 12540 19630 12560
rect 19390 12538 19414 12540
rect 19470 12538 19494 12540
rect 19550 12538 19574 12540
rect 19412 12486 19414 12538
rect 19476 12486 19488 12538
rect 19550 12486 19552 12538
rect 19390 12484 19414 12486
rect 19470 12484 19494 12486
rect 19550 12484 19574 12486
rect 19334 12464 19630 12484
rect 19800 12238 19828 12718
rect 20628 12442 20656 13262
rect 21168 12640 21220 12646
rect 21168 12582 21220 12588
rect 21718 12608 21774 12617
rect 20616 12436 20668 12442
rect 20616 12378 20668 12384
rect 21180 12238 21208 12582
rect 21718 12543 21774 12552
rect 21352 12436 21404 12442
rect 21352 12378 21404 12384
rect 19788 12232 19840 12238
rect 19788 12174 19840 12180
rect 21168 12232 21220 12238
rect 21168 12174 21220 12180
rect 21180 11830 21208 12174
rect 21364 11898 21392 12378
rect 21732 12170 21760 12543
rect 21720 12164 21772 12170
rect 21720 12106 21772 12112
rect 21352 11892 21404 11898
rect 21352 11834 21404 11840
rect 21168 11824 21220 11830
rect 21168 11766 21220 11772
rect 19052 11688 19104 11694
rect 19052 11630 19104 11636
rect 19236 11688 19288 11694
rect 19236 11630 19288 11636
rect 19064 11354 19092 11630
rect 19788 11620 19840 11626
rect 19788 11562 19840 11568
rect 19334 11452 19630 11472
rect 19390 11450 19414 11452
rect 19470 11450 19494 11452
rect 19550 11450 19574 11452
rect 19412 11398 19414 11450
rect 19476 11398 19488 11450
rect 19550 11398 19552 11450
rect 19390 11396 19414 11398
rect 19470 11396 19494 11398
rect 19550 11396 19574 11398
rect 19334 11376 19630 11396
rect 19800 11354 19828 11562
rect 20248 11552 20300 11558
rect 20248 11494 20300 11500
rect 20432 11552 20484 11558
rect 20432 11494 20484 11500
rect 18868 11348 18920 11354
rect 18868 11290 18920 11296
rect 19052 11348 19104 11354
rect 19052 11290 19104 11296
rect 19788 11348 19840 11354
rect 19788 11290 19840 11296
rect 19800 11082 19828 11290
rect 20260 11150 20288 11494
rect 20248 11144 20300 11150
rect 20248 11086 20300 11092
rect 19788 11076 19840 11082
rect 19788 11018 19840 11024
rect 19236 11008 19288 11014
rect 19236 10950 19288 10956
rect 19248 10130 19276 10950
rect 19696 10600 19748 10606
rect 19696 10542 19748 10548
rect 19334 10364 19630 10384
rect 19390 10362 19414 10364
rect 19470 10362 19494 10364
rect 19550 10362 19574 10364
rect 19412 10310 19414 10362
rect 19476 10310 19488 10362
rect 19550 10310 19552 10362
rect 19390 10308 19414 10310
rect 19470 10308 19494 10310
rect 19550 10308 19574 10310
rect 19334 10288 19630 10308
rect 19236 10124 19288 10130
rect 19236 10066 19288 10072
rect 19052 9988 19104 9994
rect 19052 9930 19104 9936
rect 18868 9920 18920 9926
rect 18868 9862 18920 9868
rect 18880 9625 18908 9862
rect 18958 9752 19014 9761
rect 18958 9687 19014 9696
rect 18866 9616 18922 9625
rect 18866 9551 18922 9560
rect 18868 9376 18920 9382
rect 18868 9318 18920 9324
rect 18880 8430 18908 9318
rect 18972 9178 19000 9687
rect 19064 9450 19092 9930
rect 19248 9722 19276 10066
rect 19708 10062 19736 10542
rect 20260 10418 20288 11086
rect 20444 10690 20472 11494
rect 21180 11286 21208 11766
rect 21168 11280 21220 11286
rect 21168 11222 21220 11228
rect 21074 10976 21130 10985
rect 21074 10911 21130 10920
rect 20352 10662 20472 10690
rect 20352 10606 20380 10662
rect 20340 10600 20392 10606
rect 20340 10542 20392 10548
rect 20984 10600 21036 10606
rect 20984 10542 21036 10548
rect 20432 10464 20484 10470
rect 20260 10390 20380 10418
rect 20432 10406 20484 10412
rect 19696 10056 19748 10062
rect 19696 9998 19748 10004
rect 20352 9926 20380 10390
rect 20444 10062 20472 10406
rect 20996 10130 21024 10542
rect 21088 10266 21116 10911
rect 21536 10464 21588 10470
rect 21536 10406 21588 10412
rect 21076 10260 21128 10266
rect 21076 10202 21128 10208
rect 20984 10124 21036 10130
rect 20984 10066 21036 10072
rect 20432 10056 20484 10062
rect 20432 9998 20484 10004
rect 20340 9920 20392 9926
rect 20340 9862 20392 9868
rect 19236 9716 19288 9722
rect 19236 9658 19288 9664
rect 20352 9518 20380 9862
rect 20340 9512 20392 9518
rect 20340 9454 20392 9460
rect 20444 9450 20472 9998
rect 20616 9920 20668 9926
rect 20616 9862 20668 9868
rect 20628 9761 20656 9862
rect 20614 9752 20670 9761
rect 20614 9687 20670 9696
rect 19052 9444 19104 9450
rect 19052 9386 19104 9392
rect 20432 9444 20484 9450
rect 20432 9386 20484 9392
rect 20248 9376 20300 9382
rect 20248 9318 20300 9324
rect 19334 9276 19630 9296
rect 19390 9274 19414 9276
rect 19470 9274 19494 9276
rect 19550 9274 19574 9276
rect 19412 9222 19414 9274
rect 19476 9222 19488 9274
rect 19550 9222 19552 9274
rect 19390 9220 19414 9222
rect 19470 9220 19494 9222
rect 19550 9220 19574 9222
rect 19334 9200 19630 9220
rect 20260 9178 20288 9318
rect 20444 9178 20472 9386
rect 20996 9382 21024 10066
rect 21088 9722 21116 10202
rect 21548 10198 21576 10406
rect 21536 10192 21588 10198
rect 21536 10134 21588 10140
rect 22008 9722 22036 19246
rect 23650 18728 23706 18737
rect 23650 18663 23706 18672
rect 23664 17377 23692 18663
rect 24001 18524 24297 18544
rect 24057 18522 24081 18524
rect 24137 18522 24161 18524
rect 24217 18522 24241 18524
rect 24079 18470 24081 18522
rect 24143 18470 24155 18522
rect 24217 18470 24219 18522
rect 24057 18468 24081 18470
rect 24137 18468 24161 18470
rect 24217 18468 24241 18470
rect 24001 18448 24297 18468
rect 23926 18048 23982 18057
rect 23926 17983 23982 17992
rect 23650 17368 23706 17377
rect 23650 17303 23706 17312
rect 23940 17241 23968 17983
rect 24400 17649 24428 19343
rect 24386 17640 24442 17649
rect 24386 17575 24442 17584
rect 24001 17436 24297 17456
rect 24057 17434 24081 17436
rect 24137 17434 24161 17436
rect 24217 17434 24241 17436
rect 24079 17382 24081 17434
rect 24143 17382 24155 17434
rect 24217 17382 24219 17434
rect 24057 17380 24081 17382
rect 24137 17380 24161 17382
rect 24217 17380 24241 17382
rect 24001 17360 24297 17380
rect 23926 17232 23982 17241
rect 23926 17167 23982 17176
rect 24001 16348 24297 16368
rect 24057 16346 24081 16348
rect 24137 16346 24161 16348
rect 24217 16346 24241 16348
rect 24079 16294 24081 16346
rect 24143 16294 24155 16346
rect 24217 16294 24219 16346
rect 24057 16292 24081 16294
rect 24137 16292 24161 16294
rect 24217 16292 24241 16294
rect 24001 16272 24297 16292
rect 24001 15260 24297 15280
rect 24057 15258 24081 15260
rect 24137 15258 24161 15260
rect 24217 15258 24241 15260
rect 24079 15206 24081 15258
rect 24143 15206 24155 15258
rect 24217 15206 24219 15258
rect 24057 15204 24081 15206
rect 24137 15204 24161 15206
rect 24217 15204 24241 15206
rect 24001 15184 24297 15204
rect 23834 14648 23890 14657
rect 24492 14618 24520 22063
rect 23834 14583 23890 14592
rect 24480 14612 24532 14618
rect 23560 13388 23612 13394
rect 23560 13330 23612 13336
rect 23572 12782 23600 13330
rect 23848 13025 23876 14583
rect 24480 14554 24532 14560
rect 24388 14476 24440 14482
rect 24388 14418 24440 14424
rect 24001 14172 24297 14192
rect 24057 14170 24081 14172
rect 24137 14170 24161 14172
rect 24217 14170 24241 14172
rect 24079 14118 24081 14170
rect 24143 14118 24155 14170
rect 24217 14118 24219 14170
rect 24057 14116 24081 14118
rect 24137 14116 24161 14118
rect 24217 14116 24241 14118
rect 24001 14096 24297 14116
rect 24400 13954 24428 14418
rect 24308 13926 24428 13954
rect 24308 13734 24336 13926
rect 24296 13728 24348 13734
rect 24296 13670 24348 13676
rect 24308 13530 24336 13670
rect 24296 13524 24348 13530
rect 24296 13466 24348 13472
rect 24478 13288 24534 13297
rect 24478 13223 24534 13232
rect 24001 13084 24297 13104
rect 24057 13082 24081 13084
rect 24137 13082 24161 13084
rect 24217 13082 24241 13084
rect 24079 13030 24081 13082
rect 24143 13030 24155 13082
rect 24217 13030 24219 13082
rect 24057 13028 24081 13030
rect 24137 13028 24161 13030
rect 24217 13028 24241 13030
rect 23834 13016 23890 13025
rect 24001 13008 24297 13028
rect 23834 12951 23890 12960
rect 23560 12776 23612 12782
rect 23558 12744 23560 12753
rect 23612 12744 23614 12753
rect 23558 12679 23614 12688
rect 23190 12608 23246 12617
rect 23190 12543 23246 12552
rect 22088 12368 22140 12374
rect 22088 12310 22140 12316
rect 22100 11898 22128 12310
rect 22088 11892 22140 11898
rect 22088 11834 22140 11840
rect 22364 11008 22416 11014
rect 22364 10950 22416 10956
rect 22376 10674 22404 10950
rect 23204 10690 23232 12543
rect 24001 11996 24297 12016
rect 24057 11994 24081 11996
rect 24137 11994 24161 11996
rect 24217 11994 24241 11996
rect 24079 11942 24081 11994
rect 24143 11942 24155 11994
rect 24217 11942 24219 11994
rect 24057 11940 24081 11942
rect 24137 11940 24161 11942
rect 24217 11940 24241 11942
rect 24001 11920 24297 11940
rect 23742 11792 23798 11801
rect 23742 11727 23798 11736
rect 22364 10668 22416 10674
rect 22364 10610 22416 10616
rect 23112 10662 23232 10690
rect 22376 10266 22404 10610
rect 23112 10606 23140 10662
rect 23100 10600 23152 10606
rect 23756 10577 23784 11727
rect 24492 11694 24520 13223
rect 24480 11688 24532 11694
rect 24480 11630 24532 11636
rect 24480 11552 24532 11558
rect 24480 11494 24532 11500
rect 24001 10908 24297 10928
rect 24057 10906 24081 10908
rect 24137 10906 24161 10908
rect 24217 10906 24241 10908
rect 24079 10854 24081 10906
rect 24143 10854 24155 10906
rect 24217 10854 24219 10906
rect 24057 10852 24081 10854
rect 24137 10852 24161 10854
rect 24217 10852 24241 10854
rect 24001 10832 24297 10852
rect 23100 10542 23152 10548
rect 23742 10568 23798 10577
rect 23742 10503 23798 10512
rect 23926 10568 23982 10577
rect 23926 10503 23982 10512
rect 22364 10260 22416 10266
rect 22364 10202 22416 10208
rect 23190 10024 23246 10033
rect 23190 9959 23246 9968
rect 21076 9716 21128 9722
rect 21076 9658 21128 9664
rect 21996 9716 22048 9722
rect 21996 9658 22048 9664
rect 22272 9716 22324 9722
rect 22272 9658 22324 9664
rect 20984 9376 21036 9382
rect 20984 9318 21036 9324
rect 21352 9376 21404 9382
rect 21352 9318 21404 9324
rect 18960 9172 19012 9178
rect 18960 9114 19012 9120
rect 20248 9172 20300 9178
rect 20248 9114 20300 9120
rect 20432 9172 20484 9178
rect 20432 9114 20484 9120
rect 18868 8424 18920 8430
rect 18868 8366 18920 8372
rect 18972 8090 19000 9114
rect 19420 8968 19472 8974
rect 19420 8910 19472 8916
rect 19432 8430 19460 8910
rect 19052 8424 19104 8430
rect 19052 8366 19104 8372
rect 19420 8424 19472 8430
rect 19420 8366 19472 8372
rect 19064 8294 19092 8366
rect 19052 8288 19104 8294
rect 19052 8230 19104 8236
rect 21260 8288 21312 8294
rect 21260 8230 21312 8236
rect 18960 8084 19012 8090
rect 18960 8026 19012 8032
rect 19064 7342 19092 8230
rect 19334 8188 19630 8208
rect 19390 8186 19414 8188
rect 19470 8186 19494 8188
rect 19550 8186 19574 8188
rect 19412 8134 19414 8186
rect 19476 8134 19488 8186
rect 19550 8134 19552 8186
rect 19390 8132 19414 8134
rect 19470 8132 19494 8134
rect 19550 8132 19574 8134
rect 19334 8112 19630 8132
rect 21272 7886 21300 8230
rect 21364 7954 21392 9318
rect 21352 7948 21404 7954
rect 21352 7890 21404 7896
rect 19236 7880 19288 7886
rect 19236 7822 19288 7828
rect 21076 7880 21128 7886
rect 21076 7822 21128 7828
rect 21260 7880 21312 7886
rect 21260 7822 21312 7828
rect 19052 7336 19104 7342
rect 19052 7278 19104 7284
rect 19248 7002 19276 7822
rect 20616 7744 20668 7750
rect 20616 7686 20668 7692
rect 19972 7200 20024 7206
rect 19972 7142 20024 7148
rect 20432 7200 20484 7206
rect 20432 7142 20484 7148
rect 19334 7100 19630 7120
rect 19390 7098 19414 7100
rect 19470 7098 19494 7100
rect 19550 7098 19574 7100
rect 19412 7046 19414 7098
rect 19476 7046 19488 7098
rect 19550 7046 19552 7098
rect 19390 7044 19414 7046
rect 19470 7044 19494 7046
rect 19550 7044 19574 7046
rect 19334 7024 19630 7044
rect 19236 6996 19288 7002
rect 19236 6938 19288 6944
rect 19144 6792 19196 6798
rect 19144 6734 19196 6740
rect 19052 6724 19104 6730
rect 19052 6666 19104 6672
rect 18960 6112 19012 6118
rect 18960 6054 19012 6060
rect 18774 3632 18830 3641
rect 18774 3567 18830 3576
rect 18972 3074 19000 6054
rect 19064 5914 19092 6666
rect 19156 6458 19184 6734
rect 19248 6458 19276 6938
rect 19694 6896 19750 6905
rect 19694 6831 19750 6840
rect 19144 6452 19196 6458
rect 19144 6394 19196 6400
rect 19236 6452 19288 6458
rect 19236 6394 19288 6400
rect 19234 6352 19290 6361
rect 19234 6287 19236 6296
rect 19288 6287 19290 6296
rect 19236 6258 19288 6264
rect 19334 6012 19630 6032
rect 19390 6010 19414 6012
rect 19470 6010 19494 6012
rect 19550 6010 19574 6012
rect 19412 5958 19414 6010
rect 19476 5958 19488 6010
rect 19550 5958 19552 6010
rect 19390 5956 19414 5958
rect 19470 5956 19494 5958
rect 19550 5956 19574 5958
rect 19334 5936 19630 5956
rect 19052 5908 19104 5914
rect 19052 5850 19104 5856
rect 19708 5778 19736 6831
rect 19984 6798 20012 7142
rect 19972 6792 20024 6798
rect 19972 6734 20024 6740
rect 19984 6458 20012 6734
rect 20444 6730 20472 7142
rect 20628 6934 20656 7686
rect 21088 7546 21116 7822
rect 21076 7540 21128 7546
rect 21076 7482 21128 7488
rect 21272 7478 21300 7822
rect 21260 7472 21312 7478
rect 21260 7414 21312 7420
rect 21364 7206 21392 7890
rect 21352 7200 21404 7206
rect 21352 7142 21404 7148
rect 20616 6928 20668 6934
rect 20616 6870 20668 6876
rect 20432 6724 20484 6730
rect 20432 6666 20484 6672
rect 19972 6452 20024 6458
rect 19972 6394 20024 6400
rect 19984 5914 20012 6394
rect 20444 6254 20472 6666
rect 20432 6248 20484 6254
rect 20432 6190 20484 6196
rect 19972 5908 20024 5914
rect 19972 5850 20024 5856
rect 21364 5778 21392 7142
rect 22284 7002 22312 9658
rect 23204 7562 23232 9959
rect 23940 8537 23968 10503
rect 24492 10169 24520 11494
rect 24478 10160 24534 10169
rect 24478 10095 24534 10104
rect 27238 10160 27294 10169
rect 27238 10095 27294 10104
rect 24001 9820 24297 9840
rect 24057 9818 24081 9820
rect 24137 9818 24161 9820
rect 24217 9818 24241 9820
rect 24079 9766 24081 9818
rect 24143 9766 24155 9818
rect 24217 9766 24219 9818
rect 24057 9764 24081 9766
rect 24137 9764 24161 9766
rect 24217 9764 24241 9766
rect 24001 9744 24297 9764
rect 24001 8732 24297 8752
rect 24057 8730 24081 8732
rect 24137 8730 24161 8732
rect 24217 8730 24241 8732
rect 24079 8678 24081 8730
rect 24143 8678 24155 8730
rect 24217 8678 24219 8730
rect 24057 8676 24081 8678
rect 24137 8676 24161 8678
rect 24217 8676 24241 8678
rect 24001 8656 24297 8676
rect 23926 8528 23982 8537
rect 23926 8463 23982 8472
rect 24478 7848 24534 7857
rect 24478 7783 24534 7792
rect 24001 7644 24297 7664
rect 24057 7642 24081 7644
rect 24137 7642 24161 7644
rect 24217 7642 24241 7644
rect 24079 7590 24081 7642
rect 24143 7590 24155 7642
rect 24217 7590 24219 7642
rect 24057 7588 24081 7590
rect 24137 7588 24161 7590
rect 24217 7588 24241 7590
rect 24001 7568 24297 7588
rect 23112 7546 23232 7562
rect 23100 7540 23232 7546
rect 23152 7534 23232 7540
rect 23100 7482 23152 7488
rect 22272 6996 22324 7002
rect 22272 6938 22324 6944
rect 21536 6860 21588 6866
rect 21536 6802 21588 6808
rect 21548 6118 21576 6802
rect 21536 6112 21588 6118
rect 21536 6054 21588 6060
rect 22180 6112 22232 6118
rect 22180 6054 22232 6060
rect 21534 5808 21590 5817
rect 19696 5772 19748 5778
rect 19696 5714 19748 5720
rect 20984 5772 21036 5778
rect 20984 5714 21036 5720
rect 21352 5772 21404 5778
rect 21534 5743 21590 5752
rect 21352 5714 21404 5720
rect 19708 5370 19736 5714
rect 19788 5568 19840 5574
rect 19788 5510 19840 5516
rect 19696 5364 19748 5370
rect 19696 5306 19748 5312
rect 19334 4924 19630 4944
rect 19390 4922 19414 4924
rect 19470 4922 19494 4924
rect 19550 4922 19574 4924
rect 19412 4870 19414 4922
rect 19476 4870 19488 4922
rect 19550 4870 19552 4922
rect 19390 4868 19414 4870
rect 19470 4868 19494 4870
rect 19550 4868 19574 4870
rect 19334 4848 19630 4868
rect 19334 3836 19630 3856
rect 19390 3834 19414 3836
rect 19470 3834 19494 3836
rect 19550 3834 19574 3836
rect 19412 3782 19414 3834
rect 19476 3782 19488 3834
rect 19550 3782 19552 3834
rect 19390 3780 19414 3782
rect 19470 3780 19494 3782
rect 19550 3780 19574 3782
rect 19334 3760 19630 3780
rect 18972 3046 19092 3074
rect 19064 480 19092 3046
rect 19334 2748 19630 2768
rect 19390 2746 19414 2748
rect 19470 2746 19494 2748
rect 19550 2746 19574 2748
rect 19412 2694 19414 2746
rect 19476 2694 19488 2746
rect 19550 2694 19552 2746
rect 19390 2692 19414 2694
rect 19470 2692 19494 2694
rect 19550 2692 19574 2694
rect 19334 2672 19630 2692
rect 19800 480 19828 5510
rect 20996 5030 21024 5714
rect 21444 5704 21496 5710
rect 21444 5646 21496 5652
rect 20156 5024 20208 5030
rect 20156 4966 20208 4972
rect 20984 5024 21036 5030
rect 20984 4966 21036 4972
rect 21260 5024 21312 5030
rect 21260 4966 21312 4972
rect 20168 4729 20196 4966
rect 20154 4720 20210 4729
rect 20154 4655 20210 4664
rect 20616 4684 20668 4690
rect 20616 4626 20668 4632
rect 20628 4282 20656 4626
rect 20616 4276 20668 4282
rect 20616 4218 20668 4224
rect 20996 3505 21024 4966
rect 21272 4690 21300 4966
rect 21456 4729 21484 5646
rect 21442 4720 21498 4729
rect 21260 4684 21312 4690
rect 21442 4655 21498 4664
rect 21260 4626 21312 4632
rect 21548 4146 21576 5743
rect 22192 5710 22220 6054
rect 22180 5704 22232 5710
rect 22180 5646 22232 5652
rect 21720 5568 21772 5574
rect 21720 5510 21772 5516
rect 21732 5234 21760 5510
rect 22192 5370 22220 5646
rect 22180 5364 22232 5370
rect 22180 5306 22232 5312
rect 22284 5234 22312 6938
rect 24001 6556 24297 6576
rect 24057 6554 24081 6556
rect 24137 6554 24161 6556
rect 24217 6554 24241 6556
rect 24079 6502 24081 6554
rect 24143 6502 24155 6554
rect 24217 6502 24219 6554
rect 24057 6500 24081 6502
rect 24137 6500 24161 6502
rect 24217 6500 24241 6502
rect 24001 6480 24297 6500
rect 24386 6488 24442 6497
rect 24386 6423 24442 6432
rect 24001 5468 24297 5488
rect 24057 5466 24081 5468
rect 24137 5466 24161 5468
rect 24217 5466 24241 5468
rect 24079 5414 24081 5466
rect 24143 5414 24155 5466
rect 24217 5414 24219 5466
rect 24057 5412 24081 5414
rect 24137 5412 24161 5414
rect 24217 5412 24241 5414
rect 24001 5392 24297 5412
rect 21720 5228 21772 5234
rect 21720 5170 21772 5176
rect 21812 5228 21864 5234
rect 21812 5170 21864 5176
rect 22272 5228 22324 5234
rect 22272 5170 22324 5176
rect 21628 5092 21680 5098
rect 21628 5034 21680 5040
rect 21640 4826 21668 5034
rect 21732 4826 21760 5170
rect 21628 4820 21680 4826
rect 21628 4762 21680 4768
rect 21720 4820 21772 4826
rect 21720 4762 21772 4768
rect 21824 4758 21852 5170
rect 24294 5128 24350 5137
rect 24294 5063 24350 5072
rect 21812 4752 21864 4758
rect 21812 4694 21864 4700
rect 24308 4690 24336 5063
rect 24400 4706 24428 6423
rect 24492 6361 24520 7783
rect 24478 6352 24534 6361
rect 24478 6287 24534 6296
rect 24296 4684 24348 4690
rect 24400 4678 24520 4706
rect 24296 4626 24348 4632
rect 24308 4570 24336 4626
rect 21812 4548 21864 4554
rect 24308 4542 24428 4570
rect 21812 4490 21864 4496
rect 21626 4176 21682 4185
rect 21536 4140 21588 4146
rect 21626 4111 21682 4120
rect 21536 4082 21588 4088
rect 21076 3936 21128 3942
rect 21076 3878 21128 3884
rect 20982 3496 21038 3505
rect 20982 3431 21038 3440
rect 20432 2304 20484 2310
rect 20432 2246 20484 2252
rect 20444 480 20472 2246
rect 21088 480 21116 3878
rect 21640 2650 21668 4111
rect 21824 4078 21852 4490
rect 23192 4480 23244 4486
rect 23192 4422 23244 4428
rect 21812 4072 21864 4078
rect 21812 4014 21864 4020
rect 22456 4004 22508 4010
rect 22456 3946 22508 3952
rect 21812 3188 21864 3194
rect 21812 3130 21864 3136
rect 21628 2644 21680 2650
rect 21628 2586 21680 2592
rect 21824 480 21852 3130
rect 22468 480 22496 3946
rect 23204 3210 23232 4422
rect 24001 4380 24297 4400
rect 24057 4378 24081 4380
rect 24137 4378 24161 4380
rect 24217 4378 24241 4380
rect 24079 4326 24081 4378
rect 24143 4326 24155 4378
rect 24217 4326 24219 4378
rect 24057 4324 24081 4326
rect 24137 4324 24161 4326
rect 24217 4324 24241 4326
rect 24001 4304 24297 4324
rect 24400 4282 24428 4542
rect 24388 4276 24440 4282
rect 24388 4218 24440 4224
rect 24492 4185 24520 4678
rect 24478 4176 24534 4185
rect 24478 4111 24534 4120
rect 23928 4072 23980 4078
rect 23928 4014 23980 4020
rect 23652 3392 23704 3398
rect 23652 3334 23704 3340
rect 23112 3194 23232 3210
rect 23100 3188 23232 3194
rect 23152 3182 23232 3188
rect 23100 3130 23152 3136
rect 23664 3097 23692 3334
rect 23650 3088 23706 3097
rect 23650 3023 23706 3032
rect 23664 2990 23692 3023
rect 23652 2984 23704 2990
rect 22730 2952 22786 2961
rect 23652 2926 23704 2932
rect 22730 2887 22786 2896
rect 22744 2650 22772 2887
rect 23836 2848 23888 2854
rect 23836 2790 23888 2796
rect 22732 2644 22784 2650
rect 22732 2586 22784 2592
rect 23284 2440 23336 2446
rect 23284 2382 23336 2388
rect 23192 2304 23244 2310
rect 23192 2246 23244 2252
rect 23204 480 23232 2246
rect 23296 1057 23324 2382
rect 23282 1048 23338 1057
rect 23282 983 23338 992
rect 23848 480 23876 2790
rect 6 0 62 480
rect 650 0 706 480
rect 1294 0 1350 480
rect 2030 0 2086 480
rect 2674 0 2730 480
rect 3410 0 3466 480
rect 4054 0 4110 480
rect 4698 0 4754 480
rect 5434 0 5490 480
rect 6078 0 6134 480
rect 6814 0 6870 480
rect 7458 0 7514 480
rect 8102 0 8158 480
rect 8838 0 8894 480
rect 9482 0 9538 480
rect 10218 0 10274 480
rect 10862 0 10918 480
rect 11598 0 11654 480
rect 12242 0 12298 480
rect 12886 0 12942 480
rect 13622 0 13678 480
rect 14266 0 14322 480
rect 15002 0 15058 480
rect 15646 0 15702 480
rect 16290 0 16346 480
rect 17026 0 17082 480
rect 17670 0 17726 480
rect 18406 0 18462 480
rect 19050 0 19106 480
rect 19786 0 19842 480
rect 20430 0 20486 480
rect 21074 0 21130 480
rect 21810 0 21866 480
rect 22454 0 22510 480
rect 23190 0 23246 480
rect 23834 0 23890 480
rect 23940 377 23968 4014
rect 24480 3936 24532 3942
rect 24480 3878 24532 3884
rect 24388 3596 24440 3602
rect 24388 3538 24440 3544
rect 24001 3292 24297 3312
rect 24057 3290 24081 3292
rect 24137 3290 24161 3292
rect 24217 3290 24241 3292
rect 24079 3238 24081 3290
rect 24143 3238 24155 3290
rect 24217 3238 24219 3290
rect 24057 3236 24081 3238
rect 24137 3236 24161 3238
rect 24217 3236 24241 3238
rect 24001 3216 24297 3236
rect 24400 3194 24428 3538
rect 24492 3369 24520 3878
rect 25216 3392 25268 3398
rect 24478 3360 24534 3369
rect 25216 3334 25268 3340
rect 26594 3360 26650 3369
rect 24478 3295 24534 3304
rect 24478 3224 24534 3233
rect 24388 3188 24440 3194
rect 24478 3159 24534 3168
rect 24388 3130 24440 3136
rect 24400 3074 24428 3130
rect 24308 3046 24428 3074
rect 24308 2530 24336 3046
rect 24492 2938 24520 3159
rect 24400 2910 24520 2938
rect 24400 2650 24428 2910
rect 24480 2848 24532 2854
rect 24480 2790 24532 2796
rect 24388 2644 24440 2650
rect 24388 2586 24440 2592
rect 24308 2502 24428 2530
rect 24001 2204 24297 2224
rect 24057 2202 24081 2204
rect 24137 2202 24161 2204
rect 24217 2202 24241 2204
rect 24079 2150 24081 2202
rect 24143 2150 24155 2202
rect 24217 2150 24219 2202
rect 24057 2148 24081 2150
rect 24137 2148 24161 2150
rect 24217 2148 24241 2150
rect 24001 2128 24297 2148
rect 24400 1737 24428 2502
rect 24386 1728 24442 1737
rect 24386 1663 24442 1672
rect 24492 480 24520 2790
rect 25228 480 25256 3334
rect 26594 3295 26650 3304
rect 25858 2952 25914 2961
rect 25858 2887 25914 2896
rect 25308 2848 25360 2854
rect 25306 2816 25308 2825
rect 25360 2816 25362 2825
rect 25306 2751 25362 2760
rect 25872 480 25900 2887
rect 26608 480 26636 3295
rect 27252 480 27280 10095
rect 23926 368 23982 377
rect 23926 303 23982 312
rect 24478 0 24534 480
rect 25214 0 25270 480
rect 25858 0 25914 480
rect 26594 0 26650 480
rect 27238 0 27294 480
<< via2 >>
rect 2030 23044 2086 23080
rect 2030 23024 2032 23044
rect 2032 23024 2084 23044
rect 2084 23024 2086 23044
rect 650 3984 706 4040
rect 6 3440 62 3496
rect 2674 22480 2730 22536
rect 4054 22344 4110 22400
rect 3962 21956 4018 21992
rect 3962 21936 3964 21956
rect 3964 21936 4016 21956
rect 4016 21936 4018 21956
rect 1294 3032 1350 3088
rect 10001 25594 10057 25596
rect 10081 25594 10137 25596
rect 10161 25594 10217 25596
rect 10241 25594 10297 25596
rect 10001 25542 10027 25594
rect 10027 25542 10057 25594
rect 10081 25542 10091 25594
rect 10091 25542 10137 25594
rect 10161 25542 10207 25594
rect 10207 25542 10217 25594
rect 10241 25542 10271 25594
rect 10271 25542 10297 25594
rect 10001 25540 10057 25542
rect 10081 25540 10137 25542
rect 10161 25540 10217 25542
rect 10241 25540 10297 25542
rect 5334 25050 5390 25052
rect 5414 25050 5470 25052
rect 5494 25050 5550 25052
rect 5574 25050 5630 25052
rect 5334 24998 5360 25050
rect 5360 24998 5390 25050
rect 5414 24998 5424 25050
rect 5424 24998 5470 25050
rect 5494 24998 5540 25050
rect 5540 24998 5550 25050
rect 5574 24998 5604 25050
rect 5604 24998 5630 25050
rect 5334 24996 5390 24998
rect 5414 24996 5470 24998
rect 5494 24996 5550 24998
rect 5574 24996 5630 24998
rect 10001 24506 10057 24508
rect 10081 24506 10137 24508
rect 10161 24506 10217 24508
rect 10241 24506 10297 24508
rect 10001 24454 10027 24506
rect 10027 24454 10057 24506
rect 10081 24454 10091 24506
rect 10091 24454 10137 24506
rect 10161 24454 10207 24506
rect 10207 24454 10217 24506
rect 10241 24454 10271 24506
rect 10271 24454 10297 24506
rect 10001 24452 10057 24454
rect 10081 24452 10137 24454
rect 10161 24452 10217 24454
rect 10241 24452 10297 24454
rect 5334 23962 5390 23964
rect 5414 23962 5470 23964
rect 5494 23962 5550 23964
rect 5574 23962 5630 23964
rect 5334 23910 5360 23962
rect 5360 23910 5390 23962
rect 5414 23910 5424 23962
rect 5424 23910 5470 23962
rect 5494 23910 5540 23962
rect 5540 23910 5550 23962
rect 5574 23910 5604 23962
rect 5604 23910 5630 23962
rect 5334 23908 5390 23910
rect 5414 23908 5470 23910
rect 5494 23908 5550 23910
rect 5574 23908 5630 23910
rect 10001 23418 10057 23420
rect 10081 23418 10137 23420
rect 10161 23418 10217 23420
rect 10241 23418 10297 23420
rect 10001 23366 10027 23418
rect 10027 23366 10057 23418
rect 10081 23366 10091 23418
rect 10091 23366 10137 23418
rect 10161 23366 10207 23418
rect 10207 23366 10217 23418
rect 10241 23366 10271 23418
rect 10271 23366 10297 23418
rect 10001 23364 10057 23366
rect 10081 23364 10137 23366
rect 10161 23364 10217 23366
rect 10241 23364 10297 23366
rect 5710 22888 5766 22944
rect 5334 22874 5390 22876
rect 5414 22874 5470 22876
rect 5494 22874 5550 22876
rect 5574 22874 5630 22876
rect 5334 22822 5360 22874
rect 5360 22822 5390 22874
rect 5414 22822 5424 22874
rect 5424 22822 5470 22874
rect 5494 22822 5540 22874
rect 5540 22822 5550 22874
rect 5574 22822 5604 22874
rect 5604 22822 5630 22874
rect 5334 22820 5390 22822
rect 5414 22820 5470 22822
rect 5494 22820 5550 22822
rect 5574 22820 5630 22822
rect 5710 22344 5766 22400
rect 10001 22330 10057 22332
rect 10081 22330 10137 22332
rect 10161 22330 10217 22332
rect 10241 22330 10297 22332
rect 10001 22278 10027 22330
rect 10027 22278 10057 22330
rect 10081 22278 10091 22330
rect 10091 22278 10137 22330
rect 10161 22278 10207 22330
rect 10207 22278 10217 22330
rect 10241 22278 10271 22330
rect 10271 22278 10297 22330
rect 10001 22276 10057 22278
rect 10081 22276 10137 22278
rect 10161 22276 10217 22278
rect 10241 22276 10297 22278
rect 5334 21786 5390 21788
rect 5414 21786 5470 21788
rect 5494 21786 5550 21788
rect 5574 21786 5630 21788
rect 5334 21734 5360 21786
rect 5360 21734 5390 21786
rect 5414 21734 5424 21786
rect 5424 21734 5470 21786
rect 5494 21734 5540 21786
rect 5540 21734 5550 21786
rect 5574 21734 5604 21786
rect 5604 21734 5630 21786
rect 5334 21732 5390 21734
rect 5414 21732 5470 21734
rect 5494 21732 5550 21734
rect 5574 21732 5630 21734
rect 10001 21242 10057 21244
rect 10081 21242 10137 21244
rect 10161 21242 10217 21244
rect 10241 21242 10297 21244
rect 10001 21190 10027 21242
rect 10027 21190 10057 21242
rect 10081 21190 10091 21242
rect 10091 21190 10137 21242
rect 10161 21190 10207 21242
rect 10207 21190 10217 21242
rect 10241 21190 10271 21242
rect 10271 21190 10297 21242
rect 10001 21188 10057 21190
rect 10081 21188 10137 21190
rect 10161 21188 10217 21190
rect 10241 21188 10297 21190
rect 5710 20848 5766 20904
rect 5334 20698 5390 20700
rect 5414 20698 5470 20700
rect 5494 20698 5550 20700
rect 5574 20698 5630 20700
rect 5334 20646 5360 20698
rect 5360 20646 5390 20698
rect 5414 20646 5424 20698
rect 5424 20646 5470 20698
rect 5494 20646 5540 20698
rect 5540 20646 5550 20698
rect 5574 20646 5604 20698
rect 5604 20646 5630 20698
rect 5334 20644 5390 20646
rect 5414 20644 5470 20646
rect 5494 20644 5550 20646
rect 5574 20644 5630 20646
rect 10001 20154 10057 20156
rect 10081 20154 10137 20156
rect 10161 20154 10217 20156
rect 10241 20154 10297 20156
rect 10001 20102 10027 20154
rect 10027 20102 10057 20154
rect 10081 20102 10091 20154
rect 10091 20102 10137 20154
rect 10161 20102 10207 20154
rect 10207 20102 10217 20154
rect 10241 20102 10271 20154
rect 10271 20102 10297 20154
rect 10001 20100 10057 20102
rect 10081 20100 10137 20102
rect 10161 20100 10217 20102
rect 10241 20100 10297 20102
rect 6722 19896 6778 19952
rect 5334 19610 5390 19612
rect 5414 19610 5470 19612
rect 5494 19610 5550 19612
rect 5574 19610 5630 19612
rect 5334 19558 5360 19610
rect 5360 19558 5390 19610
rect 5414 19558 5424 19610
rect 5424 19558 5470 19610
rect 5494 19558 5540 19610
rect 5540 19558 5550 19610
rect 5574 19558 5604 19610
rect 5604 19558 5630 19610
rect 5334 19556 5390 19558
rect 5414 19556 5470 19558
rect 5494 19556 5550 19558
rect 5574 19556 5630 19558
rect 4330 13776 4386 13832
rect 4698 3576 4754 3632
rect 5334 18522 5390 18524
rect 5414 18522 5470 18524
rect 5494 18522 5550 18524
rect 5574 18522 5630 18524
rect 5334 18470 5360 18522
rect 5360 18470 5390 18522
rect 5414 18470 5424 18522
rect 5424 18470 5470 18522
rect 5494 18470 5540 18522
rect 5540 18470 5550 18522
rect 5574 18470 5604 18522
rect 5604 18470 5630 18522
rect 5334 18468 5390 18470
rect 5414 18468 5470 18470
rect 5494 18468 5550 18470
rect 5574 18468 5630 18470
rect 5334 17434 5390 17436
rect 5414 17434 5470 17436
rect 5494 17434 5550 17436
rect 5574 17434 5630 17436
rect 5334 17382 5360 17434
rect 5360 17382 5390 17434
rect 5414 17382 5424 17434
rect 5424 17382 5470 17434
rect 5494 17382 5540 17434
rect 5540 17382 5550 17434
rect 5574 17382 5604 17434
rect 5604 17382 5630 17434
rect 5334 17380 5390 17382
rect 5414 17380 5470 17382
rect 5494 17380 5550 17382
rect 5574 17380 5630 17382
rect 5334 16346 5390 16348
rect 5414 16346 5470 16348
rect 5494 16346 5550 16348
rect 5574 16346 5630 16348
rect 5334 16294 5360 16346
rect 5360 16294 5390 16346
rect 5414 16294 5424 16346
rect 5424 16294 5470 16346
rect 5494 16294 5540 16346
rect 5540 16294 5550 16346
rect 5574 16294 5604 16346
rect 5604 16294 5630 16346
rect 5334 16292 5390 16294
rect 5414 16292 5470 16294
rect 5494 16292 5550 16294
rect 5574 16292 5630 16294
rect 5334 15258 5390 15260
rect 5414 15258 5470 15260
rect 5494 15258 5550 15260
rect 5574 15258 5630 15260
rect 5334 15206 5360 15258
rect 5360 15206 5390 15258
rect 5414 15206 5424 15258
rect 5424 15206 5470 15258
rect 5494 15206 5540 15258
rect 5540 15206 5550 15258
rect 5574 15206 5604 15258
rect 5604 15206 5630 15258
rect 5334 15204 5390 15206
rect 5414 15204 5470 15206
rect 5494 15204 5550 15206
rect 5574 15204 5630 15206
rect 5334 14170 5390 14172
rect 5414 14170 5470 14172
rect 5494 14170 5550 14172
rect 5574 14170 5630 14172
rect 5334 14118 5360 14170
rect 5360 14118 5390 14170
rect 5414 14118 5424 14170
rect 5424 14118 5470 14170
rect 5494 14118 5540 14170
rect 5540 14118 5550 14170
rect 5574 14118 5604 14170
rect 5604 14118 5630 14170
rect 5334 14116 5390 14118
rect 5414 14116 5470 14118
rect 5494 14116 5550 14118
rect 5574 14116 5630 14118
rect 5334 13082 5390 13084
rect 5414 13082 5470 13084
rect 5494 13082 5550 13084
rect 5574 13082 5630 13084
rect 5334 13030 5360 13082
rect 5360 13030 5390 13082
rect 5414 13030 5424 13082
rect 5424 13030 5470 13082
rect 5494 13030 5540 13082
rect 5540 13030 5550 13082
rect 5574 13030 5604 13082
rect 5604 13030 5630 13082
rect 5334 13028 5390 13030
rect 5414 13028 5470 13030
rect 5494 13028 5550 13030
rect 5574 13028 5630 13030
rect 5334 11994 5390 11996
rect 5414 11994 5470 11996
rect 5494 11994 5550 11996
rect 5574 11994 5630 11996
rect 5334 11942 5360 11994
rect 5360 11942 5390 11994
rect 5414 11942 5424 11994
rect 5424 11942 5470 11994
rect 5494 11942 5540 11994
rect 5540 11942 5550 11994
rect 5574 11942 5604 11994
rect 5604 11942 5630 11994
rect 5334 11940 5390 11942
rect 5414 11940 5470 11942
rect 5494 11940 5550 11942
rect 5574 11940 5630 11942
rect 5334 10906 5390 10908
rect 5414 10906 5470 10908
rect 5494 10906 5550 10908
rect 5574 10906 5630 10908
rect 5334 10854 5360 10906
rect 5360 10854 5390 10906
rect 5414 10854 5424 10906
rect 5424 10854 5470 10906
rect 5494 10854 5540 10906
rect 5540 10854 5550 10906
rect 5574 10854 5604 10906
rect 5604 10854 5630 10906
rect 5334 10852 5390 10854
rect 5414 10852 5470 10854
rect 5494 10852 5550 10854
rect 5574 10852 5630 10854
rect 5334 9818 5390 9820
rect 5414 9818 5470 9820
rect 5494 9818 5550 9820
rect 5574 9818 5630 9820
rect 5334 9766 5360 9818
rect 5360 9766 5390 9818
rect 5414 9766 5424 9818
rect 5424 9766 5470 9818
rect 5494 9766 5540 9818
rect 5540 9766 5550 9818
rect 5574 9766 5604 9818
rect 5604 9766 5630 9818
rect 5334 9764 5390 9766
rect 5414 9764 5470 9766
rect 5494 9764 5550 9766
rect 5574 9764 5630 9766
rect 5334 8730 5390 8732
rect 5414 8730 5470 8732
rect 5494 8730 5550 8732
rect 5574 8730 5630 8732
rect 5334 8678 5360 8730
rect 5360 8678 5390 8730
rect 5414 8678 5424 8730
rect 5424 8678 5470 8730
rect 5494 8678 5540 8730
rect 5540 8678 5550 8730
rect 5574 8678 5604 8730
rect 5604 8678 5630 8730
rect 5334 8676 5390 8678
rect 5414 8676 5470 8678
rect 5494 8676 5550 8678
rect 5574 8676 5630 8678
rect 5334 7642 5390 7644
rect 5414 7642 5470 7644
rect 5494 7642 5550 7644
rect 5574 7642 5630 7644
rect 5334 7590 5360 7642
rect 5360 7590 5390 7642
rect 5414 7590 5424 7642
rect 5424 7590 5470 7642
rect 5494 7590 5540 7642
rect 5540 7590 5550 7642
rect 5574 7590 5604 7642
rect 5604 7590 5630 7642
rect 5334 7588 5390 7590
rect 5414 7588 5470 7590
rect 5494 7588 5550 7590
rect 5574 7588 5630 7590
rect 5334 6554 5390 6556
rect 5414 6554 5470 6556
rect 5494 6554 5550 6556
rect 5574 6554 5630 6556
rect 5334 6502 5360 6554
rect 5360 6502 5390 6554
rect 5414 6502 5424 6554
rect 5424 6502 5470 6554
rect 5494 6502 5540 6554
rect 5540 6502 5550 6554
rect 5574 6502 5604 6554
rect 5604 6502 5630 6554
rect 5334 6500 5390 6502
rect 5414 6500 5470 6502
rect 5494 6500 5550 6502
rect 5574 6500 5630 6502
rect 5334 5466 5390 5468
rect 5414 5466 5470 5468
rect 5494 5466 5550 5468
rect 5574 5466 5630 5468
rect 5334 5414 5360 5466
rect 5360 5414 5390 5466
rect 5414 5414 5424 5466
rect 5424 5414 5470 5466
rect 5494 5414 5540 5466
rect 5540 5414 5550 5466
rect 5574 5414 5604 5466
rect 5604 5414 5630 5466
rect 5334 5412 5390 5414
rect 5414 5412 5470 5414
rect 5494 5412 5550 5414
rect 5574 5412 5630 5414
rect 5334 4378 5390 4380
rect 5414 4378 5470 4380
rect 5494 4378 5550 4380
rect 5574 4378 5630 4380
rect 5334 4326 5360 4378
rect 5360 4326 5390 4378
rect 5414 4326 5424 4378
rect 5424 4326 5470 4378
rect 5494 4326 5540 4378
rect 5540 4326 5550 4378
rect 5574 4326 5604 4378
rect 5604 4326 5630 4378
rect 5334 4324 5390 4326
rect 5414 4324 5470 4326
rect 5494 4324 5550 4326
rect 5574 4324 5630 4326
rect 6814 19352 6870 19408
rect 10001 19066 10057 19068
rect 10081 19066 10137 19068
rect 10161 19066 10217 19068
rect 10241 19066 10297 19068
rect 10001 19014 10027 19066
rect 10027 19014 10057 19066
rect 10081 19014 10091 19066
rect 10091 19014 10137 19066
rect 10161 19014 10207 19066
rect 10207 19014 10217 19066
rect 10241 19014 10271 19066
rect 10271 19014 10297 19066
rect 10001 19012 10057 19014
rect 10081 19012 10137 19014
rect 10161 19012 10217 19014
rect 10241 19012 10297 19014
rect 5334 3290 5390 3292
rect 5414 3290 5470 3292
rect 5494 3290 5550 3292
rect 5574 3290 5630 3292
rect 5334 3238 5360 3290
rect 5360 3238 5390 3290
rect 5414 3238 5424 3290
rect 5424 3238 5470 3290
rect 5494 3238 5540 3290
rect 5540 3238 5550 3290
rect 5574 3238 5604 3290
rect 5604 3238 5630 3290
rect 5334 3236 5390 3238
rect 5414 3236 5470 3238
rect 5494 3236 5550 3238
rect 5574 3236 5630 3238
rect 5334 2202 5390 2204
rect 5414 2202 5470 2204
rect 5494 2202 5550 2204
rect 5574 2202 5630 2204
rect 5334 2150 5360 2202
rect 5360 2150 5390 2202
rect 5414 2150 5424 2202
rect 5424 2150 5470 2202
rect 5494 2150 5540 2202
rect 5540 2150 5550 2202
rect 5574 2150 5604 2202
rect 5604 2150 5630 2202
rect 5334 2148 5390 2150
rect 5414 2148 5470 2150
rect 5494 2148 5550 2150
rect 5574 2148 5630 2150
rect 10001 17978 10057 17980
rect 10081 17978 10137 17980
rect 10161 17978 10217 17980
rect 10241 17978 10297 17980
rect 10001 17926 10027 17978
rect 10027 17926 10057 17978
rect 10081 17926 10091 17978
rect 10091 17926 10137 17978
rect 10161 17926 10207 17978
rect 10207 17926 10217 17978
rect 10241 17926 10271 17978
rect 10271 17926 10297 17978
rect 10001 17924 10057 17926
rect 10081 17924 10137 17926
rect 10161 17924 10217 17926
rect 10241 17924 10297 17926
rect 7458 17604 7514 17640
rect 7458 17584 7460 17604
rect 7460 17584 7512 17604
rect 7512 17584 7514 17604
rect 9574 17176 9630 17232
rect 8102 17040 8158 17096
rect 8010 15136 8066 15192
rect 10001 16890 10057 16892
rect 10081 16890 10137 16892
rect 10161 16890 10217 16892
rect 10241 16890 10297 16892
rect 10001 16838 10027 16890
rect 10027 16838 10057 16890
rect 10081 16838 10091 16890
rect 10091 16838 10137 16890
rect 10161 16838 10207 16890
rect 10207 16838 10217 16890
rect 10241 16838 10271 16890
rect 10271 16838 10297 16890
rect 10001 16836 10057 16838
rect 10081 16836 10137 16838
rect 10161 16836 10217 16838
rect 10241 16836 10297 16838
rect 9482 16632 9538 16688
rect 10001 15802 10057 15804
rect 10081 15802 10137 15804
rect 10161 15802 10217 15804
rect 10241 15802 10297 15804
rect 10001 15750 10027 15802
rect 10027 15750 10057 15802
rect 10081 15750 10091 15802
rect 10091 15750 10137 15802
rect 10161 15750 10207 15802
rect 10207 15750 10217 15802
rect 10241 15750 10271 15802
rect 10271 15750 10297 15802
rect 10001 15748 10057 15750
rect 10081 15748 10137 15750
rect 10161 15748 10217 15750
rect 10241 15748 10297 15750
rect 9850 15136 9906 15192
rect 10001 14714 10057 14716
rect 10081 14714 10137 14716
rect 10161 14714 10217 14716
rect 10241 14714 10297 14716
rect 10001 14662 10027 14714
rect 10027 14662 10057 14714
rect 10081 14662 10091 14714
rect 10091 14662 10137 14714
rect 10161 14662 10207 14714
rect 10207 14662 10217 14714
rect 10241 14662 10271 14714
rect 10271 14662 10297 14714
rect 10001 14660 10057 14662
rect 10081 14660 10137 14662
rect 10161 14660 10217 14662
rect 10241 14660 10297 14662
rect 10001 13626 10057 13628
rect 10081 13626 10137 13628
rect 10161 13626 10217 13628
rect 10241 13626 10297 13628
rect 10001 13574 10027 13626
rect 10027 13574 10057 13626
rect 10081 13574 10091 13626
rect 10091 13574 10137 13626
rect 10161 13574 10207 13626
rect 10207 13574 10217 13626
rect 10241 13574 10271 13626
rect 10271 13574 10297 13626
rect 10001 13572 10057 13574
rect 10081 13572 10137 13574
rect 10161 13572 10217 13574
rect 10241 13572 10297 13574
rect 10001 12538 10057 12540
rect 10081 12538 10137 12540
rect 10161 12538 10217 12540
rect 10241 12538 10297 12540
rect 10001 12486 10027 12538
rect 10027 12486 10057 12538
rect 10081 12486 10091 12538
rect 10091 12486 10137 12538
rect 10161 12486 10207 12538
rect 10207 12486 10217 12538
rect 10241 12486 10271 12538
rect 10271 12486 10297 12538
rect 10001 12484 10057 12486
rect 10081 12484 10137 12486
rect 10161 12484 10217 12486
rect 10241 12484 10297 12486
rect 10001 11450 10057 11452
rect 10081 11450 10137 11452
rect 10161 11450 10217 11452
rect 10241 11450 10297 11452
rect 10001 11398 10027 11450
rect 10027 11398 10057 11450
rect 10081 11398 10091 11450
rect 10091 11398 10137 11450
rect 10161 11398 10207 11450
rect 10207 11398 10217 11450
rect 10241 11398 10271 11450
rect 10271 11398 10297 11450
rect 10001 11396 10057 11398
rect 10081 11396 10137 11398
rect 10161 11396 10217 11398
rect 10241 11396 10297 11398
rect 9390 11192 9446 11248
rect 10001 10362 10057 10364
rect 10081 10362 10137 10364
rect 10161 10362 10217 10364
rect 10241 10362 10297 10364
rect 10001 10310 10027 10362
rect 10027 10310 10057 10362
rect 10081 10310 10091 10362
rect 10091 10310 10137 10362
rect 10161 10310 10207 10362
rect 10207 10310 10217 10362
rect 10241 10310 10271 10362
rect 10271 10310 10297 10362
rect 10001 10308 10057 10310
rect 10081 10308 10137 10310
rect 10161 10308 10217 10310
rect 10241 10308 10297 10310
rect 10001 9274 10057 9276
rect 10081 9274 10137 9276
rect 10161 9274 10217 9276
rect 10241 9274 10297 9276
rect 10001 9222 10027 9274
rect 10027 9222 10057 9274
rect 10081 9222 10091 9274
rect 10091 9222 10137 9274
rect 10161 9222 10207 9274
rect 10207 9222 10217 9274
rect 10241 9222 10271 9274
rect 10271 9222 10297 9274
rect 10001 9220 10057 9222
rect 10081 9220 10137 9222
rect 10161 9220 10217 9222
rect 10241 9220 10297 9222
rect 10001 8186 10057 8188
rect 10081 8186 10137 8188
rect 10161 8186 10217 8188
rect 10241 8186 10297 8188
rect 10001 8134 10027 8186
rect 10027 8134 10057 8186
rect 10081 8134 10091 8186
rect 10091 8134 10137 8186
rect 10161 8134 10207 8186
rect 10207 8134 10217 8186
rect 10241 8134 10271 8186
rect 10271 8134 10297 8186
rect 10001 8132 10057 8134
rect 10081 8132 10137 8134
rect 10161 8132 10217 8134
rect 10241 8132 10297 8134
rect 10001 7098 10057 7100
rect 10081 7098 10137 7100
rect 10161 7098 10217 7100
rect 10241 7098 10297 7100
rect 10001 7046 10027 7098
rect 10027 7046 10057 7098
rect 10081 7046 10091 7098
rect 10091 7046 10137 7098
rect 10161 7046 10207 7098
rect 10207 7046 10217 7098
rect 10241 7046 10271 7098
rect 10271 7046 10297 7098
rect 10001 7044 10057 7046
rect 10081 7044 10137 7046
rect 10161 7044 10217 7046
rect 10241 7044 10297 7046
rect 10001 6010 10057 6012
rect 10081 6010 10137 6012
rect 10161 6010 10217 6012
rect 10241 6010 10297 6012
rect 10001 5958 10027 6010
rect 10027 5958 10057 6010
rect 10081 5958 10091 6010
rect 10091 5958 10137 6010
rect 10161 5958 10207 6010
rect 10207 5958 10217 6010
rect 10241 5958 10271 6010
rect 10271 5958 10297 6010
rect 10001 5956 10057 5958
rect 10081 5956 10137 5958
rect 10161 5956 10217 5958
rect 10241 5956 10297 5958
rect 10001 4922 10057 4924
rect 10081 4922 10137 4924
rect 10161 4922 10217 4924
rect 10241 4922 10297 4924
rect 10001 4870 10027 4922
rect 10027 4870 10057 4922
rect 10081 4870 10091 4922
rect 10091 4870 10137 4922
rect 10161 4870 10207 4922
rect 10207 4870 10217 4922
rect 10241 4870 10271 4922
rect 10271 4870 10297 4922
rect 10001 4868 10057 4870
rect 10081 4868 10137 4870
rect 10161 4868 10217 4870
rect 10241 4868 10297 4870
rect 10001 3834 10057 3836
rect 10081 3834 10137 3836
rect 10161 3834 10217 3836
rect 10241 3834 10297 3836
rect 10001 3782 10027 3834
rect 10027 3782 10057 3834
rect 10081 3782 10091 3834
rect 10091 3782 10137 3834
rect 10161 3782 10207 3834
rect 10207 3782 10217 3834
rect 10241 3782 10271 3834
rect 10271 3782 10297 3834
rect 10001 3780 10057 3782
rect 10081 3780 10137 3782
rect 10161 3780 10217 3782
rect 10241 3780 10297 3782
rect 10862 15408 10918 15464
rect 10770 11464 10826 11520
rect 11046 3984 11102 4040
rect 14668 25050 14724 25052
rect 14748 25050 14804 25052
rect 14828 25050 14884 25052
rect 14908 25050 14964 25052
rect 14668 24998 14694 25050
rect 14694 24998 14724 25050
rect 14748 24998 14758 25050
rect 14758 24998 14804 25050
rect 14828 24998 14874 25050
rect 14874 24998 14884 25050
rect 14908 24998 14938 25050
rect 14938 24998 14964 25050
rect 14668 24996 14724 24998
rect 14748 24996 14804 24998
rect 14828 24996 14884 24998
rect 14908 24996 14964 24998
rect 14668 23962 14724 23964
rect 14748 23962 14804 23964
rect 14828 23962 14884 23964
rect 14908 23962 14964 23964
rect 14668 23910 14694 23962
rect 14694 23910 14724 23962
rect 14748 23910 14758 23962
rect 14758 23910 14804 23962
rect 14828 23910 14874 23962
rect 14874 23910 14884 23962
rect 14908 23910 14938 23962
rect 14938 23910 14964 23962
rect 14668 23908 14724 23910
rect 14748 23908 14804 23910
rect 14828 23908 14884 23910
rect 14908 23908 14964 23910
rect 14450 22924 14452 22944
rect 14452 22924 14504 22944
rect 14504 22924 14506 22944
rect 14450 22888 14506 22924
rect 15094 22924 15096 22944
rect 15096 22924 15148 22944
rect 15148 22924 15150 22944
rect 15094 22888 15150 22924
rect 14668 22874 14724 22876
rect 14748 22874 14804 22876
rect 14828 22874 14884 22876
rect 14908 22874 14964 22876
rect 14668 22822 14694 22874
rect 14694 22822 14724 22874
rect 14748 22822 14758 22874
rect 14758 22822 14804 22874
rect 14828 22822 14874 22874
rect 14874 22822 14884 22874
rect 14908 22822 14938 22874
rect 14938 22822 14964 22874
rect 14668 22820 14724 22822
rect 14748 22820 14804 22822
rect 14828 22820 14884 22822
rect 14908 22820 14964 22822
rect 14668 21786 14724 21788
rect 14748 21786 14804 21788
rect 14828 21786 14884 21788
rect 14908 21786 14964 21788
rect 14668 21734 14694 21786
rect 14694 21734 14724 21786
rect 14748 21734 14758 21786
rect 14758 21734 14804 21786
rect 14828 21734 14874 21786
rect 14874 21734 14884 21786
rect 14908 21734 14938 21786
rect 14938 21734 14964 21786
rect 14668 21732 14724 21734
rect 14748 21732 14804 21734
rect 14828 21732 14884 21734
rect 14908 21732 14964 21734
rect 14174 20984 14230 21040
rect 14668 20698 14724 20700
rect 14748 20698 14804 20700
rect 14828 20698 14884 20700
rect 14908 20698 14964 20700
rect 14668 20646 14694 20698
rect 14694 20646 14724 20698
rect 14748 20646 14758 20698
rect 14758 20646 14804 20698
rect 14828 20646 14874 20698
rect 14874 20646 14884 20698
rect 14908 20646 14938 20698
rect 14938 20646 14964 20698
rect 14668 20644 14724 20646
rect 14748 20644 14804 20646
rect 14828 20644 14884 20646
rect 14908 20644 14964 20646
rect 14174 20576 14230 20632
rect 14668 19610 14724 19612
rect 14748 19610 14804 19612
rect 14828 19610 14884 19612
rect 14908 19610 14964 19612
rect 14668 19558 14694 19610
rect 14694 19558 14724 19610
rect 14748 19558 14758 19610
rect 14758 19558 14804 19610
rect 14828 19558 14874 19610
rect 14874 19558 14884 19610
rect 14908 19558 14938 19610
rect 14938 19558 14964 19610
rect 14668 19556 14724 19558
rect 14748 19556 14804 19558
rect 14828 19556 14884 19558
rect 14908 19556 14964 19558
rect 14668 18522 14724 18524
rect 14748 18522 14804 18524
rect 14828 18522 14884 18524
rect 14908 18522 14964 18524
rect 14668 18470 14694 18522
rect 14694 18470 14724 18522
rect 14748 18470 14758 18522
rect 14758 18470 14804 18522
rect 14828 18470 14874 18522
rect 14874 18470 14884 18522
rect 14908 18470 14938 18522
rect 14938 18470 14964 18522
rect 14668 18468 14724 18470
rect 14748 18468 14804 18470
rect 14828 18468 14884 18470
rect 14908 18468 14964 18470
rect 14668 17434 14724 17436
rect 14748 17434 14804 17436
rect 14828 17434 14884 17436
rect 14908 17434 14964 17436
rect 14668 17382 14694 17434
rect 14694 17382 14724 17434
rect 14748 17382 14758 17434
rect 14758 17382 14804 17434
rect 14828 17382 14874 17434
rect 14874 17382 14884 17434
rect 14908 17382 14938 17434
rect 14938 17382 14964 17434
rect 14668 17380 14724 17382
rect 14748 17380 14804 17382
rect 14828 17380 14884 17382
rect 14908 17380 14964 17382
rect 16750 17312 16806 17368
rect 19334 25594 19390 25596
rect 19414 25594 19470 25596
rect 19494 25594 19550 25596
rect 19574 25594 19630 25596
rect 19334 25542 19360 25594
rect 19360 25542 19390 25594
rect 19414 25542 19424 25594
rect 19424 25542 19470 25594
rect 19494 25542 19540 25594
rect 19540 25542 19550 25594
rect 19574 25542 19604 25594
rect 19604 25542 19630 25594
rect 19334 25540 19390 25542
rect 19414 25540 19470 25542
rect 19494 25540 19550 25542
rect 19574 25540 19630 25542
rect 23834 27512 23890 27568
rect 24478 26832 24534 26888
rect 23834 26152 23890 26208
rect 24478 25472 24534 25528
rect 24001 25050 24057 25052
rect 24081 25050 24137 25052
rect 24161 25050 24217 25052
rect 24241 25050 24297 25052
rect 24001 24998 24027 25050
rect 24027 24998 24057 25050
rect 24081 24998 24091 25050
rect 24091 24998 24137 25050
rect 24161 24998 24207 25050
rect 24207 24998 24217 25050
rect 24241 24998 24271 25050
rect 24271 24998 24297 25050
rect 24001 24996 24057 24998
rect 24081 24996 24137 24998
rect 24161 24996 24217 24998
rect 24241 24996 24297 24998
rect 19334 24506 19390 24508
rect 19414 24506 19470 24508
rect 19494 24506 19550 24508
rect 19574 24506 19630 24508
rect 19334 24454 19360 24506
rect 19360 24454 19390 24506
rect 19414 24454 19424 24506
rect 19424 24454 19470 24506
rect 19494 24454 19540 24506
rect 19540 24454 19550 24506
rect 19574 24454 19604 24506
rect 19604 24454 19630 24506
rect 19334 24452 19390 24454
rect 19414 24452 19470 24454
rect 19494 24452 19550 24454
rect 19574 24452 19630 24454
rect 19334 23418 19390 23420
rect 19414 23418 19470 23420
rect 19494 23418 19550 23420
rect 19574 23418 19630 23420
rect 19334 23366 19360 23418
rect 19360 23366 19390 23418
rect 19414 23366 19424 23418
rect 19424 23366 19470 23418
rect 19494 23366 19540 23418
rect 19540 23366 19550 23418
rect 19574 23366 19604 23418
rect 19604 23366 19630 23418
rect 19334 23364 19390 23366
rect 19414 23364 19470 23366
rect 19494 23364 19550 23366
rect 19574 23364 19630 23366
rect 19334 22330 19390 22332
rect 19414 22330 19470 22332
rect 19494 22330 19550 22332
rect 19574 22330 19630 22332
rect 19334 22278 19360 22330
rect 19360 22278 19390 22330
rect 19414 22278 19424 22330
rect 19424 22278 19470 22330
rect 19494 22278 19540 22330
rect 19540 22278 19550 22330
rect 19574 22278 19604 22330
rect 19604 22278 19630 22330
rect 19334 22276 19390 22278
rect 19414 22276 19470 22278
rect 19494 22276 19550 22278
rect 19574 22276 19630 22278
rect 19334 21242 19390 21244
rect 19414 21242 19470 21244
rect 19494 21242 19550 21244
rect 19574 21242 19630 21244
rect 19334 21190 19360 21242
rect 19360 21190 19390 21242
rect 19414 21190 19424 21242
rect 19424 21190 19470 21242
rect 19494 21190 19540 21242
rect 19540 21190 19550 21242
rect 19574 21190 19604 21242
rect 19604 21190 19630 21242
rect 19334 21188 19390 21190
rect 19414 21188 19470 21190
rect 19494 21188 19550 21190
rect 19574 21188 19630 21190
rect 19334 20154 19390 20156
rect 19414 20154 19470 20156
rect 19494 20154 19550 20156
rect 19574 20154 19630 20156
rect 19334 20102 19360 20154
rect 19360 20102 19390 20154
rect 19414 20102 19424 20154
rect 19424 20102 19470 20154
rect 19494 20102 19540 20154
rect 19540 20102 19550 20154
rect 19574 20102 19604 20154
rect 19604 20102 19630 20154
rect 19334 20100 19390 20102
rect 19414 20100 19470 20102
rect 19494 20100 19550 20102
rect 19574 20100 19630 20102
rect 19786 20032 19842 20088
rect 19786 19352 19842 19408
rect 23834 24792 23890 24848
rect 23374 23432 23430 23488
rect 24478 24112 24534 24168
rect 24001 23962 24057 23964
rect 24081 23962 24137 23964
rect 24161 23962 24217 23964
rect 24241 23962 24297 23964
rect 24001 23910 24027 23962
rect 24027 23910 24057 23962
rect 24081 23910 24091 23962
rect 24091 23910 24137 23962
rect 24161 23910 24207 23962
rect 24207 23910 24217 23962
rect 24241 23910 24271 23962
rect 24271 23910 24297 23962
rect 24001 23908 24057 23910
rect 24081 23908 24137 23910
rect 24161 23908 24217 23910
rect 24241 23908 24297 23910
rect 23834 23024 23890 23080
rect 24001 22874 24057 22876
rect 24081 22874 24137 22876
rect 24161 22874 24217 22876
rect 24241 22874 24297 22876
rect 24001 22822 24027 22874
rect 24027 22822 24057 22874
rect 24081 22822 24091 22874
rect 24091 22822 24137 22874
rect 24161 22822 24207 22874
rect 24207 22822 24217 22874
rect 24241 22822 24271 22874
rect 24271 22822 24297 22874
rect 24001 22820 24057 22822
rect 24081 22820 24137 22822
rect 24161 22820 24217 22822
rect 24241 22820 24297 22822
rect 24478 22480 24534 22536
rect 24478 22072 24534 22128
rect 23374 21936 23430 21992
rect 24001 21786 24057 21788
rect 24081 21786 24137 21788
rect 24161 21786 24217 21788
rect 24241 21786 24297 21788
rect 24001 21734 24027 21786
rect 24027 21734 24057 21786
rect 24081 21734 24091 21786
rect 24091 21734 24137 21786
rect 24161 21734 24207 21786
rect 24207 21734 24217 21786
rect 24241 21734 24271 21786
rect 24271 21734 24297 21786
rect 24001 21732 24057 21734
rect 24081 21732 24137 21734
rect 24161 21732 24217 21734
rect 24241 21732 24297 21734
rect 24386 20712 24442 20768
rect 24001 20698 24057 20700
rect 24081 20698 24137 20700
rect 24161 20698 24217 20700
rect 24241 20698 24297 20700
rect 24001 20646 24027 20698
rect 24027 20646 24057 20698
rect 24081 20646 24091 20698
rect 24091 20646 24137 20698
rect 24161 20646 24207 20698
rect 24207 20646 24217 20698
rect 24241 20646 24271 20698
rect 24271 20646 24297 20698
rect 24001 20644 24057 20646
rect 24081 20644 24137 20646
rect 24161 20644 24217 20646
rect 24241 20644 24297 20646
rect 24386 19896 24442 19952
rect 24001 19610 24057 19612
rect 24081 19610 24137 19612
rect 24161 19610 24217 19612
rect 24241 19610 24297 19612
rect 24001 19558 24027 19610
rect 24027 19558 24057 19610
rect 24081 19558 24091 19610
rect 24091 19558 24137 19610
rect 24161 19558 24207 19610
rect 24207 19558 24217 19610
rect 24241 19558 24271 19610
rect 24271 19558 24297 19610
rect 24001 19556 24057 19558
rect 24081 19556 24137 19558
rect 24161 19556 24217 19558
rect 24241 19556 24297 19558
rect 24386 19352 24442 19408
rect 19334 19066 19390 19068
rect 19414 19066 19470 19068
rect 19494 19066 19550 19068
rect 19574 19066 19630 19068
rect 19334 19014 19360 19066
rect 19360 19014 19390 19066
rect 19414 19014 19424 19066
rect 19424 19014 19470 19066
rect 19494 19014 19540 19066
rect 19540 19014 19550 19066
rect 19574 19014 19604 19066
rect 19604 19014 19630 19066
rect 19334 19012 19390 19014
rect 19414 19012 19470 19014
rect 19494 19012 19550 19014
rect 19574 19012 19630 19014
rect 19334 17978 19390 17980
rect 19414 17978 19470 17980
rect 19494 17978 19550 17980
rect 19574 17978 19630 17980
rect 19334 17926 19360 17978
rect 19360 17926 19390 17978
rect 19414 17926 19424 17978
rect 19424 17926 19470 17978
rect 19494 17926 19540 17978
rect 19540 17926 19550 17978
rect 19574 17926 19604 17978
rect 19604 17926 19630 17978
rect 19334 17924 19390 17926
rect 19414 17924 19470 17926
rect 19494 17924 19550 17926
rect 19574 17924 19630 17926
rect 16750 17040 16806 17096
rect 14668 16346 14724 16348
rect 14748 16346 14804 16348
rect 14828 16346 14884 16348
rect 14908 16346 14964 16348
rect 14668 16294 14694 16346
rect 14694 16294 14724 16346
rect 14748 16294 14758 16346
rect 14758 16294 14804 16346
rect 14828 16294 14874 16346
rect 14874 16294 14884 16346
rect 14908 16294 14938 16346
rect 14938 16294 14964 16346
rect 14668 16292 14724 16294
rect 14748 16292 14804 16294
rect 14828 16292 14884 16294
rect 14908 16292 14964 16294
rect 12426 13776 12482 13832
rect 12794 13796 12850 13832
rect 12794 13776 12796 13796
rect 12796 13776 12848 13796
rect 12848 13776 12850 13796
rect 12334 12688 12390 12744
rect 10494 3032 10550 3088
rect 10001 2746 10057 2748
rect 10081 2746 10137 2748
rect 10161 2746 10217 2748
rect 10241 2746 10297 2748
rect 10001 2694 10027 2746
rect 10027 2694 10057 2746
rect 10081 2694 10091 2746
rect 10091 2694 10137 2746
rect 10161 2694 10207 2746
rect 10207 2694 10217 2746
rect 10241 2694 10271 2746
rect 10271 2694 10297 2746
rect 10001 2692 10057 2694
rect 10081 2692 10137 2694
rect 10161 2692 10217 2694
rect 10241 2692 10297 2694
rect 17946 15408 18002 15464
rect 14668 15258 14724 15260
rect 14748 15258 14804 15260
rect 14828 15258 14884 15260
rect 14908 15258 14964 15260
rect 14668 15206 14694 15258
rect 14694 15206 14724 15258
rect 14748 15206 14758 15258
rect 14758 15206 14804 15258
rect 14828 15206 14874 15258
rect 14874 15206 14884 15258
rect 14908 15206 14938 15258
rect 14938 15206 14964 15258
rect 14668 15204 14724 15206
rect 14748 15204 14804 15206
rect 14828 15204 14884 15206
rect 14908 15204 14964 15206
rect 14668 14170 14724 14172
rect 14748 14170 14804 14172
rect 14828 14170 14884 14172
rect 14908 14170 14964 14172
rect 14668 14118 14694 14170
rect 14694 14118 14724 14170
rect 14748 14118 14758 14170
rect 14758 14118 14804 14170
rect 14828 14118 14874 14170
rect 14874 14118 14884 14170
rect 14908 14118 14938 14170
rect 14938 14118 14964 14170
rect 14668 14116 14724 14118
rect 14748 14116 14804 14118
rect 14828 14116 14884 14118
rect 14908 14116 14964 14118
rect 15462 13912 15518 13968
rect 14668 13082 14724 13084
rect 14748 13082 14804 13084
rect 14828 13082 14884 13084
rect 14908 13082 14964 13084
rect 14668 13030 14694 13082
rect 14694 13030 14724 13082
rect 14748 13030 14758 13082
rect 14758 13030 14804 13082
rect 14828 13030 14874 13082
rect 14874 13030 14884 13082
rect 14908 13030 14938 13082
rect 14938 13030 14964 13082
rect 14668 13028 14724 13030
rect 14748 13028 14804 13030
rect 14828 13028 14884 13030
rect 14908 13028 14964 13030
rect 14668 11994 14724 11996
rect 14748 11994 14804 11996
rect 14828 11994 14884 11996
rect 14908 11994 14964 11996
rect 14668 11942 14694 11994
rect 14694 11942 14724 11994
rect 14748 11942 14758 11994
rect 14758 11942 14804 11994
rect 14828 11942 14874 11994
rect 14874 11942 14884 11994
rect 14908 11942 14938 11994
rect 14938 11942 14964 11994
rect 14668 11940 14724 11942
rect 14748 11940 14804 11942
rect 14828 11940 14884 11942
rect 14908 11940 14964 11942
rect 14542 11500 14544 11520
rect 14544 11500 14596 11520
rect 14596 11500 14598 11520
rect 14542 11464 14598 11500
rect 17486 11192 17542 11248
rect 14668 10906 14724 10908
rect 14748 10906 14804 10908
rect 14828 10906 14884 10908
rect 14908 10906 14964 10908
rect 14668 10854 14694 10906
rect 14694 10854 14724 10906
rect 14748 10854 14758 10906
rect 14758 10854 14804 10906
rect 14828 10854 14874 10906
rect 14874 10854 14884 10906
rect 14908 10854 14938 10906
rect 14938 10854 14964 10906
rect 14668 10852 14724 10854
rect 14748 10852 14804 10854
rect 14828 10852 14884 10854
rect 14908 10852 14964 10854
rect 15278 10532 15334 10568
rect 15278 10512 15280 10532
rect 15280 10512 15332 10532
rect 15332 10512 15334 10532
rect 14668 9818 14724 9820
rect 14748 9818 14804 9820
rect 14828 9818 14884 9820
rect 14908 9818 14964 9820
rect 14668 9766 14694 9818
rect 14694 9766 14724 9818
rect 14748 9766 14758 9818
rect 14758 9766 14804 9818
rect 14828 9766 14874 9818
rect 14874 9766 14884 9818
rect 14908 9766 14938 9818
rect 14938 9766 14964 9818
rect 14668 9764 14724 9766
rect 14748 9764 14804 9766
rect 14828 9764 14884 9766
rect 14908 9764 14964 9766
rect 14910 9580 14966 9616
rect 14910 9560 14912 9580
rect 14912 9560 14964 9580
rect 14964 9560 14966 9580
rect 18406 9016 18462 9072
rect 14668 8730 14724 8732
rect 14748 8730 14804 8732
rect 14828 8730 14884 8732
rect 14908 8730 14964 8732
rect 14668 8678 14694 8730
rect 14694 8678 14724 8730
rect 14748 8678 14758 8730
rect 14758 8678 14804 8730
rect 14828 8678 14874 8730
rect 14874 8678 14884 8730
rect 14908 8678 14938 8730
rect 14938 8678 14964 8730
rect 14668 8676 14724 8678
rect 14748 8676 14804 8678
rect 14828 8676 14884 8678
rect 14908 8676 14964 8678
rect 16014 8508 16016 8528
rect 16016 8508 16068 8528
rect 16068 8508 16070 8528
rect 16014 8472 16070 8508
rect 14668 7642 14724 7644
rect 14748 7642 14804 7644
rect 14828 7642 14884 7644
rect 14908 7642 14964 7644
rect 14668 7590 14694 7642
rect 14694 7590 14724 7642
rect 14748 7590 14758 7642
rect 14758 7590 14804 7642
rect 14828 7590 14874 7642
rect 14874 7590 14884 7642
rect 14908 7590 14938 7642
rect 14938 7590 14964 7642
rect 14668 7588 14724 7590
rect 14748 7588 14804 7590
rect 14828 7588 14884 7590
rect 14908 7588 14964 7590
rect 14668 6554 14724 6556
rect 14748 6554 14804 6556
rect 14828 6554 14884 6556
rect 14908 6554 14964 6556
rect 14668 6502 14694 6554
rect 14694 6502 14724 6554
rect 14748 6502 14758 6554
rect 14758 6502 14804 6554
rect 14828 6502 14874 6554
rect 14874 6502 14884 6554
rect 14908 6502 14938 6554
rect 14938 6502 14964 6554
rect 14668 6500 14724 6502
rect 14748 6500 14804 6502
rect 14828 6500 14884 6502
rect 14908 6500 14964 6502
rect 14668 5466 14724 5468
rect 14748 5466 14804 5468
rect 14828 5466 14884 5468
rect 14908 5466 14964 5468
rect 14668 5414 14694 5466
rect 14694 5414 14724 5466
rect 14748 5414 14758 5466
rect 14758 5414 14804 5466
rect 14828 5414 14874 5466
rect 14874 5414 14884 5466
rect 14908 5414 14938 5466
rect 14938 5414 14964 5466
rect 14668 5412 14724 5414
rect 14748 5412 14804 5414
rect 14828 5412 14884 5414
rect 14908 5412 14964 5414
rect 14668 4378 14724 4380
rect 14748 4378 14804 4380
rect 14828 4378 14884 4380
rect 14908 4378 14964 4380
rect 14668 4326 14694 4378
rect 14694 4326 14724 4378
rect 14748 4326 14758 4378
rect 14758 4326 14804 4378
rect 14828 4326 14874 4378
rect 14874 4326 14884 4378
rect 14908 4326 14938 4378
rect 14938 4326 14964 4378
rect 14668 4324 14724 4326
rect 14748 4324 14804 4326
rect 14828 4324 14884 4326
rect 14908 4324 14964 4326
rect 14668 3290 14724 3292
rect 14748 3290 14804 3292
rect 14828 3290 14884 3292
rect 14908 3290 14964 3292
rect 14668 3238 14694 3290
rect 14694 3238 14724 3290
rect 14748 3238 14758 3290
rect 14758 3238 14804 3290
rect 14828 3238 14874 3290
rect 14874 3238 14884 3290
rect 14908 3238 14938 3290
rect 14938 3238 14964 3290
rect 14668 3236 14724 3238
rect 14748 3236 14804 3238
rect 14828 3236 14884 3238
rect 14908 3236 14964 3238
rect 14668 2202 14724 2204
rect 14748 2202 14804 2204
rect 14828 2202 14884 2204
rect 14908 2202 14964 2204
rect 14668 2150 14694 2202
rect 14694 2150 14724 2202
rect 14748 2150 14758 2202
rect 14758 2150 14804 2202
rect 14828 2150 14874 2202
rect 14874 2150 14884 2202
rect 14908 2150 14938 2202
rect 14938 2150 14964 2202
rect 14668 2148 14724 2150
rect 14748 2148 14804 2150
rect 14828 2148 14884 2150
rect 14908 2148 14964 2150
rect 17854 7928 17910 7984
rect 19334 16890 19390 16892
rect 19414 16890 19470 16892
rect 19494 16890 19550 16892
rect 19574 16890 19630 16892
rect 19334 16838 19360 16890
rect 19360 16838 19390 16890
rect 19414 16838 19424 16890
rect 19424 16838 19470 16890
rect 19494 16838 19540 16890
rect 19540 16838 19550 16890
rect 19574 16838 19604 16890
rect 19604 16838 19630 16890
rect 19334 16836 19390 16838
rect 19414 16836 19470 16838
rect 19494 16836 19550 16838
rect 19574 16836 19630 16838
rect 19694 16632 19750 16688
rect 19334 15802 19390 15804
rect 19414 15802 19470 15804
rect 19494 15802 19550 15804
rect 19574 15802 19630 15804
rect 19334 15750 19360 15802
rect 19360 15750 19390 15802
rect 19414 15750 19424 15802
rect 19424 15750 19470 15802
rect 19494 15750 19540 15802
rect 19540 15750 19550 15802
rect 19574 15750 19604 15802
rect 19604 15750 19630 15802
rect 19334 15748 19390 15750
rect 19414 15748 19470 15750
rect 19494 15748 19550 15750
rect 19574 15748 19630 15750
rect 21718 15544 21774 15600
rect 21718 15272 21774 15328
rect 19334 14714 19390 14716
rect 19414 14714 19470 14716
rect 19494 14714 19550 14716
rect 19574 14714 19630 14716
rect 19334 14662 19360 14714
rect 19360 14662 19390 14714
rect 19414 14662 19424 14714
rect 19424 14662 19470 14714
rect 19494 14662 19540 14714
rect 19540 14662 19550 14714
rect 19574 14662 19604 14714
rect 19604 14662 19630 14714
rect 19334 14660 19390 14662
rect 19414 14660 19470 14662
rect 19494 14660 19550 14662
rect 19574 14660 19630 14662
rect 19334 13626 19390 13628
rect 19414 13626 19470 13628
rect 19494 13626 19550 13628
rect 19574 13626 19630 13628
rect 19334 13574 19360 13626
rect 19360 13574 19390 13626
rect 19414 13574 19424 13626
rect 19424 13574 19470 13626
rect 19494 13574 19540 13626
rect 19540 13574 19550 13626
rect 19574 13574 19604 13626
rect 19604 13574 19630 13626
rect 19334 13572 19390 13574
rect 19414 13572 19470 13574
rect 19494 13572 19550 13574
rect 19574 13572 19630 13574
rect 19334 12538 19390 12540
rect 19414 12538 19470 12540
rect 19494 12538 19550 12540
rect 19574 12538 19630 12540
rect 19334 12486 19360 12538
rect 19360 12486 19390 12538
rect 19414 12486 19424 12538
rect 19424 12486 19470 12538
rect 19494 12486 19540 12538
rect 19540 12486 19550 12538
rect 19574 12486 19604 12538
rect 19604 12486 19630 12538
rect 19334 12484 19390 12486
rect 19414 12484 19470 12486
rect 19494 12484 19550 12486
rect 19574 12484 19630 12486
rect 21718 12552 21774 12608
rect 19334 11450 19390 11452
rect 19414 11450 19470 11452
rect 19494 11450 19550 11452
rect 19574 11450 19630 11452
rect 19334 11398 19360 11450
rect 19360 11398 19390 11450
rect 19414 11398 19424 11450
rect 19424 11398 19470 11450
rect 19494 11398 19540 11450
rect 19540 11398 19550 11450
rect 19574 11398 19604 11450
rect 19604 11398 19630 11450
rect 19334 11396 19390 11398
rect 19414 11396 19470 11398
rect 19494 11396 19550 11398
rect 19574 11396 19630 11398
rect 19334 10362 19390 10364
rect 19414 10362 19470 10364
rect 19494 10362 19550 10364
rect 19574 10362 19630 10364
rect 19334 10310 19360 10362
rect 19360 10310 19390 10362
rect 19414 10310 19424 10362
rect 19424 10310 19470 10362
rect 19494 10310 19540 10362
rect 19540 10310 19550 10362
rect 19574 10310 19604 10362
rect 19604 10310 19630 10362
rect 19334 10308 19390 10310
rect 19414 10308 19470 10310
rect 19494 10308 19550 10310
rect 19574 10308 19630 10310
rect 18958 9696 19014 9752
rect 18866 9560 18922 9616
rect 21074 10920 21130 10976
rect 20614 9696 20670 9752
rect 19334 9274 19390 9276
rect 19414 9274 19470 9276
rect 19494 9274 19550 9276
rect 19574 9274 19630 9276
rect 19334 9222 19360 9274
rect 19360 9222 19390 9274
rect 19414 9222 19424 9274
rect 19424 9222 19470 9274
rect 19494 9222 19540 9274
rect 19540 9222 19550 9274
rect 19574 9222 19604 9274
rect 19604 9222 19630 9274
rect 19334 9220 19390 9222
rect 19414 9220 19470 9222
rect 19494 9220 19550 9222
rect 19574 9220 19630 9222
rect 23650 18672 23706 18728
rect 24001 18522 24057 18524
rect 24081 18522 24137 18524
rect 24161 18522 24217 18524
rect 24241 18522 24297 18524
rect 24001 18470 24027 18522
rect 24027 18470 24057 18522
rect 24081 18470 24091 18522
rect 24091 18470 24137 18522
rect 24161 18470 24207 18522
rect 24207 18470 24217 18522
rect 24241 18470 24271 18522
rect 24271 18470 24297 18522
rect 24001 18468 24057 18470
rect 24081 18468 24137 18470
rect 24161 18468 24217 18470
rect 24241 18468 24297 18470
rect 23926 17992 23982 18048
rect 23650 17312 23706 17368
rect 24386 17584 24442 17640
rect 24001 17434 24057 17436
rect 24081 17434 24137 17436
rect 24161 17434 24217 17436
rect 24241 17434 24297 17436
rect 24001 17382 24027 17434
rect 24027 17382 24057 17434
rect 24081 17382 24091 17434
rect 24091 17382 24137 17434
rect 24161 17382 24207 17434
rect 24207 17382 24217 17434
rect 24241 17382 24271 17434
rect 24271 17382 24297 17434
rect 24001 17380 24057 17382
rect 24081 17380 24137 17382
rect 24161 17380 24217 17382
rect 24241 17380 24297 17382
rect 23926 17176 23982 17232
rect 24001 16346 24057 16348
rect 24081 16346 24137 16348
rect 24161 16346 24217 16348
rect 24241 16346 24297 16348
rect 24001 16294 24027 16346
rect 24027 16294 24057 16346
rect 24081 16294 24091 16346
rect 24091 16294 24137 16346
rect 24161 16294 24207 16346
rect 24207 16294 24217 16346
rect 24241 16294 24271 16346
rect 24271 16294 24297 16346
rect 24001 16292 24057 16294
rect 24081 16292 24137 16294
rect 24161 16292 24217 16294
rect 24241 16292 24297 16294
rect 24001 15258 24057 15260
rect 24081 15258 24137 15260
rect 24161 15258 24217 15260
rect 24241 15258 24297 15260
rect 24001 15206 24027 15258
rect 24027 15206 24057 15258
rect 24081 15206 24091 15258
rect 24091 15206 24137 15258
rect 24161 15206 24207 15258
rect 24207 15206 24217 15258
rect 24241 15206 24271 15258
rect 24271 15206 24297 15258
rect 24001 15204 24057 15206
rect 24081 15204 24137 15206
rect 24161 15204 24217 15206
rect 24241 15204 24297 15206
rect 23834 14592 23890 14648
rect 24001 14170 24057 14172
rect 24081 14170 24137 14172
rect 24161 14170 24217 14172
rect 24241 14170 24297 14172
rect 24001 14118 24027 14170
rect 24027 14118 24057 14170
rect 24081 14118 24091 14170
rect 24091 14118 24137 14170
rect 24161 14118 24207 14170
rect 24207 14118 24217 14170
rect 24241 14118 24271 14170
rect 24271 14118 24297 14170
rect 24001 14116 24057 14118
rect 24081 14116 24137 14118
rect 24161 14116 24217 14118
rect 24241 14116 24297 14118
rect 24478 13232 24534 13288
rect 24001 13082 24057 13084
rect 24081 13082 24137 13084
rect 24161 13082 24217 13084
rect 24241 13082 24297 13084
rect 24001 13030 24027 13082
rect 24027 13030 24057 13082
rect 24081 13030 24091 13082
rect 24091 13030 24137 13082
rect 24161 13030 24207 13082
rect 24207 13030 24217 13082
rect 24241 13030 24271 13082
rect 24271 13030 24297 13082
rect 24001 13028 24057 13030
rect 24081 13028 24137 13030
rect 24161 13028 24217 13030
rect 24241 13028 24297 13030
rect 23834 12960 23890 13016
rect 23558 12724 23560 12744
rect 23560 12724 23612 12744
rect 23612 12724 23614 12744
rect 23558 12688 23614 12724
rect 23190 12552 23246 12608
rect 24001 11994 24057 11996
rect 24081 11994 24137 11996
rect 24161 11994 24217 11996
rect 24241 11994 24297 11996
rect 24001 11942 24027 11994
rect 24027 11942 24057 11994
rect 24081 11942 24091 11994
rect 24091 11942 24137 11994
rect 24161 11942 24207 11994
rect 24207 11942 24217 11994
rect 24241 11942 24271 11994
rect 24271 11942 24297 11994
rect 24001 11940 24057 11942
rect 24081 11940 24137 11942
rect 24161 11940 24217 11942
rect 24241 11940 24297 11942
rect 23742 11736 23798 11792
rect 24001 10906 24057 10908
rect 24081 10906 24137 10908
rect 24161 10906 24217 10908
rect 24241 10906 24297 10908
rect 24001 10854 24027 10906
rect 24027 10854 24057 10906
rect 24081 10854 24091 10906
rect 24091 10854 24137 10906
rect 24161 10854 24207 10906
rect 24207 10854 24217 10906
rect 24241 10854 24271 10906
rect 24271 10854 24297 10906
rect 24001 10852 24057 10854
rect 24081 10852 24137 10854
rect 24161 10852 24217 10854
rect 24241 10852 24297 10854
rect 23742 10512 23798 10568
rect 23926 10512 23982 10568
rect 23190 9968 23246 10024
rect 19334 8186 19390 8188
rect 19414 8186 19470 8188
rect 19494 8186 19550 8188
rect 19574 8186 19630 8188
rect 19334 8134 19360 8186
rect 19360 8134 19390 8186
rect 19414 8134 19424 8186
rect 19424 8134 19470 8186
rect 19494 8134 19540 8186
rect 19540 8134 19550 8186
rect 19574 8134 19604 8186
rect 19604 8134 19630 8186
rect 19334 8132 19390 8134
rect 19414 8132 19470 8134
rect 19494 8132 19550 8134
rect 19574 8132 19630 8134
rect 19334 7098 19390 7100
rect 19414 7098 19470 7100
rect 19494 7098 19550 7100
rect 19574 7098 19630 7100
rect 19334 7046 19360 7098
rect 19360 7046 19390 7098
rect 19414 7046 19424 7098
rect 19424 7046 19470 7098
rect 19494 7046 19540 7098
rect 19540 7046 19550 7098
rect 19574 7046 19604 7098
rect 19604 7046 19630 7098
rect 19334 7044 19390 7046
rect 19414 7044 19470 7046
rect 19494 7044 19550 7046
rect 19574 7044 19630 7046
rect 18774 3576 18830 3632
rect 19694 6840 19750 6896
rect 19234 6316 19290 6352
rect 19234 6296 19236 6316
rect 19236 6296 19288 6316
rect 19288 6296 19290 6316
rect 19334 6010 19390 6012
rect 19414 6010 19470 6012
rect 19494 6010 19550 6012
rect 19574 6010 19630 6012
rect 19334 5958 19360 6010
rect 19360 5958 19390 6010
rect 19414 5958 19424 6010
rect 19424 5958 19470 6010
rect 19494 5958 19540 6010
rect 19540 5958 19550 6010
rect 19574 5958 19604 6010
rect 19604 5958 19630 6010
rect 19334 5956 19390 5958
rect 19414 5956 19470 5958
rect 19494 5956 19550 5958
rect 19574 5956 19630 5958
rect 24478 10104 24534 10160
rect 27238 10104 27294 10160
rect 24001 9818 24057 9820
rect 24081 9818 24137 9820
rect 24161 9818 24217 9820
rect 24241 9818 24297 9820
rect 24001 9766 24027 9818
rect 24027 9766 24057 9818
rect 24081 9766 24091 9818
rect 24091 9766 24137 9818
rect 24161 9766 24207 9818
rect 24207 9766 24217 9818
rect 24241 9766 24271 9818
rect 24271 9766 24297 9818
rect 24001 9764 24057 9766
rect 24081 9764 24137 9766
rect 24161 9764 24217 9766
rect 24241 9764 24297 9766
rect 24001 8730 24057 8732
rect 24081 8730 24137 8732
rect 24161 8730 24217 8732
rect 24241 8730 24297 8732
rect 24001 8678 24027 8730
rect 24027 8678 24057 8730
rect 24081 8678 24091 8730
rect 24091 8678 24137 8730
rect 24161 8678 24207 8730
rect 24207 8678 24217 8730
rect 24241 8678 24271 8730
rect 24271 8678 24297 8730
rect 24001 8676 24057 8678
rect 24081 8676 24137 8678
rect 24161 8676 24217 8678
rect 24241 8676 24297 8678
rect 23926 8472 23982 8528
rect 24478 7792 24534 7848
rect 24001 7642 24057 7644
rect 24081 7642 24137 7644
rect 24161 7642 24217 7644
rect 24241 7642 24297 7644
rect 24001 7590 24027 7642
rect 24027 7590 24057 7642
rect 24081 7590 24091 7642
rect 24091 7590 24137 7642
rect 24161 7590 24207 7642
rect 24207 7590 24217 7642
rect 24241 7590 24271 7642
rect 24271 7590 24297 7642
rect 24001 7588 24057 7590
rect 24081 7588 24137 7590
rect 24161 7588 24217 7590
rect 24241 7588 24297 7590
rect 21534 5752 21590 5808
rect 19334 4922 19390 4924
rect 19414 4922 19470 4924
rect 19494 4922 19550 4924
rect 19574 4922 19630 4924
rect 19334 4870 19360 4922
rect 19360 4870 19390 4922
rect 19414 4870 19424 4922
rect 19424 4870 19470 4922
rect 19494 4870 19540 4922
rect 19540 4870 19550 4922
rect 19574 4870 19604 4922
rect 19604 4870 19630 4922
rect 19334 4868 19390 4870
rect 19414 4868 19470 4870
rect 19494 4868 19550 4870
rect 19574 4868 19630 4870
rect 19334 3834 19390 3836
rect 19414 3834 19470 3836
rect 19494 3834 19550 3836
rect 19574 3834 19630 3836
rect 19334 3782 19360 3834
rect 19360 3782 19390 3834
rect 19414 3782 19424 3834
rect 19424 3782 19470 3834
rect 19494 3782 19540 3834
rect 19540 3782 19550 3834
rect 19574 3782 19604 3834
rect 19604 3782 19630 3834
rect 19334 3780 19390 3782
rect 19414 3780 19470 3782
rect 19494 3780 19550 3782
rect 19574 3780 19630 3782
rect 19334 2746 19390 2748
rect 19414 2746 19470 2748
rect 19494 2746 19550 2748
rect 19574 2746 19630 2748
rect 19334 2694 19360 2746
rect 19360 2694 19390 2746
rect 19414 2694 19424 2746
rect 19424 2694 19470 2746
rect 19494 2694 19540 2746
rect 19540 2694 19550 2746
rect 19574 2694 19604 2746
rect 19604 2694 19630 2746
rect 19334 2692 19390 2694
rect 19414 2692 19470 2694
rect 19494 2692 19550 2694
rect 19574 2692 19630 2694
rect 20154 4664 20210 4720
rect 21442 4664 21498 4720
rect 24001 6554 24057 6556
rect 24081 6554 24137 6556
rect 24161 6554 24217 6556
rect 24241 6554 24297 6556
rect 24001 6502 24027 6554
rect 24027 6502 24057 6554
rect 24081 6502 24091 6554
rect 24091 6502 24137 6554
rect 24161 6502 24207 6554
rect 24207 6502 24217 6554
rect 24241 6502 24271 6554
rect 24271 6502 24297 6554
rect 24001 6500 24057 6502
rect 24081 6500 24137 6502
rect 24161 6500 24217 6502
rect 24241 6500 24297 6502
rect 24386 6432 24442 6488
rect 24001 5466 24057 5468
rect 24081 5466 24137 5468
rect 24161 5466 24217 5468
rect 24241 5466 24297 5468
rect 24001 5414 24027 5466
rect 24027 5414 24057 5466
rect 24081 5414 24091 5466
rect 24091 5414 24137 5466
rect 24161 5414 24207 5466
rect 24207 5414 24217 5466
rect 24241 5414 24271 5466
rect 24271 5414 24297 5466
rect 24001 5412 24057 5414
rect 24081 5412 24137 5414
rect 24161 5412 24217 5414
rect 24241 5412 24297 5414
rect 24294 5072 24350 5128
rect 24478 6296 24534 6352
rect 21626 4120 21682 4176
rect 20982 3440 21038 3496
rect 24001 4378 24057 4380
rect 24081 4378 24137 4380
rect 24161 4378 24217 4380
rect 24241 4378 24297 4380
rect 24001 4326 24027 4378
rect 24027 4326 24057 4378
rect 24081 4326 24091 4378
rect 24091 4326 24137 4378
rect 24161 4326 24207 4378
rect 24207 4326 24217 4378
rect 24241 4326 24271 4378
rect 24271 4326 24297 4378
rect 24001 4324 24057 4326
rect 24081 4324 24137 4326
rect 24161 4324 24217 4326
rect 24241 4324 24297 4326
rect 24478 4120 24534 4176
rect 23650 3032 23706 3088
rect 22730 2896 22786 2952
rect 23282 992 23338 1048
rect 24001 3290 24057 3292
rect 24081 3290 24137 3292
rect 24161 3290 24217 3292
rect 24241 3290 24297 3292
rect 24001 3238 24027 3290
rect 24027 3238 24057 3290
rect 24081 3238 24091 3290
rect 24091 3238 24137 3290
rect 24161 3238 24207 3290
rect 24207 3238 24217 3290
rect 24241 3238 24271 3290
rect 24271 3238 24297 3290
rect 24001 3236 24057 3238
rect 24081 3236 24137 3238
rect 24161 3236 24217 3238
rect 24241 3236 24297 3238
rect 24478 3304 24534 3360
rect 24478 3168 24534 3224
rect 24001 2202 24057 2204
rect 24081 2202 24137 2204
rect 24161 2202 24217 2204
rect 24241 2202 24297 2204
rect 24001 2150 24027 2202
rect 24027 2150 24057 2202
rect 24081 2150 24091 2202
rect 24091 2150 24137 2202
rect 24161 2150 24207 2202
rect 24207 2150 24217 2202
rect 24241 2150 24271 2202
rect 24271 2150 24297 2202
rect 24001 2148 24057 2150
rect 24081 2148 24137 2150
rect 24161 2148 24217 2150
rect 24241 2148 24297 2150
rect 24386 1672 24442 1728
rect 26594 3304 26650 3360
rect 25858 2896 25914 2952
rect 25306 2796 25308 2816
rect 25308 2796 25360 2816
rect 25360 2796 25362 2816
rect 25306 2760 25362 2796
rect 23926 312 23982 368
<< metal3 >>
rect 23829 27570 23895 27573
rect 27232 27570 27712 27600
rect 23829 27568 27712 27570
rect 23829 27512 23834 27568
rect 23890 27512 27712 27568
rect 23829 27510 27712 27512
rect 23829 27507 23895 27510
rect 27232 27480 27712 27510
rect 24473 26890 24539 26893
rect 27232 26890 27712 26920
rect 24473 26888 27712 26890
rect 24473 26832 24478 26888
rect 24534 26832 27712 26888
rect 24473 26830 27712 26832
rect 24473 26827 24539 26830
rect 27232 26800 27712 26830
rect 23829 26210 23895 26213
rect 27232 26210 27712 26240
rect 23829 26208 27712 26210
rect 23829 26152 23834 26208
rect 23890 26152 27712 26208
rect 23829 26150 27712 26152
rect 23829 26147 23895 26150
rect 27232 26120 27712 26150
rect 9989 25600 10309 25601
rect 9989 25536 9997 25600
rect 10061 25536 10077 25600
rect 10141 25536 10157 25600
rect 10221 25536 10237 25600
rect 10301 25536 10309 25600
rect 9989 25535 10309 25536
rect 19322 25600 19642 25601
rect 19322 25536 19330 25600
rect 19394 25536 19410 25600
rect 19474 25536 19490 25600
rect 19554 25536 19570 25600
rect 19634 25536 19642 25600
rect 19322 25535 19642 25536
rect 24473 25530 24539 25533
rect 27232 25530 27712 25560
rect 24473 25528 27712 25530
rect 24473 25472 24478 25528
rect 24534 25472 27712 25528
rect 24473 25470 27712 25472
rect 24473 25467 24539 25470
rect 27232 25440 27712 25470
rect 5322 25056 5642 25057
rect 5322 24992 5330 25056
rect 5394 24992 5410 25056
rect 5474 24992 5490 25056
rect 5554 24992 5570 25056
rect 5634 24992 5642 25056
rect 5322 24991 5642 24992
rect 14656 25056 14976 25057
rect 14656 24992 14664 25056
rect 14728 24992 14744 25056
rect 14808 24992 14824 25056
rect 14888 24992 14904 25056
rect 14968 24992 14976 25056
rect 14656 24991 14976 24992
rect 23989 25056 24309 25057
rect 23989 24992 23997 25056
rect 24061 24992 24077 25056
rect 24141 24992 24157 25056
rect 24221 24992 24237 25056
rect 24301 24992 24309 25056
rect 23989 24991 24309 24992
rect 23829 24850 23895 24853
rect 27232 24850 27712 24880
rect 23829 24848 27712 24850
rect 23829 24792 23834 24848
rect 23890 24792 27712 24848
rect 23829 24790 27712 24792
rect 23829 24787 23895 24790
rect 27232 24760 27712 24790
rect 9989 24512 10309 24513
rect 9989 24448 9997 24512
rect 10061 24448 10077 24512
rect 10141 24448 10157 24512
rect 10221 24448 10237 24512
rect 10301 24448 10309 24512
rect 9989 24447 10309 24448
rect 19322 24512 19642 24513
rect 19322 24448 19330 24512
rect 19394 24448 19410 24512
rect 19474 24448 19490 24512
rect 19554 24448 19570 24512
rect 19634 24448 19642 24512
rect 19322 24447 19642 24448
rect 24473 24170 24539 24173
rect 27232 24170 27712 24200
rect 24473 24168 27712 24170
rect 24473 24112 24478 24168
rect 24534 24112 27712 24168
rect 24473 24110 27712 24112
rect 24473 24107 24539 24110
rect 27232 24080 27712 24110
rect 5322 23968 5642 23969
rect 5322 23904 5330 23968
rect 5394 23904 5410 23968
rect 5474 23904 5490 23968
rect 5554 23904 5570 23968
rect 5634 23904 5642 23968
rect 5322 23903 5642 23904
rect 14656 23968 14976 23969
rect 14656 23904 14664 23968
rect 14728 23904 14744 23968
rect 14808 23904 14824 23968
rect 14888 23904 14904 23968
rect 14968 23904 14976 23968
rect 14656 23903 14976 23904
rect 23989 23968 24309 23969
rect 23989 23904 23997 23968
rect 24061 23904 24077 23968
rect 24141 23904 24157 23968
rect 24221 23904 24237 23968
rect 24301 23904 24309 23968
rect 23989 23903 24309 23904
rect 23369 23490 23435 23493
rect 27232 23490 27712 23520
rect 23369 23488 27712 23490
rect 23369 23432 23374 23488
rect 23430 23432 27712 23488
rect 23369 23430 27712 23432
rect 23369 23427 23435 23430
rect 9989 23424 10309 23425
rect 9989 23360 9997 23424
rect 10061 23360 10077 23424
rect 10141 23360 10157 23424
rect 10221 23360 10237 23424
rect 10301 23360 10309 23424
rect 9989 23359 10309 23360
rect 19322 23424 19642 23425
rect 19322 23360 19330 23424
rect 19394 23360 19410 23424
rect 19474 23360 19490 23424
rect 19554 23360 19570 23424
rect 19634 23360 19642 23424
rect 27232 23400 27712 23430
rect 19322 23359 19642 23360
rect 2025 23082 2091 23085
rect 23829 23082 23895 23085
rect 2025 23080 23895 23082
rect 2025 23024 2030 23080
rect 2086 23024 23834 23080
rect 23890 23024 23895 23080
rect 2025 23022 23895 23024
rect 2025 23019 2091 23022
rect 23829 23019 23895 23022
rect 5705 22946 5771 22949
rect 14445 22946 14511 22949
rect 5705 22944 14511 22946
rect 5705 22888 5710 22944
rect 5766 22888 14450 22944
rect 14506 22888 14511 22944
rect 5705 22886 14511 22888
rect 5705 22883 5771 22886
rect 14445 22883 14511 22886
rect 15089 22946 15155 22949
rect 15089 22944 23754 22946
rect 15089 22888 15094 22944
rect 15150 22888 23754 22944
rect 15089 22886 23754 22888
rect 15089 22883 15155 22886
rect 5322 22880 5642 22881
rect 5322 22816 5330 22880
rect 5394 22816 5410 22880
rect 5474 22816 5490 22880
rect 5554 22816 5570 22880
rect 5634 22816 5642 22880
rect 5322 22815 5642 22816
rect 14656 22880 14976 22881
rect 14656 22816 14664 22880
rect 14728 22816 14744 22880
rect 14808 22816 14824 22880
rect 14888 22816 14904 22880
rect 14968 22816 14976 22880
rect 14656 22815 14976 22816
rect 23694 22674 23754 22886
rect 23989 22880 24309 22881
rect 23989 22816 23997 22880
rect 24061 22816 24077 22880
rect 24141 22816 24157 22880
rect 24221 22816 24237 22880
rect 24301 22816 24309 22880
rect 23989 22815 24309 22816
rect 27232 22810 27712 22840
rect 24430 22750 27712 22810
rect 24430 22674 24490 22750
rect 27232 22720 27712 22750
rect 23694 22614 24490 22674
rect 2669 22538 2735 22541
rect 24473 22538 24539 22541
rect 2669 22536 24539 22538
rect 2669 22480 2674 22536
rect 2730 22480 24478 22536
rect 24534 22480 24539 22536
rect 2669 22478 24539 22480
rect 2669 22475 2735 22478
rect 24473 22475 24539 22478
rect 4049 22402 4115 22405
rect 5705 22402 5771 22405
rect 4049 22400 5771 22402
rect 4049 22344 4054 22400
rect 4110 22344 5710 22400
rect 5766 22344 5771 22400
rect 4049 22342 5771 22344
rect 4049 22339 4115 22342
rect 5705 22339 5771 22342
rect 9989 22336 10309 22337
rect 9989 22272 9997 22336
rect 10061 22272 10077 22336
rect 10141 22272 10157 22336
rect 10221 22272 10237 22336
rect 10301 22272 10309 22336
rect 9989 22271 10309 22272
rect 19322 22336 19642 22337
rect 19322 22272 19330 22336
rect 19394 22272 19410 22336
rect 19474 22272 19490 22336
rect 19554 22272 19570 22336
rect 19634 22272 19642 22336
rect 19322 22271 19642 22272
rect 24473 22130 24539 22133
rect 27232 22130 27712 22160
rect 24473 22128 27712 22130
rect 24473 22072 24478 22128
rect 24534 22072 27712 22128
rect 24473 22070 27712 22072
rect 24473 22067 24539 22070
rect 27232 22040 27712 22070
rect 3957 21994 4023 21997
rect 23369 21994 23435 21997
rect 3957 21992 23435 21994
rect 3957 21936 3962 21992
rect 4018 21936 23374 21992
rect 23430 21936 23435 21992
rect 3957 21934 23435 21936
rect 3957 21931 4023 21934
rect 23369 21931 23435 21934
rect 5322 21792 5642 21793
rect 5322 21728 5330 21792
rect 5394 21728 5410 21792
rect 5474 21728 5490 21792
rect 5554 21728 5570 21792
rect 5634 21728 5642 21792
rect 5322 21727 5642 21728
rect 14656 21792 14976 21793
rect 14656 21728 14664 21792
rect 14728 21728 14744 21792
rect 14808 21728 14824 21792
rect 14888 21728 14904 21792
rect 14968 21728 14976 21792
rect 14656 21727 14976 21728
rect 23989 21792 24309 21793
rect 23989 21728 23997 21792
rect 24061 21728 24077 21792
rect 24141 21728 24157 21792
rect 24221 21728 24237 21792
rect 24301 21728 24309 21792
rect 23989 21727 24309 21728
rect 27232 21450 27712 21480
rect 27190 21360 27712 21450
rect 9989 21248 10309 21249
rect 9989 21184 9997 21248
rect 10061 21184 10077 21248
rect 10141 21184 10157 21248
rect 10221 21184 10237 21248
rect 10301 21184 10309 21248
rect 9989 21183 10309 21184
rect 19322 21248 19642 21249
rect 19322 21184 19330 21248
rect 19394 21184 19410 21248
rect 19474 21184 19490 21248
rect 19554 21184 19570 21248
rect 19634 21184 19642 21248
rect 19322 21183 19642 21184
rect 14169 21042 14235 21045
rect 27190 21042 27250 21360
rect 14169 21040 27250 21042
rect 14169 20984 14174 21040
rect 14230 20984 27250 21040
rect 14169 20982 27250 20984
rect 14169 20979 14235 20982
rect 5705 20906 5771 20909
rect 9334 20906 9340 20908
rect 5705 20904 9340 20906
rect 5705 20848 5710 20904
rect 5766 20848 9340 20904
rect 5705 20846 9340 20848
rect 5705 20843 5771 20846
rect 9334 20844 9340 20846
rect 9404 20844 9410 20908
rect 24381 20770 24447 20773
rect 27232 20770 27712 20800
rect 24381 20768 27712 20770
rect 24381 20712 24386 20768
rect 24442 20712 27712 20768
rect 24381 20710 27712 20712
rect 24381 20707 24447 20710
rect 5322 20704 5642 20705
rect 5322 20640 5330 20704
rect 5394 20640 5410 20704
rect 5474 20640 5490 20704
rect 5554 20640 5570 20704
rect 5634 20640 5642 20704
rect 5322 20639 5642 20640
rect 14656 20704 14976 20705
rect 14656 20640 14664 20704
rect 14728 20640 14744 20704
rect 14808 20640 14824 20704
rect 14888 20640 14904 20704
rect 14968 20640 14976 20704
rect 14656 20639 14976 20640
rect 23989 20704 24309 20705
rect 23989 20640 23997 20704
rect 24061 20640 24077 20704
rect 24141 20640 24157 20704
rect 24221 20640 24237 20704
rect 24301 20640 24309 20704
rect 27232 20680 27712 20710
rect 23989 20639 24309 20640
rect 9334 20572 9340 20636
rect 9404 20634 9410 20636
rect 14169 20634 14235 20637
rect 9404 20632 14235 20634
rect 9404 20576 14174 20632
rect 14230 20576 14235 20632
rect 9404 20574 14235 20576
rect 9404 20572 9410 20574
rect 14169 20571 14235 20574
rect 9989 20160 10309 20161
rect 9989 20096 9997 20160
rect 10061 20096 10077 20160
rect 10141 20096 10157 20160
rect 10221 20096 10237 20160
rect 10301 20096 10309 20160
rect 9989 20095 10309 20096
rect 19322 20160 19642 20161
rect 19322 20096 19330 20160
rect 19394 20096 19410 20160
rect 19474 20096 19490 20160
rect 19554 20096 19570 20160
rect 19634 20096 19642 20160
rect 19322 20095 19642 20096
rect 19781 20090 19847 20093
rect 27232 20090 27712 20120
rect 19781 20088 27712 20090
rect 19781 20032 19786 20088
rect 19842 20032 27712 20088
rect 19781 20030 27712 20032
rect 19781 20027 19847 20030
rect 27232 20000 27712 20030
rect 6717 19954 6783 19957
rect 24381 19954 24447 19957
rect 6717 19952 24447 19954
rect 6717 19896 6722 19952
rect 6778 19896 24386 19952
rect 24442 19896 24447 19952
rect 6717 19894 24447 19896
rect 6717 19891 6783 19894
rect 24381 19891 24447 19894
rect 5322 19616 5642 19617
rect 5322 19552 5330 19616
rect 5394 19552 5410 19616
rect 5474 19552 5490 19616
rect 5554 19552 5570 19616
rect 5634 19552 5642 19616
rect 5322 19551 5642 19552
rect 14656 19616 14976 19617
rect 14656 19552 14664 19616
rect 14728 19552 14744 19616
rect 14808 19552 14824 19616
rect 14888 19552 14904 19616
rect 14968 19552 14976 19616
rect 14656 19551 14976 19552
rect 23989 19616 24309 19617
rect 23989 19552 23997 19616
rect 24061 19552 24077 19616
rect 24141 19552 24157 19616
rect 24221 19552 24237 19616
rect 24301 19552 24309 19616
rect 23989 19551 24309 19552
rect 6809 19410 6875 19413
rect 19781 19410 19847 19413
rect 6809 19408 19847 19410
rect 6809 19352 6814 19408
rect 6870 19352 19786 19408
rect 19842 19352 19847 19408
rect 6809 19350 19847 19352
rect 6809 19347 6875 19350
rect 19781 19347 19847 19350
rect 24381 19410 24447 19413
rect 27232 19410 27712 19440
rect 24381 19408 27712 19410
rect 24381 19352 24386 19408
rect 24442 19352 27712 19408
rect 24381 19350 27712 19352
rect 24381 19347 24447 19350
rect 27232 19320 27712 19350
rect 9989 19072 10309 19073
rect 9989 19008 9997 19072
rect 10061 19008 10077 19072
rect 10141 19008 10157 19072
rect 10221 19008 10237 19072
rect 10301 19008 10309 19072
rect 9989 19007 10309 19008
rect 19322 19072 19642 19073
rect 19322 19008 19330 19072
rect 19394 19008 19410 19072
rect 19474 19008 19490 19072
rect 19554 19008 19570 19072
rect 19634 19008 19642 19072
rect 19322 19007 19642 19008
rect 23645 18730 23711 18733
rect 27232 18730 27712 18760
rect 23645 18728 27712 18730
rect 23645 18672 23650 18728
rect 23706 18672 27712 18728
rect 23645 18670 27712 18672
rect 23645 18667 23711 18670
rect 27232 18640 27712 18670
rect 5322 18528 5642 18529
rect 5322 18464 5330 18528
rect 5394 18464 5410 18528
rect 5474 18464 5490 18528
rect 5554 18464 5570 18528
rect 5634 18464 5642 18528
rect 5322 18463 5642 18464
rect 14656 18528 14976 18529
rect 14656 18464 14664 18528
rect 14728 18464 14744 18528
rect 14808 18464 14824 18528
rect 14888 18464 14904 18528
rect 14968 18464 14976 18528
rect 14656 18463 14976 18464
rect 23989 18528 24309 18529
rect 23989 18464 23997 18528
rect 24061 18464 24077 18528
rect 24141 18464 24157 18528
rect 24221 18464 24237 18528
rect 24301 18464 24309 18528
rect 23989 18463 24309 18464
rect 23921 18050 23987 18053
rect 27232 18050 27712 18080
rect 23921 18048 27712 18050
rect 23921 17992 23926 18048
rect 23982 17992 27712 18048
rect 23921 17990 27712 17992
rect 23921 17987 23987 17990
rect 9989 17984 10309 17985
rect 9989 17920 9997 17984
rect 10061 17920 10077 17984
rect 10141 17920 10157 17984
rect 10221 17920 10237 17984
rect 10301 17920 10309 17984
rect 9989 17919 10309 17920
rect 19322 17984 19642 17985
rect 19322 17920 19330 17984
rect 19394 17920 19410 17984
rect 19474 17920 19490 17984
rect 19554 17920 19570 17984
rect 19634 17920 19642 17984
rect 27232 17960 27712 17990
rect 19322 17919 19642 17920
rect 7453 17642 7519 17645
rect 24381 17642 24447 17645
rect 7453 17640 24447 17642
rect 7453 17584 7458 17640
rect 7514 17584 24386 17640
rect 24442 17584 24447 17640
rect 7453 17582 24447 17584
rect 7453 17579 7519 17582
rect 24381 17579 24447 17582
rect 5322 17440 5642 17441
rect 5322 17376 5330 17440
rect 5394 17376 5410 17440
rect 5474 17376 5490 17440
rect 5554 17376 5570 17440
rect 5634 17376 5642 17440
rect 5322 17375 5642 17376
rect 14656 17440 14976 17441
rect 14656 17376 14664 17440
rect 14728 17376 14744 17440
rect 14808 17376 14824 17440
rect 14888 17376 14904 17440
rect 14968 17376 14976 17440
rect 14656 17375 14976 17376
rect 23989 17440 24309 17441
rect 23989 17376 23997 17440
rect 24061 17376 24077 17440
rect 24141 17376 24157 17440
rect 24221 17376 24237 17440
rect 24301 17376 24309 17440
rect 23989 17375 24309 17376
rect 16745 17370 16811 17373
rect 23645 17370 23711 17373
rect 27232 17370 27712 17400
rect 16745 17368 23711 17370
rect 16745 17312 16750 17368
rect 16806 17312 23650 17368
rect 23706 17312 23711 17368
rect 16745 17310 23711 17312
rect 16745 17307 16811 17310
rect 23645 17307 23711 17310
rect 24614 17310 27712 17370
rect 9569 17234 9635 17237
rect 23921 17234 23987 17237
rect 9569 17232 23987 17234
rect 9569 17176 9574 17232
rect 9630 17176 23926 17232
rect 23982 17176 23987 17232
rect 9569 17174 23987 17176
rect 9569 17171 9635 17174
rect 23921 17171 23987 17174
rect 8097 17098 8163 17101
rect 16745 17098 16811 17101
rect 24614 17098 24674 17310
rect 27232 17280 27712 17310
rect 8097 17096 16811 17098
rect 8097 17040 8102 17096
rect 8158 17040 16750 17096
rect 16806 17040 16811 17096
rect 8097 17038 16811 17040
rect 8097 17035 8163 17038
rect 16745 17035 16811 17038
rect 16886 17038 24674 17098
rect 9989 16896 10309 16897
rect 9989 16832 9997 16896
rect 10061 16832 10077 16896
rect 10141 16832 10157 16896
rect 10221 16832 10237 16896
rect 10301 16832 10309 16896
rect 9989 16831 10309 16832
rect 9477 16690 9543 16693
rect 16886 16690 16946 17038
rect 19322 16896 19642 16897
rect 19322 16832 19330 16896
rect 19394 16832 19410 16896
rect 19474 16832 19490 16896
rect 19554 16832 19570 16896
rect 19634 16832 19642 16896
rect 19322 16831 19642 16832
rect 9477 16688 16946 16690
rect 9477 16632 9482 16688
rect 9538 16632 16946 16688
rect 9477 16630 16946 16632
rect 19689 16690 19755 16693
rect 27232 16690 27712 16720
rect 19689 16688 27712 16690
rect 19689 16632 19694 16688
rect 19750 16632 27712 16688
rect 19689 16630 27712 16632
rect 9477 16627 9543 16630
rect 19689 16627 19755 16630
rect 27232 16600 27712 16630
rect 5322 16352 5642 16353
rect 5322 16288 5330 16352
rect 5394 16288 5410 16352
rect 5474 16288 5490 16352
rect 5554 16288 5570 16352
rect 5634 16288 5642 16352
rect 5322 16287 5642 16288
rect 14656 16352 14976 16353
rect 14656 16288 14664 16352
rect 14728 16288 14744 16352
rect 14808 16288 14824 16352
rect 14888 16288 14904 16352
rect 14968 16288 14976 16352
rect 14656 16287 14976 16288
rect 23989 16352 24309 16353
rect 23989 16288 23997 16352
rect 24061 16288 24077 16352
rect 24141 16288 24157 16352
rect 24221 16288 24237 16352
rect 24301 16288 24309 16352
rect 23989 16287 24309 16288
rect 27232 16010 27712 16040
rect 27190 15920 27712 16010
rect 9989 15808 10309 15809
rect 9989 15744 9997 15808
rect 10061 15744 10077 15808
rect 10141 15744 10157 15808
rect 10221 15744 10237 15808
rect 10301 15744 10309 15808
rect 9989 15743 10309 15744
rect 19322 15808 19642 15809
rect 19322 15744 19330 15808
rect 19394 15744 19410 15808
rect 19474 15744 19490 15808
rect 19554 15744 19570 15808
rect 19634 15744 19642 15808
rect 19322 15743 19642 15744
rect 21713 15602 21779 15605
rect 27190 15602 27250 15920
rect 21713 15600 27250 15602
rect 21713 15544 21718 15600
rect 21774 15544 27250 15600
rect 21713 15542 27250 15544
rect 21713 15539 21779 15542
rect 10857 15466 10923 15469
rect 17941 15466 18007 15469
rect 10857 15464 16946 15466
rect 10857 15408 10862 15464
rect 10918 15408 16946 15464
rect 10857 15406 16946 15408
rect 10857 15403 10923 15406
rect 16886 15330 16946 15406
rect 17941 15464 24674 15466
rect 17941 15408 17946 15464
rect 18002 15408 24674 15464
rect 17941 15406 24674 15408
rect 17941 15403 18007 15406
rect 21713 15330 21779 15333
rect 16886 15328 21779 15330
rect 16886 15272 21718 15328
rect 21774 15272 21779 15328
rect 16886 15270 21779 15272
rect 24614 15330 24674 15406
rect 27232 15330 27712 15360
rect 24614 15270 27712 15330
rect 21713 15267 21779 15270
rect 5322 15264 5642 15265
rect 5322 15200 5330 15264
rect 5394 15200 5410 15264
rect 5474 15200 5490 15264
rect 5554 15200 5570 15264
rect 5634 15200 5642 15264
rect 5322 15199 5642 15200
rect 14656 15264 14976 15265
rect 14656 15200 14664 15264
rect 14728 15200 14744 15264
rect 14808 15200 14824 15264
rect 14888 15200 14904 15264
rect 14968 15200 14976 15264
rect 14656 15199 14976 15200
rect 23989 15264 24309 15265
rect 23989 15200 23997 15264
rect 24061 15200 24077 15264
rect 24141 15200 24157 15264
rect 24221 15200 24237 15264
rect 24301 15200 24309 15264
rect 27232 15240 27712 15270
rect 23989 15199 24309 15200
rect 8005 15194 8071 15197
rect 9845 15194 9911 15197
rect 8005 15192 9911 15194
rect 8005 15136 8010 15192
rect 8066 15136 9850 15192
rect 9906 15136 9911 15192
rect 8005 15134 9911 15136
rect 8005 15131 8071 15134
rect 9845 15131 9911 15134
rect 9989 14720 10309 14721
rect 9989 14656 9997 14720
rect 10061 14656 10077 14720
rect 10141 14656 10157 14720
rect 10221 14656 10237 14720
rect 10301 14656 10309 14720
rect 9989 14655 10309 14656
rect 19322 14720 19642 14721
rect 19322 14656 19330 14720
rect 19394 14656 19410 14720
rect 19474 14656 19490 14720
rect 19554 14656 19570 14720
rect 19634 14656 19642 14720
rect 19322 14655 19642 14656
rect 23829 14650 23895 14653
rect 27232 14650 27712 14680
rect 23829 14648 27712 14650
rect 23829 14592 23834 14648
rect 23890 14592 27712 14648
rect 23829 14590 27712 14592
rect 23829 14587 23895 14590
rect 27232 14560 27712 14590
rect 5322 14176 5642 14177
rect 5322 14112 5330 14176
rect 5394 14112 5410 14176
rect 5474 14112 5490 14176
rect 5554 14112 5570 14176
rect 5634 14112 5642 14176
rect 5322 14111 5642 14112
rect 14656 14176 14976 14177
rect 14656 14112 14664 14176
rect 14728 14112 14744 14176
rect 14808 14112 14824 14176
rect 14888 14112 14904 14176
rect 14968 14112 14976 14176
rect 14656 14111 14976 14112
rect 23989 14176 24309 14177
rect 23989 14112 23997 14176
rect 24061 14112 24077 14176
rect 24141 14112 24157 14176
rect 24221 14112 24237 14176
rect 24301 14112 24309 14176
rect 23989 14111 24309 14112
rect 15457 13970 15523 13973
rect 27232 13970 27712 14000
rect 15457 13968 27712 13970
rect 15457 13912 15462 13968
rect 15518 13912 27712 13968
rect 15457 13910 27712 13912
rect 15457 13907 15523 13910
rect 27232 13880 27712 13910
rect 4325 13834 4391 13837
rect 12421 13834 12487 13837
rect 12789 13834 12855 13837
rect 4325 13832 12855 13834
rect 4325 13776 4330 13832
rect 4386 13776 12426 13832
rect 12482 13776 12794 13832
rect 12850 13776 12855 13832
rect 4325 13774 12855 13776
rect 4325 13771 4391 13774
rect 12421 13771 12487 13774
rect 12789 13771 12855 13774
rect 9989 13632 10309 13633
rect 9989 13568 9997 13632
rect 10061 13568 10077 13632
rect 10141 13568 10157 13632
rect 10221 13568 10237 13632
rect 10301 13568 10309 13632
rect 9989 13567 10309 13568
rect 19322 13632 19642 13633
rect 19322 13568 19330 13632
rect 19394 13568 19410 13632
rect 19474 13568 19490 13632
rect 19554 13568 19570 13632
rect 19634 13568 19642 13632
rect 19322 13567 19642 13568
rect 24473 13290 24539 13293
rect 27232 13290 27712 13320
rect 24473 13288 27712 13290
rect 24473 13232 24478 13288
rect 24534 13232 27712 13288
rect 24473 13230 27712 13232
rect 24473 13227 24539 13230
rect 27232 13200 27712 13230
rect 5322 13088 5642 13089
rect 5322 13024 5330 13088
rect 5394 13024 5410 13088
rect 5474 13024 5490 13088
rect 5554 13024 5570 13088
rect 5634 13024 5642 13088
rect 5322 13023 5642 13024
rect 14656 13088 14976 13089
rect 14656 13024 14664 13088
rect 14728 13024 14744 13088
rect 14808 13024 14824 13088
rect 14888 13024 14904 13088
rect 14968 13024 14976 13088
rect 14656 13023 14976 13024
rect 23989 13088 24309 13089
rect 23989 13024 23997 13088
rect 24061 13024 24077 13088
rect 24141 13024 24157 13088
rect 24221 13024 24237 13088
rect 24301 13024 24309 13088
rect 23989 13023 24309 13024
rect 23829 13018 23895 13021
rect 22590 13016 23895 13018
rect 22590 12960 23834 13016
rect 23890 12960 23895 13016
rect 22590 12958 23895 12960
rect 12329 12746 12395 12749
rect 22590 12746 22650 12958
rect 23829 12955 23895 12958
rect 23553 12746 23619 12749
rect 12329 12744 22650 12746
rect 12329 12688 12334 12744
rect 12390 12688 22650 12744
rect 12329 12686 22650 12688
rect 22774 12744 23619 12746
rect 22774 12688 23558 12744
rect 23614 12688 23619 12744
rect 22774 12686 23619 12688
rect 12329 12683 12395 12686
rect 21713 12610 21779 12613
rect 22774 12610 22834 12686
rect 23553 12683 23619 12686
rect 21713 12608 22834 12610
rect 21713 12552 21718 12608
rect 21774 12552 22834 12608
rect 21713 12550 22834 12552
rect 23185 12610 23251 12613
rect 27232 12610 27712 12640
rect 23185 12608 27712 12610
rect 23185 12552 23190 12608
rect 23246 12552 27712 12608
rect 23185 12550 27712 12552
rect 21713 12547 21779 12550
rect 23185 12547 23251 12550
rect 9989 12544 10309 12545
rect 9989 12480 9997 12544
rect 10061 12480 10077 12544
rect 10141 12480 10157 12544
rect 10221 12480 10237 12544
rect 10301 12480 10309 12544
rect 9989 12479 10309 12480
rect 19322 12544 19642 12545
rect 19322 12480 19330 12544
rect 19394 12480 19410 12544
rect 19474 12480 19490 12544
rect 19554 12480 19570 12544
rect 19634 12480 19642 12544
rect 27232 12520 27712 12550
rect 19322 12479 19642 12480
rect 5322 12000 5642 12001
rect 5322 11936 5330 12000
rect 5394 11936 5410 12000
rect 5474 11936 5490 12000
rect 5554 11936 5570 12000
rect 5634 11936 5642 12000
rect 5322 11935 5642 11936
rect 14656 12000 14976 12001
rect 14656 11936 14664 12000
rect 14728 11936 14744 12000
rect 14808 11936 14824 12000
rect 14888 11936 14904 12000
rect 14968 11936 14976 12000
rect 14656 11935 14976 11936
rect 23989 12000 24309 12001
rect 23989 11936 23997 12000
rect 24061 11936 24077 12000
rect 24141 11936 24157 12000
rect 24221 11936 24237 12000
rect 24301 11936 24309 12000
rect 23989 11935 24309 11936
rect 27232 11930 27712 11960
rect 24430 11870 27712 11930
rect 23737 11794 23803 11797
rect 24430 11794 24490 11870
rect 27232 11840 27712 11870
rect 23737 11792 24490 11794
rect 23737 11736 23742 11792
rect 23798 11736 24490 11792
rect 23737 11734 24490 11736
rect 23737 11731 23803 11734
rect 10765 11522 10831 11525
rect 14537 11522 14603 11525
rect 10765 11520 14603 11522
rect 10765 11464 10770 11520
rect 10826 11464 14542 11520
rect 14598 11464 14603 11520
rect 10765 11462 14603 11464
rect 10765 11459 10831 11462
rect 14537 11459 14603 11462
rect 9989 11456 10309 11457
rect 9989 11392 9997 11456
rect 10061 11392 10077 11456
rect 10141 11392 10157 11456
rect 10221 11392 10237 11456
rect 10301 11392 10309 11456
rect 9989 11391 10309 11392
rect 19322 11456 19642 11457
rect 19322 11392 19330 11456
rect 19394 11392 19410 11456
rect 19474 11392 19490 11456
rect 19554 11392 19570 11456
rect 19634 11392 19642 11456
rect 19322 11391 19642 11392
rect 9385 11250 9451 11253
rect 17481 11250 17547 11253
rect 27232 11250 27712 11280
rect 9385 11248 17547 11250
rect 9385 11192 9390 11248
rect 9446 11192 17486 11248
rect 17542 11192 17547 11248
rect 9385 11190 17547 11192
rect 9385 11187 9451 11190
rect 17481 11187 17547 11190
rect 23694 11190 27712 11250
rect 21069 10978 21135 10981
rect 23694 10978 23754 11190
rect 27232 11160 27712 11190
rect 21069 10976 23754 10978
rect 21069 10920 21074 10976
rect 21130 10920 23754 10976
rect 21069 10918 23754 10920
rect 21069 10915 21135 10918
rect 5322 10912 5642 10913
rect 5322 10848 5330 10912
rect 5394 10848 5410 10912
rect 5474 10848 5490 10912
rect 5554 10848 5570 10912
rect 5634 10848 5642 10912
rect 5322 10847 5642 10848
rect 14656 10912 14976 10913
rect 14656 10848 14664 10912
rect 14728 10848 14744 10912
rect 14808 10848 14824 10912
rect 14888 10848 14904 10912
rect 14968 10848 14976 10912
rect 14656 10847 14976 10848
rect 23989 10912 24309 10913
rect 23989 10848 23997 10912
rect 24061 10848 24077 10912
rect 24141 10848 24157 10912
rect 24221 10848 24237 10912
rect 24301 10848 24309 10912
rect 23989 10847 24309 10848
rect 15273 10570 15339 10573
rect 23737 10570 23803 10573
rect 15273 10568 23803 10570
rect 15273 10512 15278 10568
rect 15334 10512 23742 10568
rect 23798 10512 23803 10568
rect 15273 10510 23803 10512
rect 15273 10507 15339 10510
rect 23737 10507 23803 10510
rect 23921 10570 23987 10573
rect 27232 10570 27712 10600
rect 23921 10568 27712 10570
rect 23921 10512 23926 10568
rect 23982 10512 27712 10568
rect 23921 10510 27712 10512
rect 23921 10507 23987 10510
rect 27232 10480 27712 10510
rect 9989 10368 10309 10369
rect 9989 10304 9997 10368
rect 10061 10304 10077 10368
rect 10141 10304 10157 10368
rect 10221 10304 10237 10368
rect 10301 10304 10309 10368
rect 9989 10303 10309 10304
rect 19322 10368 19642 10369
rect 19322 10304 19330 10368
rect 19394 10304 19410 10368
rect 19474 10304 19490 10368
rect 19554 10304 19570 10368
rect 19634 10304 19642 10368
rect 19322 10303 19642 10304
rect 24473 10162 24539 10165
rect 27233 10162 27299 10165
rect 24473 10160 27299 10162
rect 24473 10104 24478 10160
rect 24534 10104 27238 10160
rect 27294 10104 27299 10160
rect 24473 10102 27299 10104
rect 24473 10099 24539 10102
rect 27233 10099 27299 10102
rect 23185 10026 23251 10029
rect 23185 10024 24490 10026
rect 23185 9968 23190 10024
rect 23246 9968 24490 10024
rect 23185 9966 24490 9968
rect 23185 9963 23251 9966
rect 24430 9890 24490 9966
rect 27232 9890 27712 9920
rect 24430 9830 27712 9890
rect 5322 9824 5642 9825
rect 5322 9760 5330 9824
rect 5394 9760 5410 9824
rect 5474 9760 5490 9824
rect 5554 9760 5570 9824
rect 5634 9760 5642 9824
rect 5322 9759 5642 9760
rect 14656 9824 14976 9825
rect 14656 9760 14664 9824
rect 14728 9760 14744 9824
rect 14808 9760 14824 9824
rect 14888 9760 14904 9824
rect 14968 9760 14976 9824
rect 14656 9759 14976 9760
rect 23989 9824 24309 9825
rect 23989 9760 23997 9824
rect 24061 9760 24077 9824
rect 24141 9760 24157 9824
rect 24221 9760 24237 9824
rect 24301 9760 24309 9824
rect 27232 9800 27712 9830
rect 23989 9759 24309 9760
rect 18953 9754 19019 9757
rect 20609 9754 20675 9757
rect 18953 9752 20675 9754
rect 18953 9696 18958 9752
rect 19014 9696 20614 9752
rect 20670 9696 20675 9752
rect 18953 9694 20675 9696
rect 18953 9691 19019 9694
rect 20609 9691 20675 9694
rect 14905 9618 14971 9621
rect 18861 9618 18927 9621
rect 14905 9616 18927 9618
rect 14905 9560 14910 9616
rect 14966 9560 18866 9616
rect 18922 9560 18927 9616
rect 14905 9558 18927 9560
rect 14905 9555 14971 9558
rect 18861 9555 18927 9558
rect 9989 9280 10309 9281
rect 9989 9216 9997 9280
rect 10061 9216 10077 9280
rect 10141 9216 10157 9280
rect 10221 9216 10237 9280
rect 10301 9216 10309 9280
rect 9989 9215 10309 9216
rect 19322 9280 19642 9281
rect 19322 9216 19330 9280
rect 19394 9216 19410 9280
rect 19474 9216 19490 9280
rect 19554 9216 19570 9280
rect 19634 9216 19642 9280
rect 19322 9215 19642 9216
rect 27232 9210 27712 9240
rect 19784 9150 27712 9210
rect 18401 9074 18467 9077
rect 19784 9074 19844 9150
rect 27232 9120 27712 9150
rect 18401 9072 19844 9074
rect 18401 9016 18406 9072
rect 18462 9016 19844 9072
rect 18401 9014 19844 9016
rect 18401 9011 18467 9014
rect 5322 8736 5642 8737
rect 5322 8672 5330 8736
rect 5394 8672 5410 8736
rect 5474 8672 5490 8736
rect 5554 8672 5570 8736
rect 5634 8672 5642 8736
rect 5322 8671 5642 8672
rect 14656 8736 14976 8737
rect 14656 8672 14664 8736
rect 14728 8672 14744 8736
rect 14808 8672 14824 8736
rect 14888 8672 14904 8736
rect 14968 8672 14976 8736
rect 14656 8671 14976 8672
rect 23989 8736 24309 8737
rect 23989 8672 23997 8736
rect 24061 8672 24077 8736
rect 24141 8672 24157 8736
rect 24221 8672 24237 8736
rect 24301 8672 24309 8736
rect 23989 8671 24309 8672
rect 16009 8530 16075 8533
rect 23921 8530 23987 8533
rect 27232 8530 27712 8560
rect 16009 8528 23987 8530
rect 16009 8472 16014 8528
rect 16070 8472 23926 8528
rect 23982 8472 23987 8528
rect 16009 8470 23987 8472
rect 16009 8467 16075 8470
rect 23921 8467 23987 8470
rect 24430 8470 27712 8530
rect 9989 8192 10309 8193
rect 9989 8128 9997 8192
rect 10061 8128 10077 8192
rect 10141 8128 10157 8192
rect 10221 8128 10237 8192
rect 10301 8128 10309 8192
rect 9989 8127 10309 8128
rect 19322 8192 19642 8193
rect 19322 8128 19330 8192
rect 19394 8128 19410 8192
rect 19474 8128 19490 8192
rect 19554 8128 19570 8192
rect 19634 8128 19642 8192
rect 19322 8127 19642 8128
rect 17849 7986 17915 7989
rect 24430 7986 24490 8470
rect 27232 8440 27712 8470
rect 17849 7984 24490 7986
rect 17849 7928 17854 7984
rect 17910 7928 24490 7984
rect 17849 7926 24490 7928
rect 17849 7923 17915 7926
rect 24473 7850 24539 7853
rect 27232 7850 27712 7880
rect 24473 7848 27712 7850
rect 24473 7792 24478 7848
rect 24534 7792 27712 7848
rect 24473 7790 27712 7792
rect 24473 7787 24539 7790
rect 27232 7760 27712 7790
rect 5322 7648 5642 7649
rect 5322 7584 5330 7648
rect 5394 7584 5410 7648
rect 5474 7584 5490 7648
rect 5554 7584 5570 7648
rect 5634 7584 5642 7648
rect 5322 7583 5642 7584
rect 14656 7648 14976 7649
rect 14656 7584 14664 7648
rect 14728 7584 14744 7648
rect 14808 7584 14824 7648
rect 14888 7584 14904 7648
rect 14968 7584 14976 7648
rect 14656 7583 14976 7584
rect 23989 7648 24309 7649
rect 23989 7584 23997 7648
rect 24061 7584 24077 7648
rect 24141 7584 24157 7648
rect 24221 7584 24237 7648
rect 24301 7584 24309 7648
rect 23989 7583 24309 7584
rect 27232 7170 27712 7200
rect 24246 7110 27712 7170
rect 9989 7104 10309 7105
rect 9989 7040 9997 7104
rect 10061 7040 10077 7104
rect 10141 7040 10157 7104
rect 10221 7040 10237 7104
rect 10301 7040 10309 7104
rect 9989 7039 10309 7040
rect 19322 7104 19642 7105
rect 19322 7040 19330 7104
rect 19394 7040 19410 7104
rect 19474 7040 19490 7104
rect 19554 7040 19570 7104
rect 19634 7040 19642 7104
rect 19322 7039 19642 7040
rect 19689 6898 19755 6901
rect 24246 6898 24306 7110
rect 27232 7080 27712 7110
rect 19689 6896 24306 6898
rect 19689 6840 19694 6896
rect 19750 6840 24306 6896
rect 19689 6838 24306 6840
rect 19689 6835 19755 6838
rect 5322 6560 5642 6561
rect 5322 6496 5330 6560
rect 5394 6496 5410 6560
rect 5474 6496 5490 6560
rect 5554 6496 5570 6560
rect 5634 6496 5642 6560
rect 5322 6495 5642 6496
rect 14656 6560 14976 6561
rect 14656 6496 14664 6560
rect 14728 6496 14744 6560
rect 14808 6496 14824 6560
rect 14888 6496 14904 6560
rect 14968 6496 14976 6560
rect 14656 6495 14976 6496
rect 23989 6560 24309 6561
rect 23989 6496 23997 6560
rect 24061 6496 24077 6560
rect 24141 6496 24157 6560
rect 24221 6496 24237 6560
rect 24301 6496 24309 6560
rect 23989 6495 24309 6496
rect 24381 6490 24447 6493
rect 27232 6490 27712 6520
rect 24381 6488 27712 6490
rect 24381 6432 24386 6488
rect 24442 6432 27712 6488
rect 24381 6430 27712 6432
rect 24381 6427 24447 6430
rect 27232 6400 27712 6430
rect 19229 6354 19295 6357
rect 24473 6354 24539 6357
rect 19229 6352 24539 6354
rect 19229 6296 19234 6352
rect 19290 6296 24478 6352
rect 24534 6296 24539 6352
rect 19229 6294 24539 6296
rect 19229 6291 19295 6294
rect 24473 6291 24539 6294
rect 9989 6016 10309 6017
rect 9989 5952 9997 6016
rect 10061 5952 10077 6016
rect 10141 5952 10157 6016
rect 10221 5952 10237 6016
rect 10301 5952 10309 6016
rect 9989 5951 10309 5952
rect 19322 6016 19642 6017
rect 19322 5952 19330 6016
rect 19394 5952 19410 6016
rect 19474 5952 19490 6016
rect 19554 5952 19570 6016
rect 19634 5952 19642 6016
rect 19322 5951 19642 5952
rect 21529 5810 21595 5813
rect 27232 5810 27712 5840
rect 21529 5808 27712 5810
rect 21529 5752 21534 5808
rect 21590 5752 27712 5808
rect 21529 5750 27712 5752
rect 21529 5747 21595 5750
rect 27232 5720 27712 5750
rect 5322 5472 5642 5473
rect 5322 5408 5330 5472
rect 5394 5408 5410 5472
rect 5474 5408 5490 5472
rect 5554 5408 5570 5472
rect 5634 5408 5642 5472
rect 5322 5407 5642 5408
rect 14656 5472 14976 5473
rect 14656 5408 14664 5472
rect 14728 5408 14744 5472
rect 14808 5408 14824 5472
rect 14888 5408 14904 5472
rect 14968 5408 14976 5472
rect 14656 5407 14976 5408
rect 23989 5472 24309 5473
rect 23989 5408 23997 5472
rect 24061 5408 24077 5472
rect 24141 5408 24157 5472
rect 24221 5408 24237 5472
rect 24301 5408 24309 5472
rect 23989 5407 24309 5408
rect 24289 5130 24355 5133
rect 27232 5130 27712 5160
rect 24289 5128 27712 5130
rect 24289 5072 24294 5128
rect 24350 5072 27712 5128
rect 24289 5070 27712 5072
rect 24289 5067 24355 5070
rect 27232 5040 27712 5070
rect 9989 4928 10309 4929
rect 9989 4864 9997 4928
rect 10061 4864 10077 4928
rect 10141 4864 10157 4928
rect 10221 4864 10237 4928
rect 10301 4864 10309 4928
rect 9989 4863 10309 4864
rect 19322 4928 19642 4929
rect 19322 4864 19330 4928
rect 19394 4864 19410 4928
rect 19474 4864 19490 4928
rect 19554 4864 19570 4928
rect 19634 4864 19642 4928
rect 19322 4863 19642 4864
rect 20149 4722 20215 4725
rect 21437 4722 21503 4725
rect 20149 4720 24674 4722
rect 20149 4664 20154 4720
rect 20210 4664 21442 4720
rect 21498 4664 24674 4720
rect 20149 4662 24674 4664
rect 20149 4659 20215 4662
rect 21437 4659 21503 4662
rect 24614 4450 24674 4662
rect 27232 4450 27712 4480
rect 24614 4390 27712 4450
rect 5322 4384 5642 4385
rect 5322 4320 5330 4384
rect 5394 4320 5410 4384
rect 5474 4320 5490 4384
rect 5554 4320 5570 4384
rect 5634 4320 5642 4384
rect 5322 4319 5642 4320
rect 14656 4384 14976 4385
rect 14656 4320 14664 4384
rect 14728 4320 14744 4384
rect 14808 4320 14824 4384
rect 14888 4320 14904 4384
rect 14968 4320 14976 4384
rect 14656 4319 14976 4320
rect 23989 4384 24309 4385
rect 23989 4320 23997 4384
rect 24061 4320 24077 4384
rect 24141 4320 24157 4384
rect 24221 4320 24237 4384
rect 24301 4320 24309 4384
rect 27232 4360 27712 4390
rect 23989 4319 24309 4320
rect 21621 4178 21687 4181
rect 24473 4178 24539 4181
rect 21621 4176 24539 4178
rect 21621 4120 21626 4176
rect 21682 4120 24478 4176
rect 24534 4120 24539 4176
rect 21621 4118 24539 4120
rect 21621 4115 21687 4118
rect 24473 4115 24539 4118
rect 645 4042 711 4045
rect 11041 4042 11107 4045
rect 645 4040 11107 4042
rect 645 3984 650 4040
rect 706 3984 11046 4040
rect 11102 3984 11107 4040
rect 645 3982 11107 3984
rect 645 3979 711 3982
rect 11041 3979 11107 3982
rect 9989 3840 10309 3841
rect 9989 3776 9997 3840
rect 10061 3776 10077 3840
rect 10141 3776 10157 3840
rect 10221 3776 10237 3840
rect 10301 3776 10309 3840
rect 9989 3775 10309 3776
rect 19322 3840 19642 3841
rect 19322 3776 19330 3840
rect 19394 3776 19410 3840
rect 19474 3776 19490 3840
rect 19554 3776 19570 3840
rect 19634 3776 19642 3840
rect 19322 3775 19642 3776
rect 27232 3770 27712 3800
rect 26822 3710 27712 3770
rect 4693 3634 4759 3637
rect 18769 3634 18835 3637
rect 4693 3632 18835 3634
rect 4693 3576 4698 3632
rect 4754 3576 18774 3632
rect 18830 3576 18835 3632
rect 4693 3574 18835 3576
rect 4693 3571 4759 3574
rect 18769 3571 18835 3574
rect 1 3498 67 3501
rect 20977 3498 21043 3501
rect 1 3496 21043 3498
rect 1 3440 6 3496
rect 62 3440 20982 3496
rect 21038 3440 21043 3496
rect 1 3438 21043 3440
rect 1 3435 67 3438
rect 20977 3435 21043 3438
rect 24473 3362 24539 3365
rect 26589 3362 26655 3365
rect 24473 3360 26655 3362
rect 24473 3304 24478 3360
rect 24534 3304 26594 3360
rect 26650 3304 26655 3360
rect 24473 3302 26655 3304
rect 24473 3299 24539 3302
rect 26589 3299 26655 3302
rect 5322 3296 5642 3297
rect 5322 3232 5330 3296
rect 5394 3232 5410 3296
rect 5474 3232 5490 3296
rect 5554 3232 5570 3296
rect 5634 3232 5642 3296
rect 5322 3231 5642 3232
rect 14656 3296 14976 3297
rect 14656 3232 14664 3296
rect 14728 3232 14744 3296
rect 14808 3232 14824 3296
rect 14888 3232 14904 3296
rect 14968 3232 14976 3296
rect 14656 3231 14976 3232
rect 23989 3296 24309 3297
rect 23989 3232 23997 3296
rect 24061 3232 24077 3296
rect 24141 3232 24157 3296
rect 24221 3232 24237 3296
rect 24301 3232 24309 3296
rect 23989 3231 24309 3232
rect 24473 3226 24539 3229
rect 26822 3226 26882 3710
rect 27232 3680 27712 3710
rect 24473 3224 26882 3226
rect 24473 3168 24478 3224
rect 24534 3168 26882 3224
rect 24473 3166 26882 3168
rect 24473 3163 24539 3166
rect 1289 3090 1355 3093
rect 10489 3090 10555 3093
rect 1289 3088 10555 3090
rect 1289 3032 1294 3088
rect 1350 3032 10494 3088
rect 10550 3032 10555 3088
rect 1289 3030 10555 3032
rect 1289 3027 1355 3030
rect 10489 3027 10555 3030
rect 23645 3090 23711 3093
rect 27232 3090 27712 3120
rect 23645 3088 27712 3090
rect 23645 3032 23650 3088
rect 23706 3032 27712 3088
rect 23645 3030 27712 3032
rect 23645 3027 23711 3030
rect 27232 3000 27712 3030
rect 22725 2954 22791 2957
rect 25853 2954 25919 2957
rect 22725 2952 25919 2954
rect 22725 2896 22730 2952
rect 22786 2896 25858 2952
rect 25914 2896 25919 2952
rect 22725 2894 25919 2896
rect 22725 2891 22791 2894
rect 25853 2891 25919 2894
rect 25301 2818 25367 2821
rect 25301 2816 25410 2818
rect 25301 2760 25306 2816
rect 25362 2760 25410 2816
rect 25301 2755 25410 2760
rect 9989 2752 10309 2753
rect 9989 2688 9997 2752
rect 10061 2688 10077 2752
rect 10141 2688 10157 2752
rect 10221 2688 10237 2752
rect 10301 2688 10309 2752
rect 9989 2687 10309 2688
rect 19322 2752 19642 2753
rect 19322 2688 19330 2752
rect 19394 2688 19410 2752
rect 19474 2688 19490 2752
rect 19554 2688 19570 2752
rect 19634 2688 19642 2752
rect 19322 2687 19642 2688
rect 25350 2682 25410 2755
rect 25350 2622 25594 2682
rect 25534 2410 25594 2622
rect 27232 2410 27712 2440
rect 25534 2350 27712 2410
rect 27232 2320 27712 2350
rect 5322 2208 5642 2209
rect 5322 2144 5330 2208
rect 5394 2144 5410 2208
rect 5474 2144 5490 2208
rect 5554 2144 5570 2208
rect 5634 2144 5642 2208
rect 5322 2143 5642 2144
rect 14656 2208 14976 2209
rect 14656 2144 14664 2208
rect 14728 2144 14744 2208
rect 14808 2144 14824 2208
rect 14888 2144 14904 2208
rect 14968 2144 14976 2208
rect 14656 2143 14976 2144
rect 23989 2208 24309 2209
rect 23989 2144 23997 2208
rect 24061 2144 24077 2208
rect 24141 2144 24157 2208
rect 24221 2144 24237 2208
rect 24301 2144 24309 2208
rect 23989 2143 24309 2144
rect 24381 1730 24447 1733
rect 27232 1730 27712 1760
rect 24381 1728 27712 1730
rect 24381 1672 24386 1728
rect 24442 1672 27712 1728
rect 24381 1670 27712 1672
rect 24381 1667 24447 1670
rect 27232 1640 27712 1670
rect 23277 1050 23343 1053
rect 27232 1050 27712 1080
rect 23277 1048 27712 1050
rect 23277 992 23282 1048
rect 23338 992 27712 1048
rect 23277 990 27712 992
rect 23277 987 23343 990
rect 27232 960 27712 990
rect 23921 370 23987 373
rect 27232 370 27712 400
rect 23921 368 27712 370
rect 23921 312 23926 368
rect 23982 312 27712 368
rect 23921 310 27712 312
rect 23921 307 23987 310
rect 27232 280 27712 310
<< via3 >>
rect 9997 25596 10061 25600
rect 9997 25540 10001 25596
rect 10001 25540 10057 25596
rect 10057 25540 10061 25596
rect 9997 25536 10061 25540
rect 10077 25596 10141 25600
rect 10077 25540 10081 25596
rect 10081 25540 10137 25596
rect 10137 25540 10141 25596
rect 10077 25536 10141 25540
rect 10157 25596 10221 25600
rect 10157 25540 10161 25596
rect 10161 25540 10217 25596
rect 10217 25540 10221 25596
rect 10157 25536 10221 25540
rect 10237 25596 10301 25600
rect 10237 25540 10241 25596
rect 10241 25540 10297 25596
rect 10297 25540 10301 25596
rect 10237 25536 10301 25540
rect 19330 25596 19394 25600
rect 19330 25540 19334 25596
rect 19334 25540 19390 25596
rect 19390 25540 19394 25596
rect 19330 25536 19394 25540
rect 19410 25596 19474 25600
rect 19410 25540 19414 25596
rect 19414 25540 19470 25596
rect 19470 25540 19474 25596
rect 19410 25536 19474 25540
rect 19490 25596 19554 25600
rect 19490 25540 19494 25596
rect 19494 25540 19550 25596
rect 19550 25540 19554 25596
rect 19490 25536 19554 25540
rect 19570 25596 19634 25600
rect 19570 25540 19574 25596
rect 19574 25540 19630 25596
rect 19630 25540 19634 25596
rect 19570 25536 19634 25540
rect 5330 25052 5394 25056
rect 5330 24996 5334 25052
rect 5334 24996 5390 25052
rect 5390 24996 5394 25052
rect 5330 24992 5394 24996
rect 5410 25052 5474 25056
rect 5410 24996 5414 25052
rect 5414 24996 5470 25052
rect 5470 24996 5474 25052
rect 5410 24992 5474 24996
rect 5490 25052 5554 25056
rect 5490 24996 5494 25052
rect 5494 24996 5550 25052
rect 5550 24996 5554 25052
rect 5490 24992 5554 24996
rect 5570 25052 5634 25056
rect 5570 24996 5574 25052
rect 5574 24996 5630 25052
rect 5630 24996 5634 25052
rect 5570 24992 5634 24996
rect 14664 25052 14728 25056
rect 14664 24996 14668 25052
rect 14668 24996 14724 25052
rect 14724 24996 14728 25052
rect 14664 24992 14728 24996
rect 14744 25052 14808 25056
rect 14744 24996 14748 25052
rect 14748 24996 14804 25052
rect 14804 24996 14808 25052
rect 14744 24992 14808 24996
rect 14824 25052 14888 25056
rect 14824 24996 14828 25052
rect 14828 24996 14884 25052
rect 14884 24996 14888 25052
rect 14824 24992 14888 24996
rect 14904 25052 14968 25056
rect 14904 24996 14908 25052
rect 14908 24996 14964 25052
rect 14964 24996 14968 25052
rect 14904 24992 14968 24996
rect 23997 25052 24061 25056
rect 23997 24996 24001 25052
rect 24001 24996 24057 25052
rect 24057 24996 24061 25052
rect 23997 24992 24061 24996
rect 24077 25052 24141 25056
rect 24077 24996 24081 25052
rect 24081 24996 24137 25052
rect 24137 24996 24141 25052
rect 24077 24992 24141 24996
rect 24157 25052 24221 25056
rect 24157 24996 24161 25052
rect 24161 24996 24217 25052
rect 24217 24996 24221 25052
rect 24157 24992 24221 24996
rect 24237 25052 24301 25056
rect 24237 24996 24241 25052
rect 24241 24996 24297 25052
rect 24297 24996 24301 25052
rect 24237 24992 24301 24996
rect 9997 24508 10061 24512
rect 9997 24452 10001 24508
rect 10001 24452 10057 24508
rect 10057 24452 10061 24508
rect 9997 24448 10061 24452
rect 10077 24508 10141 24512
rect 10077 24452 10081 24508
rect 10081 24452 10137 24508
rect 10137 24452 10141 24508
rect 10077 24448 10141 24452
rect 10157 24508 10221 24512
rect 10157 24452 10161 24508
rect 10161 24452 10217 24508
rect 10217 24452 10221 24508
rect 10157 24448 10221 24452
rect 10237 24508 10301 24512
rect 10237 24452 10241 24508
rect 10241 24452 10297 24508
rect 10297 24452 10301 24508
rect 10237 24448 10301 24452
rect 19330 24508 19394 24512
rect 19330 24452 19334 24508
rect 19334 24452 19390 24508
rect 19390 24452 19394 24508
rect 19330 24448 19394 24452
rect 19410 24508 19474 24512
rect 19410 24452 19414 24508
rect 19414 24452 19470 24508
rect 19470 24452 19474 24508
rect 19410 24448 19474 24452
rect 19490 24508 19554 24512
rect 19490 24452 19494 24508
rect 19494 24452 19550 24508
rect 19550 24452 19554 24508
rect 19490 24448 19554 24452
rect 19570 24508 19634 24512
rect 19570 24452 19574 24508
rect 19574 24452 19630 24508
rect 19630 24452 19634 24508
rect 19570 24448 19634 24452
rect 5330 23964 5394 23968
rect 5330 23908 5334 23964
rect 5334 23908 5390 23964
rect 5390 23908 5394 23964
rect 5330 23904 5394 23908
rect 5410 23964 5474 23968
rect 5410 23908 5414 23964
rect 5414 23908 5470 23964
rect 5470 23908 5474 23964
rect 5410 23904 5474 23908
rect 5490 23964 5554 23968
rect 5490 23908 5494 23964
rect 5494 23908 5550 23964
rect 5550 23908 5554 23964
rect 5490 23904 5554 23908
rect 5570 23964 5634 23968
rect 5570 23908 5574 23964
rect 5574 23908 5630 23964
rect 5630 23908 5634 23964
rect 5570 23904 5634 23908
rect 14664 23964 14728 23968
rect 14664 23908 14668 23964
rect 14668 23908 14724 23964
rect 14724 23908 14728 23964
rect 14664 23904 14728 23908
rect 14744 23964 14808 23968
rect 14744 23908 14748 23964
rect 14748 23908 14804 23964
rect 14804 23908 14808 23964
rect 14744 23904 14808 23908
rect 14824 23964 14888 23968
rect 14824 23908 14828 23964
rect 14828 23908 14884 23964
rect 14884 23908 14888 23964
rect 14824 23904 14888 23908
rect 14904 23964 14968 23968
rect 14904 23908 14908 23964
rect 14908 23908 14964 23964
rect 14964 23908 14968 23964
rect 14904 23904 14968 23908
rect 23997 23964 24061 23968
rect 23997 23908 24001 23964
rect 24001 23908 24057 23964
rect 24057 23908 24061 23964
rect 23997 23904 24061 23908
rect 24077 23964 24141 23968
rect 24077 23908 24081 23964
rect 24081 23908 24137 23964
rect 24137 23908 24141 23964
rect 24077 23904 24141 23908
rect 24157 23964 24221 23968
rect 24157 23908 24161 23964
rect 24161 23908 24217 23964
rect 24217 23908 24221 23964
rect 24157 23904 24221 23908
rect 24237 23964 24301 23968
rect 24237 23908 24241 23964
rect 24241 23908 24297 23964
rect 24297 23908 24301 23964
rect 24237 23904 24301 23908
rect 9997 23420 10061 23424
rect 9997 23364 10001 23420
rect 10001 23364 10057 23420
rect 10057 23364 10061 23420
rect 9997 23360 10061 23364
rect 10077 23420 10141 23424
rect 10077 23364 10081 23420
rect 10081 23364 10137 23420
rect 10137 23364 10141 23420
rect 10077 23360 10141 23364
rect 10157 23420 10221 23424
rect 10157 23364 10161 23420
rect 10161 23364 10217 23420
rect 10217 23364 10221 23420
rect 10157 23360 10221 23364
rect 10237 23420 10301 23424
rect 10237 23364 10241 23420
rect 10241 23364 10297 23420
rect 10297 23364 10301 23420
rect 10237 23360 10301 23364
rect 19330 23420 19394 23424
rect 19330 23364 19334 23420
rect 19334 23364 19390 23420
rect 19390 23364 19394 23420
rect 19330 23360 19394 23364
rect 19410 23420 19474 23424
rect 19410 23364 19414 23420
rect 19414 23364 19470 23420
rect 19470 23364 19474 23420
rect 19410 23360 19474 23364
rect 19490 23420 19554 23424
rect 19490 23364 19494 23420
rect 19494 23364 19550 23420
rect 19550 23364 19554 23420
rect 19490 23360 19554 23364
rect 19570 23420 19634 23424
rect 19570 23364 19574 23420
rect 19574 23364 19630 23420
rect 19630 23364 19634 23420
rect 19570 23360 19634 23364
rect 5330 22876 5394 22880
rect 5330 22820 5334 22876
rect 5334 22820 5390 22876
rect 5390 22820 5394 22876
rect 5330 22816 5394 22820
rect 5410 22876 5474 22880
rect 5410 22820 5414 22876
rect 5414 22820 5470 22876
rect 5470 22820 5474 22876
rect 5410 22816 5474 22820
rect 5490 22876 5554 22880
rect 5490 22820 5494 22876
rect 5494 22820 5550 22876
rect 5550 22820 5554 22876
rect 5490 22816 5554 22820
rect 5570 22876 5634 22880
rect 5570 22820 5574 22876
rect 5574 22820 5630 22876
rect 5630 22820 5634 22876
rect 5570 22816 5634 22820
rect 14664 22876 14728 22880
rect 14664 22820 14668 22876
rect 14668 22820 14724 22876
rect 14724 22820 14728 22876
rect 14664 22816 14728 22820
rect 14744 22876 14808 22880
rect 14744 22820 14748 22876
rect 14748 22820 14804 22876
rect 14804 22820 14808 22876
rect 14744 22816 14808 22820
rect 14824 22876 14888 22880
rect 14824 22820 14828 22876
rect 14828 22820 14884 22876
rect 14884 22820 14888 22876
rect 14824 22816 14888 22820
rect 14904 22876 14968 22880
rect 14904 22820 14908 22876
rect 14908 22820 14964 22876
rect 14964 22820 14968 22876
rect 14904 22816 14968 22820
rect 23997 22876 24061 22880
rect 23997 22820 24001 22876
rect 24001 22820 24057 22876
rect 24057 22820 24061 22876
rect 23997 22816 24061 22820
rect 24077 22876 24141 22880
rect 24077 22820 24081 22876
rect 24081 22820 24137 22876
rect 24137 22820 24141 22876
rect 24077 22816 24141 22820
rect 24157 22876 24221 22880
rect 24157 22820 24161 22876
rect 24161 22820 24217 22876
rect 24217 22820 24221 22876
rect 24157 22816 24221 22820
rect 24237 22876 24301 22880
rect 24237 22820 24241 22876
rect 24241 22820 24297 22876
rect 24297 22820 24301 22876
rect 24237 22816 24301 22820
rect 9997 22332 10061 22336
rect 9997 22276 10001 22332
rect 10001 22276 10057 22332
rect 10057 22276 10061 22332
rect 9997 22272 10061 22276
rect 10077 22332 10141 22336
rect 10077 22276 10081 22332
rect 10081 22276 10137 22332
rect 10137 22276 10141 22332
rect 10077 22272 10141 22276
rect 10157 22332 10221 22336
rect 10157 22276 10161 22332
rect 10161 22276 10217 22332
rect 10217 22276 10221 22332
rect 10157 22272 10221 22276
rect 10237 22332 10301 22336
rect 10237 22276 10241 22332
rect 10241 22276 10297 22332
rect 10297 22276 10301 22332
rect 10237 22272 10301 22276
rect 19330 22332 19394 22336
rect 19330 22276 19334 22332
rect 19334 22276 19390 22332
rect 19390 22276 19394 22332
rect 19330 22272 19394 22276
rect 19410 22332 19474 22336
rect 19410 22276 19414 22332
rect 19414 22276 19470 22332
rect 19470 22276 19474 22332
rect 19410 22272 19474 22276
rect 19490 22332 19554 22336
rect 19490 22276 19494 22332
rect 19494 22276 19550 22332
rect 19550 22276 19554 22332
rect 19490 22272 19554 22276
rect 19570 22332 19634 22336
rect 19570 22276 19574 22332
rect 19574 22276 19630 22332
rect 19630 22276 19634 22332
rect 19570 22272 19634 22276
rect 5330 21788 5394 21792
rect 5330 21732 5334 21788
rect 5334 21732 5390 21788
rect 5390 21732 5394 21788
rect 5330 21728 5394 21732
rect 5410 21788 5474 21792
rect 5410 21732 5414 21788
rect 5414 21732 5470 21788
rect 5470 21732 5474 21788
rect 5410 21728 5474 21732
rect 5490 21788 5554 21792
rect 5490 21732 5494 21788
rect 5494 21732 5550 21788
rect 5550 21732 5554 21788
rect 5490 21728 5554 21732
rect 5570 21788 5634 21792
rect 5570 21732 5574 21788
rect 5574 21732 5630 21788
rect 5630 21732 5634 21788
rect 5570 21728 5634 21732
rect 14664 21788 14728 21792
rect 14664 21732 14668 21788
rect 14668 21732 14724 21788
rect 14724 21732 14728 21788
rect 14664 21728 14728 21732
rect 14744 21788 14808 21792
rect 14744 21732 14748 21788
rect 14748 21732 14804 21788
rect 14804 21732 14808 21788
rect 14744 21728 14808 21732
rect 14824 21788 14888 21792
rect 14824 21732 14828 21788
rect 14828 21732 14884 21788
rect 14884 21732 14888 21788
rect 14824 21728 14888 21732
rect 14904 21788 14968 21792
rect 14904 21732 14908 21788
rect 14908 21732 14964 21788
rect 14964 21732 14968 21788
rect 14904 21728 14968 21732
rect 23997 21788 24061 21792
rect 23997 21732 24001 21788
rect 24001 21732 24057 21788
rect 24057 21732 24061 21788
rect 23997 21728 24061 21732
rect 24077 21788 24141 21792
rect 24077 21732 24081 21788
rect 24081 21732 24137 21788
rect 24137 21732 24141 21788
rect 24077 21728 24141 21732
rect 24157 21788 24221 21792
rect 24157 21732 24161 21788
rect 24161 21732 24217 21788
rect 24217 21732 24221 21788
rect 24157 21728 24221 21732
rect 24237 21788 24301 21792
rect 24237 21732 24241 21788
rect 24241 21732 24297 21788
rect 24297 21732 24301 21788
rect 24237 21728 24301 21732
rect 9997 21244 10061 21248
rect 9997 21188 10001 21244
rect 10001 21188 10057 21244
rect 10057 21188 10061 21244
rect 9997 21184 10061 21188
rect 10077 21244 10141 21248
rect 10077 21188 10081 21244
rect 10081 21188 10137 21244
rect 10137 21188 10141 21244
rect 10077 21184 10141 21188
rect 10157 21244 10221 21248
rect 10157 21188 10161 21244
rect 10161 21188 10217 21244
rect 10217 21188 10221 21244
rect 10157 21184 10221 21188
rect 10237 21244 10301 21248
rect 10237 21188 10241 21244
rect 10241 21188 10297 21244
rect 10297 21188 10301 21244
rect 10237 21184 10301 21188
rect 19330 21244 19394 21248
rect 19330 21188 19334 21244
rect 19334 21188 19390 21244
rect 19390 21188 19394 21244
rect 19330 21184 19394 21188
rect 19410 21244 19474 21248
rect 19410 21188 19414 21244
rect 19414 21188 19470 21244
rect 19470 21188 19474 21244
rect 19410 21184 19474 21188
rect 19490 21244 19554 21248
rect 19490 21188 19494 21244
rect 19494 21188 19550 21244
rect 19550 21188 19554 21244
rect 19490 21184 19554 21188
rect 19570 21244 19634 21248
rect 19570 21188 19574 21244
rect 19574 21188 19630 21244
rect 19630 21188 19634 21244
rect 19570 21184 19634 21188
rect 9340 20844 9404 20908
rect 5330 20700 5394 20704
rect 5330 20644 5334 20700
rect 5334 20644 5390 20700
rect 5390 20644 5394 20700
rect 5330 20640 5394 20644
rect 5410 20700 5474 20704
rect 5410 20644 5414 20700
rect 5414 20644 5470 20700
rect 5470 20644 5474 20700
rect 5410 20640 5474 20644
rect 5490 20700 5554 20704
rect 5490 20644 5494 20700
rect 5494 20644 5550 20700
rect 5550 20644 5554 20700
rect 5490 20640 5554 20644
rect 5570 20700 5634 20704
rect 5570 20644 5574 20700
rect 5574 20644 5630 20700
rect 5630 20644 5634 20700
rect 5570 20640 5634 20644
rect 14664 20700 14728 20704
rect 14664 20644 14668 20700
rect 14668 20644 14724 20700
rect 14724 20644 14728 20700
rect 14664 20640 14728 20644
rect 14744 20700 14808 20704
rect 14744 20644 14748 20700
rect 14748 20644 14804 20700
rect 14804 20644 14808 20700
rect 14744 20640 14808 20644
rect 14824 20700 14888 20704
rect 14824 20644 14828 20700
rect 14828 20644 14884 20700
rect 14884 20644 14888 20700
rect 14824 20640 14888 20644
rect 14904 20700 14968 20704
rect 14904 20644 14908 20700
rect 14908 20644 14964 20700
rect 14964 20644 14968 20700
rect 14904 20640 14968 20644
rect 23997 20700 24061 20704
rect 23997 20644 24001 20700
rect 24001 20644 24057 20700
rect 24057 20644 24061 20700
rect 23997 20640 24061 20644
rect 24077 20700 24141 20704
rect 24077 20644 24081 20700
rect 24081 20644 24137 20700
rect 24137 20644 24141 20700
rect 24077 20640 24141 20644
rect 24157 20700 24221 20704
rect 24157 20644 24161 20700
rect 24161 20644 24217 20700
rect 24217 20644 24221 20700
rect 24157 20640 24221 20644
rect 24237 20700 24301 20704
rect 24237 20644 24241 20700
rect 24241 20644 24297 20700
rect 24297 20644 24301 20700
rect 24237 20640 24301 20644
rect 9340 20572 9404 20636
rect 9997 20156 10061 20160
rect 9997 20100 10001 20156
rect 10001 20100 10057 20156
rect 10057 20100 10061 20156
rect 9997 20096 10061 20100
rect 10077 20156 10141 20160
rect 10077 20100 10081 20156
rect 10081 20100 10137 20156
rect 10137 20100 10141 20156
rect 10077 20096 10141 20100
rect 10157 20156 10221 20160
rect 10157 20100 10161 20156
rect 10161 20100 10217 20156
rect 10217 20100 10221 20156
rect 10157 20096 10221 20100
rect 10237 20156 10301 20160
rect 10237 20100 10241 20156
rect 10241 20100 10297 20156
rect 10297 20100 10301 20156
rect 10237 20096 10301 20100
rect 19330 20156 19394 20160
rect 19330 20100 19334 20156
rect 19334 20100 19390 20156
rect 19390 20100 19394 20156
rect 19330 20096 19394 20100
rect 19410 20156 19474 20160
rect 19410 20100 19414 20156
rect 19414 20100 19470 20156
rect 19470 20100 19474 20156
rect 19410 20096 19474 20100
rect 19490 20156 19554 20160
rect 19490 20100 19494 20156
rect 19494 20100 19550 20156
rect 19550 20100 19554 20156
rect 19490 20096 19554 20100
rect 19570 20156 19634 20160
rect 19570 20100 19574 20156
rect 19574 20100 19630 20156
rect 19630 20100 19634 20156
rect 19570 20096 19634 20100
rect 5330 19612 5394 19616
rect 5330 19556 5334 19612
rect 5334 19556 5390 19612
rect 5390 19556 5394 19612
rect 5330 19552 5394 19556
rect 5410 19612 5474 19616
rect 5410 19556 5414 19612
rect 5414 19556 5470 19612
rect 5470 19556 5474 19612
rect 5410 19552 5474 19556
rect 5490 19612 5554 19616
rect 5490 19556 5494 19612
rect 5494 19556 5550 19612
rect 5550 19556 5554 19612
rect 5490 19552 5554 19556
rect 5570 19612 5634 19616
rect 5570 19556 5574 19612
rect 5574 19556 5630 19612
rect 5630 19556 5634 19612
rect 5570 19552 5634 19556
rect 14664 19612 14728 19616
rect 14664 19556 14668 19612
rect 14668 19556 14724 19612
rect 14724 19556 14728 19612
rect 14664 19552 14728 19556
rect 14744 19612 14808 19616
rect 14744 19556 14748 19612
rect 14748 19556 14804 19612
rect 14804 19556 14808 19612
rect 14744 19552 14808 19556
rect 14824 19612 14888 19616
rect 14824 19556 14828 19612
rect 14828 19556 14884 19612
rect 14884 19556 14888 19612
rect 14824 19552 14888 19556
rect 14904 19612 14968 19616
rect 14904 19556 14908 19612
rect 14908 19556 14964 19612
rect 14964 19556 14968 19612
rect 14904 19552 14968 19556
rect 23997 19612 24061 19616
rect 23997 19556 24001 19612
rect 24001 19556 24057 19612
rect 24057 19556 24061 19612
rect 23997 19552 24061 19556
rect 24077 19612 24141 19616
rect 24077 19556 24081 19612
rect 24081 19556 24137 19612
rect 24137 19556 24141 19612
rect 24077 19552 24141 19556
rect 24157 19612 24221 19616
rect 24157 19556 24161 19612
rect 24161 19556 24217 19612
rect 24217 19556 24221 19612
rect 24157 19552 24221 19556
rect 24237 19612 24301 19616
rect 24237 19556 24241 19612
rect 24241 19556 24297 19612
rect 24297 19556 24301 19612
rect 24237 19552 24301 19556
rect 9997 19068 10061 19072
rect 9997 19012 10001 19068
rect 10001 19012 10057 19068
rect 10057 19012 10061 19068
rect 9997 19008 10061 19012
rect 10077 19068 10141 19072
rect 10077 19012 10081 19068
rect 10081 19012 10137 19068
rect 10137 19012 10141 19068
rect 10077 19008 10141 19012
rect 10157 19068 10221 19072
rect 10157 19012 10161 19068
rect 10161 19012 10217 19068
rect 10217 19012 10221 19068
rect 10157 19008 10221 19012
rect 10237 19068 10301 19072
rect 10237 19012 10241 19068
rect 10241 19012 10297 19068
rect 10297 19012 10301 19068
rect 10237 19008 10301 19012
rect 19330 19068 19394 19072
rect 19330 19012 19334 19068
rect 19334 19012 19390 19068
rect 19390 19012 19394 19068
rect 19330 19008 19394 19012
rect 19410 19068 19474 19072
rect 19410 19012 19414 19068
rect 19414 19012 19470 19068
rect 19470 19012 19474 19068
rect 19410 19008 19474 19012
rect 19490 19068 19554 19072
rect 19490 19012 19494 19068
rect 19494 19012 19550 19068
rect 19550 19012 19554 19068
rect 19490 19008 19554 19012
rect 19570 19068 19634 19072
rect 19570 19012 19574 19068
rect 19574 19012 19630 19068
rect 19630 19012 19634 19068
rect 19570 19008 19634 19012
rect 5330 18524 5394 18528
rect 5330 18468 5334 18524
rect 5334 18468 5390 18524
rect 5390 18468 5394 18524
rect 5330 18464 5394 18468
rect 5410 18524 5474 18528
rect 5410 18468 5414 18524
rect 5414 18468 5470 18524
rect 5470 18468 5474 18524
rect 5410 18464 5474 18468
rect 5490 18524 5554 18528
rect 5490 18468 5494 18524
rect 5494 18468 5550 18524
rect 5550 18468 5554 18524
rect 5490 18464 5554 18468
rect 5570 18524 5634 18528
rect 5570 18468 5574 18524
rect 5574 18468 5630 18524
rect 5630 18468 5634 18524
rect 5570 18464 5634 18468
rect 14664 18524 14728 18528
rect 14664 18468 14668 18524
rect 14668 18468 14724 18524
rect 14724 18468 14728 18524
rect 14664 18464 14728 18468
rect 14744 18524 14808 18528
rect 14744 18468 14748 18524
rect 14748 18468 14804 18524
rect 14804 18468 14808 18524
rect 14744 18464 14808 18468
rect 14824 18524 14888 18528
rect 14824 18468 14828 18524
rect 14828 18468 14884 18524
rect 14884 18468 14888 18524
rect 14824 18464 14888 18468
rect 14904 18524 14968 18528
rect 14904 18468 14908 18524
rect 14908 18468 14964 18524
rect 14964 18468 14968 18524
rect 14904 18464 14968 18468
rect 23997 18524 24061 18528
rect 23997 18468 24001 18524
rect 24001 18468 24057 18524
rect 24057 18468 24061 18524
rect 23997 18464 24061 18468
rect 24077 18524 24141 18528
rect 24077 18468 24081 18524
rect 24081 18468 24137 18524
rect 24137 18468 24141 18524
rect 24077 18464 24141 18468
rect 24157 18524 24221 18528
rect 24157 18468 24161 18524
rect 24161 18468 24217 18524
rect 24217 18468 24221 18524
rect 24157 18464 24221 18468
rect 24237 18524 24301 18528
rect 24237 18468 24241 18524
rect 24241 18468 24297 18524
rect 24297 18468 24301 18524
rect 24237 18464 24301 18468
rect 9997 17980 10061 17984
rect 9997 17924 10001 17980
rect 10001 17924 10057 17980
rect 10057 17924 10061 17980
rect 9997 17920 10061 17924
rect 10077 17980 10141 17984
rect 10077 17924 10081 17980
rect 10081 17924 10137 17980
rect 10137 17924 10141 17980
rect 10077 17920 10141 17924
rect 10157 17980 10221 17984
rect 10157 17924 10161 17980
rect 10161 17924 10217 17980
rect 10217 17924 10221 17980
rect 10157 17920 10221 17924
rect 10237 17980 10301 17984
rect 10237 17924 10241 17980
rect 10241 17924 10297 17980
rect 10297 17924 10301 17980
rect 10237 17920 10301 17924
rect 19330 17980 19394 17984
rect 19330 17924 19334 17980
rect 19334 17924 19390 17980
rect 19390 17924 19394 17980
rect 19330 17920 19394 17924
rect 19410 17980 19474 17984
rect 19410 17924 19414 17980
rect 19414 17924 19470 17980
rect 19470 17924 19474 17980
rect 19410 17920 19474 17924
rect 19490 17980 19554 17984
rect 19490 17924 19494 17980
rect 19494 17924 19550 17980
rect 19550 17924 19554 17980
rect 19490 17920 19554 17924
rect 19570 17980 19634 17984
rect 19570 17924 19574 17980
rect 19574 17924 19630 17980
rect 19630 17924 19634 17980
rect 19570 17920 19634 17924
rect 5330 17436 5394 17440
rect 5330 17380 5334 17436
rect 5334 17380 5390 17436
rect 5390 17380 5394 17436
rect 5330 17376 5394 17380
rect 5410 17436 5474 17440
rect 5410 17380 5414 17436
rect 5414 17380 5470 17436
rect 5470 17380 5474 17436
rect 5410 17376 5474 17380
rect 5490 17436 5554 17440
rect 5490 17380 5494 17436
rect 5494 17380 5550 17436
rect 5550 17380 5554 17436
rect 5490 17376 5554 17380
rect 5570 17436 5634 17440
rect 5570 17380 5574 17436
rect 5574 17380 5630 17436
rect 5630 17380 5634 17436
rect 5570 17376 5634 17380
rect 14664 17436 14728 17440
rect 14664 17380 14668 17436
rect 14668 17380 14724 17436
rect 14724 17380 14728 17436
rect 14664 17376 14728 17380
rect 14744 17436 14808 17440
rect 14744 17380 14748 17436
rect 14748 17380 14804 17436
rect 14804 17380 14808 17436
rect 14744 17376 14808 17380
rect 14824 17436 14888 17440
rect 14824 17380 14828 17436
rect 14828 17380 14884 17436
rect 14884 17380 14888 17436
rect 14824 17376 14888 17380
rect 14904 17436 14968 17440
rect 14904 17380 14908 17436
rect 14908 17380 14964 17436
rect 14964 17380 14968 17436
rect 14904 17376 14968 17380
rect 23997 17436 24061 17440
rect 23997 17380 24001 17436
rect 24001 17380 24057 17436
rect 24057 17380 24061 17436
rect 23997 17376 24061 17380
rect 24077 17436 24141 17440
rect 24077 17380 24081 17436
rect 24081 17380 24137 17436
rect 24137 17380 24141 17436
rect 24077 17376 24141 17380
rect 24157 17436 24221 17440
rect 24157 17380 24161 17436
rect 24161 17380 24217 17436
rect 24217 17380 24221 17436
rect 24157 17376 24221 17380
rect 24237 17436 24301 17440
rect 24237 17380 24241 17436
rect 24241 17380 24297 17436
rect 24297 17380 24301 17436
rect 24237 17376 24301 17380
rect 9997 16892 10061 16896
rect 9997 16836 10001 16892
rect 10001 16836 10057 16892
rect 10057 16836 10061 16892
rect 9997 16832 10061 16836
rect 10077 16892 10141 16896
rect 10077 16836 10081 16892
rect 10081 16836 10137 16892
rect 10137 16836 10141 16892
rect 10077 16832 10141 16836
rect 10157 16892 10221 16896
rect 10157 16836 10161 16892
rect 10161 16836 10217 16892
rect 10217 16836 10221 16892
rect 10157 16832 10221 16836
rect 10237 16892 10301 16896
rect 10237 16836 10241 16892
rect 10241 16836 10297 16892
rect 10297 16836 10301 16892
rect 10237 16832 10301 16836
rect 19330 16892 19394 16896
rect 19330 16836 19334 16892
rect 19334 16836 19390 16892
rect 19390 16836 19394 16892
rect 19330 16832 19394 16836
rect 19410 16892 19474 16896
rect 19410 16836 19414 16892
rect 19414 16836 19470 16892
rect 19470 16836 19474 16892
rect 19410 16832 19474 16836
rect 19490 16892 19554 16896
rect 19490 16836 19494 16892
rect 19494 16836 19550 16892
rect 19550 16836 19554 16892
rect 19490 16832 19554 16836
rect 19570 16892 19634 16896
rect 19570 16836 19574 16892
rect 19574 16836 19630 16892
rect 19630 16836 19634 16892
rect 19570 16832 19634 16836
rect 5330 16348 5394 16352
rect 5330 16292 5334 16348
rect 5334 16292 5390 16348
rect 5390 16292 5394 16348
rect 5330 16288 5394 16292
rect 5410 16348 5474 16352
rect 5410 16292 5414 16348
rect 5414 16292 5470 16348
rect 5470 16292 5474 16348
rect 5410 16288 5474 16292
rect 5490 16348 5554 16352
rect 5490 16292 5494 16348
rect 5494 16292 5550 16348
rect 5550 16292 5554 16348
rect 5490 16288 5554 16292
rect 5570 16348 5634 16352
rect 5570 16292 5574 16348
rect 5574 16292 5630 16348
rect 5630 16292 5634 16348
rect 5570 16288 5634 16292
rect 14664 16348 14728 16352
rect 14664 16292 14668 16348
rect 14668 16292 14724 16348
rect 14724 16292 14728 16348
rect 14664 16288 14728 16292
rect 14744 16348 14808 16352
rect 14744 16292 14748 16348
rect 14748 16292 14804 16348
rect 14804 16292 14808 16348
rect 14744 16288 14808 16292
rect 14824 16348 14888 16352
rect 14824 16292 14828 16348
rect 14828 16292 14884 16348
rect 14884 16292 14888 16348
rect 14824 16288 14888 16292
rect 14904 16348 14968 16352
rect 14904 16292 14908 16348
rect 14908 16292 14964 16348
rect 14964 16292 14968 16348
rect 14904 16288 14968 16292
rect 23997 16348 24061 16352
rect 23997 16292 24001 16348
rect 24001 16292 24057 16348
rect 24057 16292 24061 16348
rect 23997 16288 24061 16292
rect 24077 16348 24141 16352
rect 24077 16292 24081 16348
rect 24081 16292 24137 16348
rect 24137 16292 24141 16348
rect 24077 16288 24141 16292
rect 24157 16348 24221 16352
rect 24157 16292 24161 16348
rect 24161 16292 24217 16348
rect 24217 16292 24221 16348
rect 24157 16288 24221 16292
rect 24237 16348 24301 16352
rect 24237 16292 24241 16348
rect 24241 16292 24297 16348
rect 24297 16292 24301 16348
rect 24237 16288 24301 16292
rect 9997 15804 10061 15808
rect 9997 15748 10001 15804
rect 10001 15748 10057 15804
rect 10057 15748 10061 15804
rect 9997 15744 10061 15748
rect 10077 15804 10141 15808
rect 10077 15748 10081 15804
rect 10081 15748 10137 15804
rect 10137 15748 10141 15804
rect 10077 15744 10141 15748
rect 10157 15804 10221 15808
rect 10157 15748 10161 15804
rect 10161 15748 10217 15804
rect 10217 15748 10221 15804
rect 10157 15744 10221 15748
rect 10237 15804 10301 15808
rect 10237 15748 10241 15804
rect 10241 15748 10297 15804
rect 10297 15748 10301 15804
rect 10237 15744 10301 15748
rect 19330 15804 19394 15808
rect 19330 15748 19334 15804
rect 19334 15748 19390 15804
rect 19390 15748 19394 15804
rect 19330 15744 19394 15748
rect 19410 15804 19474 15808
rect 19410 15748 19414 15804
rect 19414 15748 19470 15804
rect 19470 15748 19474 15804
rect 19410 15744 19474 15748
rect 19490 15804 19554 15808
rect 19490 15748 19494 15804
rect 19494 15748 19550 15804
rect 19550 15748 19554 15804
rect 19490 15744 19554 15748
rect 19570 15804 19634 15808
rect 19570 15748 19574 15804
rect 19574 15748 19630 15804
rect 19630 15748 19634 15804
rect 19570 15744 19634 15748
rect 5330 15260 5394 15264
rect 5330 15204 5334 15260
rect 5334 15204 5390 15260
rect 5390 15204 5394 15260
rect 5330 15200 5394 15204
rect 5410 15260 5474 15264
rect 5410 15204 5414 15260
rect 5414 15204 5470 15260
rect 5470 15204 5474 15260
rect 5410 15200 5474 15204
rect 5490 15260 5554 15264
rect 5490 15204 5494 15260
rect 5494 15204 5550 15260
rect 5550 15204 5554 15260
rect 5490 15200 5554 15204
rect 5570 15260 5634 15264
rect 5570 15204 5574 15260
rect 5574 15204 5630 15260
rect 5630 15204 5634 15260
rect 5570 15200 5634 15204
rect 14664 15260 14728 15264
rect 14664 15204 14668 15260
rect 14668 15204 14724 15260
rect 14724 15204 14728 15260
rect 14664 15200 14728 15204
rect 14744 15260 14808 15264
rect 14744 15204 14748 15260
rect 14748 15204 14804 15260
rect 14804 15204 14808 15260
rect 14744 15200 14808 15204
rect 14824 15260 14888 15264
rect 14824 15204 14828 15260
rect 14828 15204 14884 15260
rect 14884 15204 14888 15260
rect 14824 15200 14888 15204
rect 14904 15260 14968 15264
rect 14904 15204 14908 15260
rect 14908 15204 14964 15260
rect 14964 15204 14968 15260
rect 14904 15200 14968 15204
rect 23997 15260 24061 15264
rect 23997 15204 24001 15260
rect 24001 15204 24057 15260
rect 24057 15204 24061 15260
rect 23997 15200 24061 15204
rect 24077 15260 24141 15264
rect 24077 15204 24081 15260
rect 24081 15204 24137 15260
rect 24137 15204 24141 15260
rect 24077 15200 24141 15204
rect 24157 15260 24221 15264
rect 24157 15204 24161 15260
rect 24161 15204 24217 15260
rect 24217 15204 24221 15260
rect 24157 15200 24221 15204
rect 24237 15260 24301 15264
rect 24237 15204 24241 15260
rect 24241 15204 24297 15260
rect 24297 15204 24301 15260
rect 24237 15200 24301 15204
rect 9997 14716 10061 14720
rect 9997 14660 10001 14716
rect 10001 14660 10057 14716
rect 10057 14660 10061 14716
rect 9997 14656 10061 14660
rect 10077 14716 10141 14720
rect 10077 14660 10081 14716
rect 10081 14660 10137 14716
rect 10137 14660 10141 14716
rect 10077 14656 10141 14660
rect 10157 14716 10221 14720
rect 10157 14660 10161 14716
rect 10161 14660 10217 14716
rect 10217 14660 10221 14716
rect 10157 14656 10221 14660
rect 10237 14716 10301 14720
rect 10237 14660 10241 14716
rect 10241 14660 10297 14716
rect 10297 14660 10301 14716
rect 10237 14656 10301 14660
rect 19330 14716 19394 14720
rect 19330 14660 19334 14716
rect 19334 14660 19390 14716
rect 19390 14660 19394 14716
rect 19330 14656 19394 14660
rect 19410 14716 19474 14720
rect 19410 14660 19414 14716
rect 19414 14660 19470 14716
rect 19470 14660 19474 14716
rect 19410 14656 19474 14660
rect 19490 14716 19554 14720
rect 19490 14660 19494 14716
rect 19494 14660 19550 14716
rect 19550 14660 19554 14716
rect 19490 14656 19554 14660
rect 19570 14716 19634 14720
rect 19570 14660 19574 14716
rect 19574 14660 19630 14716
rect 19630 14660 19634 14716
rect 19570 14656 19634 14660
rect 5330 14172 5394 14176
rect 5330 14116 5334 14172
rect 5334 14116 5390 14172
rect 5390 14116 5394 14172
rect 5330 14112 5394 14116
rect 5410 14172 5474 14176
rect 5410 14116 5414 14172
rect 5414 14116 5470 14172
rect 5470 14116 5474 14172
rect 5410 14112 5474 14116
rect 5490 14172 5554 14176
rect 5490 14116 5494 14172
rect 5494 14116 5550 14172
rect 5550 14116 5554 14172
rect 5490 14112 5554 14116
rect 5570 14172 5634 14176
rect 5570 14116 5574 14172
rect 5574 14116 5630 14172
rect 5630 14116 5634 14172
rect 5570 14112 5634 14116
rect 14664 14172 14728 14176
rect 14664 14116 14668 14172
rect 14668 14116 14724 14172
rect 14724 14116 14728 14172
rect 14664 14112 14728 14116
rect 14744 14172 14808 14176
rect 14744 14116 14748 14172
rect 14748 14116 14804 14172
rect 14804 14116 14808 14172
rect 14744 14112 14808 14116
rect 14824 14172 14888 14176
rect 14824 14116 14828 14172
rect 14828 14116 14884 14172
rect 14884 14116 14888 14172
rect 14824 14112 14888 14116
rect 14904 14172 14968 14176
rect 14904 14116 14908 14172
rect 14908 14116 14964 14172
rect 14964 14116 14968 14172
rect 14904 14112 14968 14116
rect 23997 14172 24061 14176
rect 23997 14116 24001 14172
rect 24001 14116 24057 14172
rect 24057 14116 24061 14172
rect 23997 14112 24061 14116
rect 24077 14172 24141 14176
rect 24077 14116 24081 14172
rect 24081 14116 24137 14172
rect 24137 14116 24141 14172
rect 24077 14112 24141 14116
rect 24157 14172 24221 14176
rect 24157 14116 24161 14172
rect 24161 14116 24217 14172
rect 24217 14116 24221 14172
rect 24157 14112 24221 14116
rect 24237 14172 24301 14176
rect 24237 14116 24241 14172
rect 24241 14116 24297 14172
rect 24297 14116 24301 14172
rect 24237 14112 24301 14116
rect 9997 13628 10061 13632
rect 9997 13572 10001 13628
rect 10001 13572 10057 13628
rect 10057 13572 10061 13628
rect 9997 13568 10061 13572
rect 10077 13628 10141 13632
rect 10077 13572 10081 13628
rect 10081 13572 10137 13628
rect 10137 13572 10141 13628
rect 10077 13568 10141 13572
rect 10157 13628 10221 13632
rect 10157 13572 10161 13628
rect 10161 13572 10217 13628
rect 10217 13572 10221 13628
rect 10157 13568 10221 13572
rect 10237 13628 10301 13632
rect 10237 13572 10241 13628
rect 10241 13572 10297 13628
rect 10297 13572 10301 13628
rect 10237 13568 10301 13572
rect 19330 13628 19394 13632
rect 19330 13572 19334 13628
rect 19334 13572 19390 13628
rect 19390 13572 19394 13628
rect 19330 13568 19394 13572
rect 19410 13628 19474 13632
rect 19410 13572 19414 13628
rect 19414 13572 19470 13628
rect 19470 13572 19474 13628
rect 19410 13568 19474 13572
rect 19490 13628 19554 13632
rect 19490 13572 19494 13628
rect 19494 13572 19550 13628
rect 19550 13572 19554 13628
rect 19490 13568 19554 13572
rect 19570 13628 19634 13632
rect 19570 13572 19574 13628
rect 19574 13572 19630 13628
rect 19630 13572 19634 13628
rect 19570 13568 19634 13572
rect 5330 13084 5394 13088
rect 5330 13028 5334 13084
rect 5334 13028 5390 13084
rect 5390 13028 5394 13084
rect 5330 13024 5394 13028
rect 5410 13084 5474 13088
rect 5410 13028 5414 13084
rect 5414 13028 5470 13084
rect 5470 13028 5474 13084
rect 5410 13024 5474 13028
rect 5490 13084 5554 13088
rect 5490 13028 5494 13084
rect 5494 13028 5550 13084
rect 5550 13028 5554 13084
rect 5490 13024 5554 13028
rect 5570 13084 5634 13088
rect 5570 13028 5574 13084
rect 5574 13028 5630 13084
rect 5630 13028 5634 13084
rect 5570 13024 5634 13028
rect 14664 13084 14728 13088
rect 14664 13028 14668 13084
rect 14668 13028 14724 13084
rect 14724 13028 14728 13084
rect 14664 13024 14728 13028
rect 14744 13084 14808 13088
rect 14744 13028 14748 13084
rect 14748 13028 14804 13084
rect 14804 13028 14808 13084
rect 14744 13024 14808 13028
rect 14824 13084 14888 13088
rect 14824 13028 14828 13084
rect 14828 13028 14884 13084
rect 14884 13028 14888 13084
rect 14824 13024 14888 13028
rect 14904 13084 14968 13088
rect 14904 13028 14908 13084
rect 14908 13028 14964 13084
rect 14964 13028 14968 13084
rect 14904 13024 14968 13028
rect 23997 13084 24061 13088
rect 23997 13028 24001 13084
rect 24001 13028 24057 13084
rect 24057 13028 24061 13084
rect 23997 13024 24061 13028
rect 24077 13084 24141 13088
rect 24077 13028 24081 13084
rect 24081 13028 24137 13084
rect 24137 13028 24141 13084
rect 24077 13024 24141 13028
rect 24157 13084 24221 13088
rect 24157 13028 24161 13084
rect 24161 13028 24217 13084
rect 24217 13028 24221 13084
rect 24157 13024 24221 13028
rect 24237 13084 24301 13088
rect 24237 13028 24241 13084
rect 24241 13028 24297 13084
rect 24297 13028 24301 13084
rect 24237 13024 24301 13028
rect 9997 12540 10061 12544
rect 9997 12484 10001 12540
rect 10001 12484 10057 12540
rect 10057 12484 10061 12540
rect 9997 12480 10061 12484
rect 10077 12540 10141 12544
rect 10077 12484 10081 12540
rect 10081 12484 10137 12540
rect 10137 12484 10141 12540
rect 10077 12480 10141 12484
rect 10157 12540 10221 12544
rect 10157 12484 10161 12540
rect 10161 12484 10217 12540
rect 10217 12484 10221 12540
rect 10157 12480 10221 12484
rect 10237 12540 10301 12544
rect 10237 12484 10241 12540
rect 10241 12484 10297 12540
rect 10297 12484 10301 12540
rect 10237 12480 10301 12484
rect 19330 12540 19394 12544
rect 19330 12484 19334 12540
rect 19334 12484 19390 12540
rect 19390 12484 19394 12540
rect 19330 12480 19394 12484
rect 19410 12540 19474 12544
rect 19410 12484 19414 12540
rect 19414 12484 19470 12540
rect 19470 12484 19474 12540
rect 19410 12480 19474 12484
rect 19490 12540 19554 12544
rect 19490 12484 19494 12540
rect 19494 12484 19550 12540
rect 19550 12484 19554 12540
rect 19490 12480 19554 12484
rect 19570 12540 19634 12544
rect 19570 12484 19574 12540
rect 19574 12484 19630 12540
rect 19630 12484 19634 12540
rect 19570 12480 19634 12484
rect 5330 11996 5394 12000
rect 5330 11940 5334 11996
rect 5334 11940 5390 11996
rect 5390 11940 5394 11996
rect 5330 11936 5394 11940
rect 5410 11996 5474 12000
rect 5410 11940 5414 11996
rect 5414 11940 5470 11996
rect 5470 11940 5474 11996
rect 5410 11936 5474 11940
rect 5490 11996 5554 12000
rect 5490 11940 5494 11996
rect 5494 11940 5550 11996
rect 5550 11940 5554 11996
rect 5490 11936 5554 11940
rect 5570 11996 5634 12000
rect 5570 11940 5574 11996
rect 5574 11940 5630 11996
rect 5630 11940 5634 11996
rect 5570 11936 5634 11940
rect 14664 11996 14728 12000
rect 14664 11940 14668 11996
rect 14668 11940 14724 11996
rect 14724 11940 14728 11996
rect 14664 11936 14728 11940
rect 14744 11996 14808 12000
rect 14744 11940 14748 11996
rect 14748 11940 14804 11996
rect 14804 11940 14808 11996
rect 14744 11936 14808 11940
rect 14824 11996 14888 12000
rect 14824 11940 14828 11996
rect 14828 11940 14884 11996
rect 14884 11940 14888 11996
rect 14824 11936 14888 11940
rect 14904 11996 14968 12000
rect 14904 11940 14908 11996
rect 14908 11940 14964 11996
rect 14964 11940 14968 11996
rect 14904 11936 14968 11940
rect 23997 11996 24061 12000
rect 23997 11940 24001 11996
rect 24001 11940 24057 11996
rect 24057 11940 24061 11996
rect 23997 11936 24061 11940
rect 24077 11996 24141 12000
rect 24077 11940 24081 11996
rect 24081 11940 24137 11996
rect 24137 11940 24141 11996
rect 24077 11936 24141 11940
rect 24157 11996 24221 12000
rect 24157 11940 24161 11996
rect 24161 11940 24217 11996
rect 24217 11940 24221 11996
rect 24157 11936 24221 11940
rect 24237 11996 24301 12000
rect 24237 11940 24241 11996
rect 24241 11940 24297 11996
rect 24297 11940 24301 11996
rect 24237 11936 24301 11940
rect 9997 11452 10061 11456
rect 9997 11396 10001 11452
rect 10001 11396 10057 11452
rect 10057 11396 10061 11452
rect 9997 11392 10061 11396
rect 10077 11452 10141 11456
rect 10077 11396 10081 11452
rect 10081 11396 10137 11452
rect 10137 11396 10141 11452
rect 10077 11392 10141 11396
rect 10157 11452 10221 11456
rect 10157 11396 10161 11452
rect 10161 11396 10217 11452
rect 10217 11396 10221 11452
rect 10157 11392 10221 11396
rect 10237 11452 10301 11456
rect 10237 11396 10241 11452
rect 10241 11396 10297 11452
rect 10297 11396 10301 11452
rect 10237 11392 10301 11396
rect 19330 11452 19394 11456
rect 19330 11396 19334 11452
rect 19334 11396 19390 11452
rect 19390 11396 19394 11452
rect 19330 11392 19394 11396
rect 19410 11452 19474 11456
rect 19410 11396 19414 11452
rect 19414 11396 19470 11452
rect 19470 11396 19474 11452
rect 19410 11392 19474 11396
rect 19490 11452 19554 11456
rect 19490 11396 19494 11452
rect 19494 11396 19550 11452
rect 19550 11396 19554 11452
rect 19490 11392 19554 11396
rect 19570 11452 19634 11456
rect 19570 11396 19574 11452
rect 19574 11396 19630 11452
rect 19630 11396 19634 11452
rect 19570 11392 19634 11396
rect 5330 10908 5394 10912
rect 5330 10852 5334 10908
rect 5334 10852 5390 10908
rect 5390 10852 5394 10908
rect 5330 10848 5394 10852
rect 5410 10908 5474 10912
rect 5410 10852 5414 10908
rect 5414 10852 5470 10908
rect 5470 10852 5474 10908
rect 5410 10848 5474 10852
rect 5490 10908 5554 10912
rect 5490 10852 5494 10908
rect 5494 10852 5550 10908
rect 5550 10852 5554 10908
rect 5490 10848 5554 10852
rect 5570 10908 5634 10912
rect 5570 10852 5574 10908
rect 5574 10852 5630 10908
rect 5630 10852 5634 10908
rect 5570 10848 5634 10852
rect 14664 10908 14728 10912
rect 14664 10852 14668 10908
rect 14668 10852 14724 10908
rect 14724 10852 14728 10908
rect 14664 10848 14728 10852
rect 14744 10908 14808 10912
rect 14744 10852 14748 10908
rect 14748 10852 14804 10908
rect 14804 10852 14808 10908
rect 14744 10848 14808 10852
rect 14824 10908 14888 10912
rect 14824 10852 14828 10908
rect 14828 10852 14884 10908
rect 14884 10852 14888 10908
rect 14824 10848 14888 10852
rect 14904 10908 14968 10912
rect 14904 10852 14908 10908
rect 14908 10852 14964 10908
rect 14964 10852 14968 10908
rect 14904 10848 14968 10852
rect 23997 10908 24061 10912
rect 23997 10852 24001 10908
rect 24001 10852 24057 10908
rect 24057 10852 24061 10908
rect 23997 10848 24061 10852
rect 24077 10908 24141 10912
rect 24077 10852 24081 10908
rect 24081 10852 24137 10908
rect 24137 10852 24141 10908
rect 24077 10848 24141 10852
rect 24157 10908 24221 10912
rect 24157 10852 24161 10908
rect 24161 10852 24217 10908
rect 24217 10852 24221 10908
rect 24157 10848 24221 10852
rect 24237 10908 24301 10912
rect 24237 10852 24241 10908
rect 24241 10852 24297 10908
rect 24297 10852 24301 10908
rect 24237 10848 24301 10852
rect 9997 10364 10061 10368
rect 9997 10308 10001 10364
rect 10001 10308 10057 10364
rect 10057 10308 10061 10364
rect 9997 10304 10061 10308
rect 10077 10364 10141 10368
rect 10077 10308 10081 10364
rect 10081 10308 10137 10364
rect 10137 10308 10141 10364
rect 10077 10304 10141 10308
rect 10157 10364 10221 10368
rect 10157 10308 10161 10364
rect 10161 10308 10217 10364
rect 10217 10308 10221 10364
rect 10157 10304 10221 10308
rect 10237 10364 10301 10368
rect 10237 10308 10241 10364
rect 10241 10308 10297 10364
rect 10297 10308 10301 10364
rect 10237 10304 10301 10308
rect 19330 10364 19394 10368
rect 19330 10308 19334 10364
rect 19334 10308 19390 10364
rect 19390 10308 19394 10364
rect 19330 10304 19394 10308
rect 19410 10364 19474 10368
rect 19410 10308 19414 10364
rect 19414 10308 19470 10364
rect 19470 10308 19474 10364
rect 19410 10304 19474 10308
rect 19490 10364 19554 10368
rect 19490 10308 19494 10364
rect 19494 10308 19550 10364
rect 19550 10308 19554 10364
rect 19490 10304 19554 10308
rect 19570 10364 19634 10368
rect 19570 10308 19574 10364
rect 19574 10308 19630 10364
rect 19630 10308 19634 10364
rect 19570 10304 19634 10308
rect 5330 9820 5394 9824
rect 5330 9764 5334 9820
rect 5334 9764 5390 9820
rect 5390 9764 5394 9820
rect 5330 9760 5394 9764
rect 5410 9820 5474 9824
rect 5410 9764 5414 9820
rect 5414 9764 5470 9820
rect 5470 9764 5474 9820
rect 5410 9760 5474 9764
rect 5490 9820 5554 9824
rect 5490 9764 5494 9820
rect 5494 9764 5550 9820
rect 5550 9764 5554 9820
rect 5490 9760 5554 9764
rect 5570 9820 5634 9824
rect 5570 9764 5574 9820
rect 5574 9764 5630 9820
rect 5630 9764 5634 9820
rect 5570 9760 5634 9764
rect 14664 9820 14728 9824
rect 14664 9764 14668 9820
rect 14668 9764 14724 9820
rect 14724 9764 14728 9820
rect 14664 9760 14728 9764
rect 14744 9820 14808 9824
rect 14744 9764 14748 9820
rect 14748 9764 14804 9820
rect 14804 9764 14808 9820
rect 14744 9760 14808 9764
rect 14824 9820 14888 9824
rect 14824 9764 14828 9820
rect 14828 9764 14884 9820
rect 14884 9764 14888 9820
rect 14824 9760 14888 9764
rect 14904 9820 14968 9824
rect 14904 9764 14908 9820
rect 14908 9764 14964 9820
rect 14964 9764 14968 9820
rect 14904 9760 14968 9764
rect 23997 9820 24061 9824
rect 23997 9764 24001 9820
rect 24001 9764 24057 9820
rect 24057 9764 24061 9820
rect 23997 9760 24061 9764
rect 24077 9820 24141 9824
rect 24077 9764 24081 9820
rect 24081 9764 24137 9820
rect 24137 9764 24141 9820
rect 24077 9760 24141 9764
rect 24157 9820 24221 9824
rect 24157 9764 24161 9820
rect 24161 9764 24217 9820
rect 24217 9764 24221 9820
rect 24157 9760 24221 9764
rect 24237 9820 24301 9824
rect 24237 9764 24241 9820
rect 24241 9764 24297 9820
rect 24297 9764 24301 9820
rect 24237 9760 24301 9764
rect 9997 9276 10061 9280
rect 9997 9220 10001 9276
rect 10001 9220 10057 9276
rect 10057 9220 10061 9276
rect 9997 9216 10061 9220
rect 10077 9276 10141 9280
rect 10077 9220 10081 9276
rect 10081 9220 10137 9276
rect 10137 9220 10141 9276
rect 10077 9216 10141 9220
rect 10157 9276 10221 9280
rect 10157 9220 10161 9276
rect 10161 9220 10217 9276
rect 10217 9220 10221 9276
rect 10157 9216 10221 9220
rect 10237 9276 10301 9280
rect 10237 9220 10241 9276
rect 10241 9220 10297 9276
rect 10297 9220 10301 9276
rect 10237 9216 10301 9220
rect 19330 9276 19394 9280
rect 19330 9220 19334 9276
rect 19334 9220 19390 9276
rect 19390 9220 19394 9276
rect 19330 9216 19394 9220
rect 19410 9276 19474 9280
rect 19410 9220 19414 9276
rect 19414 9220 19470 9276
rect 19470 9220 19474 9276
rect 19410 9216 19474 9220
rect 19490 9276 19554 9280
rect 19490 9220 19494 9276
rect 19494 9220 19550 9276
rect 19550 9220 19554 9276
rect 19490 9216 19554 9220
rect 19570 9276 19634 9280
rect 19570 9220 19574 9276
rect 19574 9220 19630 9276
rect 19630 9220 19634 9276
rect 19570 9216 19634 9220
rect 5330 8732 5394 8736
rect 5330 8676 5334 8732
rect 5334 8676 5390 8732
rect 5390 8676 5394 8732
rect 5330 8672 5394 8676
rect 5410 8732 5474 8736
rect 5410 8676 5414 8732
rect 5414 8676 5470 8732
rect 5470 8676 5474 8732
rect 5410 8672 5474 8676
rect 5490 8732 5554 8736
rect 5490 8676 5494 8732
rect 5494 8676 5550 8732
rect 5550 8676 5554 8732
rect 5490 8672 5554 8676
rect 5570 8732 5634 8736
rect 5570 8676 5574 8732
rect 5574 8676 5630 8732
rect 5630 8676 5634 8732
rect 5570 8672 5634 8676
rect 14664 8732 14728 8736
rect 14664 8676 14668 8732
rect 14668 8676 14724 8732
rect 14724 8676 14728 8732
rect 14664 8672 14728 8676
rect 14744 8732 14808 8736
rect 14744 8676 14748 8732
rect 14748 8676 14804 8732
rect 14804 8676 14808 8732
rect 14744 8672 14808 8676
rect 14824 8732 14888 8736
rect 14824 8676 14828 8732
rect 14828 8676 14884 8732
rect 14884 8676 14888 8732
rect 14824 8672 14888 8676
rect 14904 8732 14968 8736
rect 14904 8676 14908 8732
rect 14908 8676 14964 8732
rect 14964 8676 14968 8732
rect 14904 8672 14968 8676
rect 23997 8732 24061 8736
rect 23997 8676 24001 8732
rect 24001 8676 24057 8732
rect 24057 8676 24061 8732
rect 23997 8672 24061 8676
rect 24077 8732 24141 8736
rect 24077 8676 24081 8732
rect 24081 8676 24137 8732
rect 24137 8676 24141 8732
rect 24077 8672 24141 8676
rect 24157 8732 24221 8736
rect 24157 8676 24161 8732
rect 24161 8676 24217 8732
rect 24217 8676 24221 8732
rect 24157 8672 24221 8676
rect 24237 8732 24301 8736
rect 24237 8676 24241 8732
rect 24241 8676 24297 8732
rect 24297 8676 24301 8732
rect 24237 8672 24301 8676
rect 9997 8188 10061 8192
rect 9997 8132 10001 8188
rect 10001 8132 10057 8188
rect 10057 8132 10061 8188
rect 9997 8128 10061 8132
rect 10077 8188 10141 8192
rect 10077 8132 10081 8188
rect 10081 8132 10137 8188
rect 10137 8132 10141 8188
rect 10077 8128 10141 8132
rect 10157 8188 10221 8192
rect 10157 8132 10161 8188
rect 10161 8132 10217 8188
rect 10217 8132 10221 8188
rect 10157 8128 10221 8132
rect 10237 8188 10301 8192
rect 10237 8132 10241 8188
rect 10241 8132 10297 8188
rect 10297 8132 10301 8188
rect 10237 8128 10301 8132
rect 19330 8188 19394 8192
rect 19330 8132 19334 8188
rect 19334 8132 19390 8188
rect 19390 8132 19394 8188
rect 19330 8128 19394 8132
rect 19410 8188 19474 8192
rect 19410 8132 19414 8188
rect 19414 8132 19470 8188
rect 19470 8132 19474 8188
rect 19410 8128 19474 8132
rect 19490 8188 19554 8192
rect 19490 8132 19494 8188
rect 19494 8132 19550 8188
rect 19550 8132 19554 8188
rect 19490 8128 19554 8132
rect 19570 8188 19634 8192
rect 19570 8132 19574 8188
rect 19574 8132 19630 8188
rect 19630 8132 19634 8188
rect 19570 8128 19634 8132
rect 5330 7644 5394 7648
rect 5330 7588 5334 7644
rect 5334 7588 5390 7644
rect 5390 7588 5394 7644
rect 5330 7584 5394 7588
rect 5410 7644 5474 7648
rect 5410 7588 5414 7644
rect 5414 7588 5470 7644
rect 5470 7588 5474 7644
rect 5410 7584 5474 7588
rect 5490 7644 5554 7648
rect 5490 7588 5494 7644
rect 5494 7588 5550 7644
rect 5550 7588 5554 7644
rect 5490 7584 5554 7588
rect 5570 7644 5634 7648
rect 5570 7588 5574 7644
rect 5574 7588 5630 7644
rect 5630 7588 5634 7644
rect 5570 7584 5634 7588
rect 14664 7644 14728 7648
rect 14664 7588 14668 7644
rect 14668 7588 14724 7644
rect 14724 7588 14728 7644
rect 14664 7584 14728 7588
rect 14744 7644 14808 7648
rect 14744 7588 14748 7644
rect 14748 7588 14804 7644
rect 14804 7588 14808 7644
rect 14744 7584 14808 7588
rect 14824 7644 14888 7648
rect 14824 7588 14828 7644
rect 14828 7588 14884 7644
rect 14884 7588 14888 7644
rect 14824 7584 14888 7588
rect 14904 7644 14968 7648
rect 14904 7588 14908 7644
rect 14908 7588 14964 7644
rect 14964 7588 14968 7644
rect 14904 7584 14968 7588
rect 23997 7644 24061 7648
rect 23997 7588 24001 7644
rect 24001 7588 24057 7644
rect 24057 7588 24061 7644
rect 23997 7584 24061 7588
rect 24077 7644 24141 7648
rect 24077 7588 24081 7644
rect 24081 7588 24137 7644
rect 24137 7588 24141 7644
rect 24077 7584 24141 7588
rect 24157 7644 24221 7648
rect 24157 7588 24161 7644
rect 24161 7588 24217 7644
rect 24217 7588 24221 7644
rect 24157 7584 24221 7588
rect 24237 7644 24301 7648
rect 24237 7588 24241 7644
rect 24241 7588 24297 7644
rect 24297 7588 24301 7644
rect 24237 7584 24301 7588
rect 9997 7100 10061 7104
rect 9997 7044 10001 7100
rect 10001 7044 10057 7100
rect 10057 7044 10061 7100
rect 9997 7040 10061 7044
rect 10077 7100 10141 7104
rect 10077 7044 10081 7100
rect 10081 7044 10137 7100
rect 10137 7044 10141 7100
rect 10077 7040 10141 7044
rect 10157 7100 10221 7104
rect 10157 7044 10161 7100
rect 10161 7044 10217 7100
rect 10217 7044 10221 7100
rect 10157 7040 10221 7044
rect 10237 7100 10301 7104
rect 10237 7044 10241 7100
rect 10241 7044 10297 7100
rect 10297 7044 10301 7100
rect 10237 7040 10301 7044
rect 19330 7100 19394 7104
rect 19330 7044 19334 7100
rect 19334 7044 19390 7100
rect 19390 7044 19394 7100
rect 19330 7040 19394 7044
rect 19410 7100 19474 7104
rect 19410 7044 19414 7100
rect 19414 7044 19470 7100
rect 19470 7044 19474 7100
rect 19410 7040 19474 7044
rect 19490 7100 19554 7104
rect 19490 7044 19494 7100
rect 19494 7044 19550 7100
rect 19550 7044 19554 7100
rect 19490 7040 19554 7044
rect 19570 7100 19634 7104
rect 19570 7044 19574 7100
rect 19574 7044 19630 7100
rect 19630 7044 19634 7100
rect 19570 7040 19634 7044
rect 5330 6556 5394 6560
rect 5330 6500 5334 6556
rect 5334 6500 5390 6556
rect 5390 6500 5394 6556
rect 5330 6496 5394 6500
rect 5410 6556 5474 6560
rect 5410 6500 5414 6556
rect 5414 6500 5470 6556
rect 5470 6500 5474 6556
rect 5410 6496 5474 6500
rect 5490 6556 5554 6560
rect 5490 6500 5494 6556
rect 5494 6500 5550 6556
rect 5550 6500 5554 6556
rect 5490 6496 5554 6500
rect 5570 6556 5634 6560
rect 5570 6500 5574 6556
rect 5574 6500 5630 6556
rect 5630 6500 5634 6556
rect 5570 6496 5634 6500
rect 14664 6556 14728 6560
rect 14664 6500 14668 6556
rect 14668 6500 14724 6556
rect 14724 6500 14728 6556
rect 14664 6496 14728 6500
rect 14744 6556 14808 6560
rect 14744 6500 14748 6556
rect 14748 6500 14804 6556
rect 14804 6500 14808 6556
rect 14744 6496 14808 6500
rect 14824 6556 14888 6560
rect 14824 6500 14828 6556
rect 14828 6500 14884 6556
rect 14884 6500 14888 6556
rect 14824 6496 14888 6500
rect 14904 6556 14968 6560
rect 14904 6500 14908 6556
rect 14908 6500 14964 6556
rect 14964 6500 14968 6556
rect 14904 6496 14968 6500
rect 23997 6556 24061 6560
rect 23997 6500 24001 6556
rect 24001 6500 24057 6556
rect 24057 6500 24061 6556
rect 23997 6496 24061 6500
rect 24077 6556 24141 6560
rect 24077 6500 24081 6556
rect 24081 6500 24137 6556
rect 24137 6500 24141 6556
rect 24077 6496 24141 6500
rect 24157 6556 24221 6560
rect 24157 6500 24161 6556
rect 24161 6500 24217 6556
rect 24217 6500 24221 6556
rect 24157 6496 24221 6500
rect 24237 6556 24301 6560
rect 24237 6500 24241 6556
rect 24241 6500 24297 6556
rect 24297 6500 24301 6556
rect 24237 6496 24301 6500
rect 9997 6012 10061 6016
rect 9997 5956 10001 6012
rect 10001 5956 10057 6012
rect 10057 5956 10061 6012
rect 9997 5952 10061 5956
rect 10077 6012 10141 6016
rect 10077 5956 10081 6012
rect 10081 5956 10137 6012
rect 10137 5956 10141 6012
rect 10077 5952 10141 5956
rect 10157 6012 10221 6016
rect 10157 5956 10161 6012
rect 10161 5956 10217 6012
rect 10217 5956 10221 6012
rect 10157 5952 10221 5956
rect 10237 6012 10301 6016
rect 10237 5956 10241 6012
rect 10241 5956 10297 6012
rect 10297 5956 10301 6012
rect 10237 5952 10301 5956
rect 19330 6012 19394 6016
rect 19330 5956 19334 6012
rect 19334 5956 19390 6012
rect 19390 5956 19394 6012
rect 19330 5952 19394 5956
rect 19410 6012 19474 6016
rect 19410 5956 19414 6012
rect 19414 5956 19470 6012
rect 19470 5956 19474 6012
rect 19410 5952 19474 5956
rect 19490 6012 19554 6016
rect 19490 5956 19494 6012
rect 19494 5956 19550 6012
rect 19550 5956 19554 6012
rect 19490 5952 19554 5956
rect 19570 6012 19634 6016
rect 19570 5956 19574 6012
rect 19574 5956 19630 6012
rect 19630 5956 19634 6012
rect 19570 5952 19634 5956
rect 5330 5468 5394 5472
rect 5330 5412 5334 5468
rect 5334 5412 5390 5468
rect 5390 5412 5394 5468
rect 5330 5408 5394 5412
rect 5410 5468 5474 5472
rect 5410 5412 5414 5468
rect 5414 5412 5470 5468
rect 5470 5412 5474 5468
rect 5410 5408 5474 5412
rect 5490 5468 5554 5472
rect 5490 5412 5494 5468
rect 5494 5412 5550 5468
rect 5550 5412 5554 5468
rect 5490 5408 5554 5412
rect 5570 5468 5634 5472
rect 5570 5412 5574 5468
rect 5574 5412 5630 5468
rect 5630 5412 5634 5468
rect 5570 5408 5634 5412
rect 14664 5468 14728 5472
rect 14664 5412 14668 5468
rect 14668 5412 14724 5468
rect 14724 5412 14728 5468
rect 14664 5408 14728 5412
rect 14744 5468 14808 5472
rect 14744 5412 14748 5468
rect 14748 5412 14804 5468
rect 14804 5412 14808 5468
rect 14744 5408 14808 5412
rect 14824 5468 14888 5472
rect 14824 5412 14828 5468
rect 14828 5412 14884 5468
rect 14884 5412 14888 5468
rect 14824 5408 14888 5412
rect 14904 5468 14968 5472
rect 14904 5412 14908 5468
rect 14908 5412 14964 5468
rect 14964 5412 14968 5468
rect 14904 5408 14968 5412
rect 23997 5468 24061 5472
rect 23997 5412 24001 5468
rect 24001 5412 24057 5468
rect 24057 5412 24061 5468
rect 23997 5408 24061 5412
rect 24077 5468 24141 5472
rect 24077 5412 24081 5468
rect 24081 5412 24137 5468
rect 24137 5412 24141 5468
rect 24077 5408 24141 5412
rect 24157 5468 24221 5472
rect 24157 5412 24161 5468
rect 24161 5412 24217 5468
rect 24217 5412 24221 5468
rect 24157 5408 24221 5412
rect 24237 5468 24301 5472
rect 24237 5412 24241 5468
rect 24241 5412 24297 5468
rect 24297 5412 24301 5468
rect 24237 5408 24301 5412
rect 9997 4924 10061 4928
rect 9997 4868 10001 4924
rect 10001 4868 10057 4924
rect 10057 4868 10061 4924
rect 9997 4864 10061 4868
rect 10077 4924 10141 4928
rect 10077 4868 10081 4924
rect 10081 4868 10137 4924
rect 10137 4868 10141 4924
rect 10077 4864 10141 4868
rect 10157 4924 10221 4928
rect 10157 4868 10161 4924
rect 10161 4868 10217 4924
rect 10217 4868 10221 4924
rect 10157 4864 10221 4868
rect 10237 4924 10301 4928
rect 10237 4868 10241 4924
rect 10241 4868 10297 4924
rect 10297 4868 10301 4924
rect 10237 4864 10301 4868
rect 19330 4924 19394 4928
rect 19330 4868 19334 4924
rect 19334 4868 19390 4924
rect 19390 4868 19394 4924
rect 19330 4864 19394 4868
rect 19410 4924 19474 4928
rect 19410 4868 19414 4924
rect 19414 4868 19470 4924
rect 19470 4868 19474 4924
rect 19410 4864 19474 4868
rect 19490 4924 19554 4928
rect 19490 4868 19494 4924
rect 19494 4868 19550 4924
rect 19550 4868 19554 4924
rect 19490 4864 19554 4868
rect 19570 4924 19634 4928
rect 19570 4868 19574 4924
rect 19574 4868 19630 4924
rect 19630 4868 19634 4924
rect 19570 4864 19634 4868
rect 5330 4380 5394 4384
rect 5330 4324 5334 4380
rect 5334 4324 5390 4380
rect 5390 4324 5394 4380
rect 5330 4320 5394 4324
rect 5410 4380 5474 4384
rect 5410 4324 5414 4380
rect 5414 4324 5470 4380
rect 5470 4324 5474 4380
rect 5410 4320 5474 4324
rect 5490 4380 5554 4384
rect 5490 4324 5494 4380
rect 5494 4324 5550 4380
rect 5550 4324 5554 4380
rect 5490 4320 5554 4324
rect 5570 4380 5634 4384
rect 5570 4324 5574 4380
rect 5574 4324 5630 4380
rect 5630 4324 5634 4380
rect 5570 4320 5634 4324
rect 14664 4380 14728 4384
rect 14664 4324 14668 4380
rect 14668 4324 14724 4380
rect 14724 4324 14728 4380
rect 14664 4320 14728 4324
rect 14744 4380 14808 4384
rect 14744 4324 14748 4380
rect 14748 4324 14804 4380
rect 14804 4324 14808 4380
rect 14744 4320 14808 4324
rect 14824 4380 14888 4384
rect 14824 4324 14828 4380
rect 14828 4324 14884 4380
rect 14884 4324 14888 4380
rect 14824 4320 14888 4324
rect 14904 4380 14968 4384
rect 14904 4324 14908 4380
rect 14908 4324 14964 4380
rect 14964 4324 14968 4380
rect 14904 4320 14968 4324
rect 23997 4380 24061 4384
rect 23997 4324 24001 4380
rect 24001 4324 24057 4380
rect 24057 4324 24061 4380
rect 23997 4320 24061 4324
rect 24077 4380 24141 4384
rect 24077 4324 24081 4380
rect 24081 4324 24137 4380
rect 24137 4324 24141 4380
rect 24077 4320 24141 4324
rect 24157 4380 24221 4384
rect 24157 4324 24161 4380
rect 24161 4324 24217 4380
rect 24217 4324 24221 4380
rect 24157 4320 24221 4324
rect 24237 4380 24301 4384
rect 24237 4324 24241 4380
rect 24241 4324 24297 4380
rect 24297 4324 24301 4380
rect 24237 4320 24301 4324
rect 9997 3836 10061 3840
rect 9997 3780 10001 3836
rect 10001 3780 10057 3836
rect 10057 3780 10061 3836
rect 9997 3776 10061 3780
rect 10077 3836 10141 3840
rect 10077 3780 10081 3836
rect 10081 3780 10137 3836
rect 10137 3780 10141 3836
rect 10077 3776 10141 3780
rect 10157 3836 10221 3840
rect 10157 3780 10161 3836
rect 10161 3780 10217 3836
rect 10217 3780 10221 3836
rect 10157 3776 10221 3780
rect 10237 3836 10301 3840
rect 10237 3780 10241 3836
rect 10241 3780 10297 3836
rect 10297 3780 10301 3836
rect 10237 3776 10301 3780
rect 19330 3836 19394 3840
rect 19330 3780 19334 3836
rect 19334 3780 19390 3836
rect 19390 3780 19394 3836
rect 19330 3776 19394 3780
rect 19410 3836 19474 3840
rect 19410 3780 19414 3836
rect 19414 3780 19470 3836
rect 19470 3780 19474 3836
rect 19410 3776 19474 3780
rect 19490 3836 19554 3840
rect 19490 3780 19494 3836
rect 19494 3780 19550 3836
rect 19550 3780 19554 3836
rect 19490 3776 19554 3780
rect 19570 3836 19634 3840
rect 19570 3780 19574 3836
rect 19574 3780 19630 3836
rect 19630 3780 19634 3836
rect 19570 3776 19634 3780
rect 5330 3292 5394 3296
rect 5330 3236 5334 3292
rect 5334 3236 5390 3292
rect 5390 3236 5394 3292
rect 5330 3232 5394 3236
rect 5410 3292 5474 3296
rect 5410 3236 5414 3292
rect 5414 3236 5470 3292
rect 5470 3236 5474 3292
rect 5410 3232 5474 3236
rect 5490 3292 5554 3296
rect 5490 3236 5494 3292
rect 5494 3236 5550 3292
rect 5550 3236 5554 3292
rect 5490 3232 5554 3236
rect 5570 3292 5634 3296
rect 5570 3236 5574 3292
rect 5574 3236 5630 3292
rect 5630 3236 5634 3292
rect 5570 3232 5634 3236
rect 14664 3292 14728 3296
rect 14664 3236 14668 3292
rect 14668 3236 14724 3292
rect 14724 3236 14728 3292
rect 14664 3232 14728 3236
rect 14744 3292 14808 3296
rect 14744 3236 14748 3292
rect 14748 3236 14804 3292
rect 14804 3236 14808 3292
rect 14744 3232 14808 3236
rect 14824 3292 14888 3296
rect 14824 3236 14828 3292
rect 14828 3236 14884 3292
rect 14884 3236 14888 3292
rect 14824 3232 14888 3236
rect 14904 3292 14968 3296
rect 14904 3236 14908 3292
rect 14908 3236 14964 3292
rect 14964 3236 14968 3292
rect 14904 3232 14968 3236
rect 23997 3292 24061 3296
rect 23997 3236 24001 3292
rect 24001 3236 24057 3292
rect 24057 3236 24061 3292
rect 23997 3232 24061 3236
rect 24077 3292 24141 3296
rect 24077 3236 24081 3292
rect 24081 3236 24137 3292
rect 24137 3236 24141 3292
rect 24077 3232 24141 3236
rect 24157 3292 24221 3296
rect 24157 3236 24161 3292
rect 24161 3236 24217 3292
rect 24217 3236 24221 3292
rect 24157 3232 24221 3236
rect 24237 3292 24301 3296
rect 24237 3236 24241 3292
rect 24241 3236 24297 3292
rect 24297 3236 24301 3292
rect 24237 3232 24301 3236
rect 9997 2748 10061 2752
rect 9997 2692 10001 2748
rect 10001 2692 10057 2748
rect 10057 2692 10061 2748
rect 9997 2688 10061 2692
rect 10077 2748 10141 2752
rect 10077 2692 10081 2748
rect 10081 2692 10137 2748
rect 10137 2692 10141 2748
rect 10077 2688 10141 2692
rect 10157 2748 10221 2752
rect 10157 2692 10161 2748
rect 10161 2692 10217 2748
rect 10217 2692 10221 2748
rect 10157 2688 10221 2692
rect 10237 2748 10301 2752
rect 10237 2692 10241 2748
rect 10241 2692 10297 2748
rect 10297 2692 10301 2748
rect 10237 2688 10301 2692
rect 19330 2748 19394 2752
rect 19330 2692 19334 2748
rect 19334 2692 19390 2748
rect 19390 2692 19394 2748
rect 19330 2688 19394 2692
rect 19410 2748 19474 2752
rect 19410 2692 19414 2748
rect 19414 2692 19470 2748
rect 19470 2692 19474 2748
rect 19410 2688 19474 2692
rect 19490 2748 19554 2752
rect 19490 2692 19494 2748
rect 19494 2692 19550 2748
rect 19550 2692 19554 2748
rect 19490 2688 19554 2692
rect 19570 2748 19634 2752
rect 19570 2692 19574 2748
rect 19574 2692 19630 2748
rect 19630 2692 19634 2748
rect 19570 2688 19634 2692
rect 5330 2204 5394 2208
rect 5330 2148 5334 2204
rect 5334 2148 5390 2204
rect 5390 2148 5394 2204
rect 5330 2144 5394 2148
rect 5410 2204 5474 2208
rect 5410 2148 5414 2204
rect 5414 2148 5470 2204
rect 5470 2148 5474 2204
rect 5410 2144 5474 2148
rect 5490 2204 5554 2208
rect 5490 2148 5494 2204
rect 5494 2148 5550 2204
rect 5550 2148 5554 2204
rect 5490 2144 5554 2148
rect 5570 2204 5634 2208
rect 5570 2148 5574 2204
rect 5574 2148 5630 2204
rect 5630 2148 5634 2204
rect 5570 2144 5634 2148
rect 14664 2204 14728 2208
rect 14664 2148 14668 2204
rect 14668 2148 14724 2204
rect 14724 2148 14728 2204
rect 14664 2144 14728 2148
rect 14744 2204 14808 2208
rect 14744 2148 14748 2204
rect 14748 2148 14804 2204
rect 14804 2148 14808 2204
rect 14744 2144 14808 2148
rect 14824 2204 14888 2208
rect 14824 2148 14828 2204
rect 14828 2148 14884 2204
rect 14884 2148 14888 2204
rect 14824 2144 14888 2148
rect 14904 2204 14968 2208
rect 14904 2148 14908 2204
rect 14908 2148 14964 2204
rect 14964 2148 14968 2204
rect 14904 2144 14968 2148
rect 23997 2204 24061 2208
rect 23997 2148 24001 2204
rect 24001 2148 24057 2204
rect 24057 2148 24061 2204
rect 23997 2144 24061 2148
rect 24077 2204 24141 2208
rect 24077 2148 24081 2204
rect 24081 2148 24137 2204
rect 24137 2148 24141 2204
rect 24077 2144 24141 2148
rect 24157 2204 24221 2208
rect 24157 2148 24161 2204
rect 24161 2148 24217 2204
rect 24217 2148 24221 2204
rect 24157 2144 24221 2148
rect 24237 2204 24301 2208
rect 24237 2148 24241 2204
rect 24241 2148 24297 2204
rect 24297 2148 24301 2204
rect 24237 2144 24301 2148
<< metal4 >>
rect 5322 25056 5643 25616
rect 5322 24992 5330 25056
rect 5394 24992 5410 25056
rect 5474 24992 5490 25056
rect 5554 24992 5570 25056
rect 5634 24992 5643 25056
rect 5322 23968 5643 24992
rect 5322 23904 5330 23968
rect 5394 23904 5410 23968
rect 5474 23904 5490 23968
rect 5554 23904 5570 23968
rect 5634 23904 5643 23968
rect 5322 22880 5643 23904
rect 5322 22816 5330 22880
rect 5394 22816 5410 22880
rect 5474 22816 5490 22880
rect 5554 22816 5570 22880
rect 5634 22816 5643 22880
rect 5322 21792 5643 22816
rect 5322 21728 5330 21792
rect 5394 21728 5410 21792
rect 5474 21728 5490 21792
rect 5554 21728 5570 21792
rect 5634 21728 5643 21792
rect 5322 20704 5643 21728
rect 9989 25600 10309 25616
rect 9989 25536 9997 25600
rect 10061 25536 10077 25600
rect 10141 25536 10157 25600
rect 10221 25536 10237 25600
rect 10301 25536 10309 25600
rect 9989 24512 10309 25536
rect 9989 24448 9997 24512
rect 10061 24448 10077 24512
rect 10141 24448 10157 24512
rect 10221 24448 10237 24512
rect 10301 24448 10309 24512
rect 9989 23424 10309 24448
rect 9989 23360 9997 23424
rect 10061 23360 10077 23424
rect 10141 23360 10157 23424
rect 10221 23360 10237 23424
rect 10301 23360 10309 23424
rect 9989 22336 10309 23360
rect 9989 22272 9997 22336
rect 10061 22272 10077 22336
rect 10141 22272 10157 22336
rect 10221 22272 10237 22336
rect 10301 22272 10309 22336
rect 9989 21248 10309 22272
rect 9989 21184 9997 21248
rect 10061 21184 10077 21248
rect 10141 21184 10157 21248
rect 10221 21184 10237 21248
rect 10301 21184 10309 21248
rect 9339 20908 9405 20909
rect 9339 20844 9340 20908
rect 9404 20844 9405 20908
rect 9339 20843 9405 20844
rect 5322 20640 5330 20704
rect 5394 20640 5410 20704
rect 5474 20640 5490 20704
rect 5554 20640 5570 20704
rect 5634 20640 5643 20704
rect 5322 19616 5643 20640
rect 9342 20637 9402 20843
rect 9339 20636 9405 20637
rect 9339 20572 9340 20636
rect 9404 20572 9405 20636
rect 9339 20571 9405 20572
rect 5322 19552 5330 19616
rect 5394 19552 5410 19616
rect 5474 19552 5490 19616
rect 5554 19552 5570 19616
rect 5634 19552 5643 19616
rect 5322 18528 5643 19552
rect 5322 18464 5330 18528
rect 5394 18464 5410 18528
rect 5474 18464 5490 18528
rect 5554 18464 5570 18528
rect 5634 18464 5643 18528
rect 5322 17440 5643 18464
rect 5322 17376 5330 17440
rect 5394 17376 5410 17440
rect 5474 17376 5490 17440
rect 5554 17376 5570 17440
rect 5634 17376 5643 17440
rect 5322 16352 5643 17376
rect 5322 16288 5330 16352
rect 5394 16288 5410 16352
rect 5474 16288 5490 16352
rect 5554 16288 5570 16352
rect 5634 16288 5643 16352
rect 5322 15264 5643 16288
rect 5322 15200 5330 15264
rect 5394 15200 5410 15264
rect 5474 15200 5490 15264
rect 5554 15200 5570 15264
rect 5634 15200 5643 15264
rect 5322 14176 5643 15200
rect 5322 14112 5330 14176
rect 5394 14112 5410 14176
rect 5474 14112 5490 14176
rect 5554 14112 5570 14176
rect 5634 14112 5643 14176
rect 5322 13088 5643 14112
rect 5322 13024 5330 13088
rect 5394 13024 5410 13088
rect 5474 13024 5490 13088
rect 5554 13024 5570 13088
rect 5634 13024 5643 13088
rect 5322 12000 5643 13024
rect 5322 11936 5330 12000
rect 5394 11936 5410 12000
rect 5474 11936 5490 12000
rect 5554 11936 5570 12000
rect 5634 11936 5643 12000
rect 5322 10912 5643 11936
rect 5322 10848 5330 10912
rect 5394 10848 5410 10912
rect 5474 10848 5490 10912
rect 5554 10848 5570 10912
rect 5634 10848 5643 10912
rect 5322 9824 5643 10848
rect 5322 9760 5330 9824
rect 5394 9760 5410 9824
rect 5474 9760 5490 9824
rect 5554 9760 5570 9824
rect 5634 9760 5643 9824
rect 5322 8736 5643 9760
rect 5322 8672 5330 8736
rect 5394 8672 5410 8736
rect 5474 8672 5490 8736
rect 5554 8672 5570 8736
rect 5634 8672 5643 8736
rect 5322 7648 5643 8672
rect 5322 7584 5330 7648
rect 5394 7584 5410 7648
rect 5474 7584 5490 7648
rect 5554 7584 5570 7648
rect 5634 7584 5643 7648
rect 5322 6560 5643 7584
rect 5322 6496 5330 6560
rect 5394 6496 5410 6560
rect 5474 6496 5490 6560
rect 5554 6496 5570 6560
rect 5634 6496 5643 6560
rect 5322 5472 5643 6496
rect 5322 5408 5330 5472
rect 5394 5408 5410 5472
rect 5474 5408 5490 5472
rect 5554 5408 5570 5472
rect 5634 5408 5643 5472
rect 5322 4384 5643 5408
rect 5322 4320 5330 4384
rect 5394 4320 5410 4384
rect 5474 4320 5490 4384
rect 5554 4320 5570 4384
rect 5634 4320 5643 4384
rect 5322 3296 5643 4320
rect 5322 3232 5330 3296
rect 5394 3232 5410 3296
rect 5474 3232 5490 3296
rect 5554 3232 5570 3296
rect 5634 3232 5643 3296
rect 5322 2208 5643 3232
rect 5322 2144 5330 2208
rect 5394 2144 5410 2208
rect 5474 2144 5490 2208
rect 5554 2144 5570 2208
rect 5634 2144 5643 2208
rect 5322 2128 5643 2144
rect 9989 20160 10309 21184
rect 9989 20096 9997 20160
rect 10061 20096 10077 20160
rect 10141 20096 10157 20160
rect 10221 20096 10237 20160
rect 10301 20096 10309 20160
rect 9989 19072 10309 20096
rect 9989 19008 9997 19072
rect 10061 19008 10077 19072
rect 10141 19008 10157 19072
rect 10221 19008 10237 19072
rect 10301 19008 10309 19072
rect 9989 17984 10309 19008
rect 9989 17920 9997 17984
rect 10061 17920 10077 17984
rect 10141 17920 10157 17984
rect 10221 17920 10237 17984
rect 10301 17920 10309 17984
rect 9989 16896 10309 17920
rect 9989 16832 9997 16896
rect 10061 16832 10077 16896
rect 10141 16832 10157 16896
rect 10221 16832 10237 16896
rect 10301 16832 10309 16896
rect 9989 15808 10309 16832
rect 9989 15744 9997 15808
rect 10061 15744 10077 15808
rect 10141 15744 10157 15808
rect 10221 15744 10237 15808
rect 10301 15744 10309 15808
rect 9989 14720 10309 15744
rect 9989 14656 9997 14720
rect 10061 14656 10077 14720
rect 10141 14656 10157 14720
rect 10221 14656 10237 14720
rect 10301 14656 10309 14720
rect 9989 13632 10309 14656
rect 9989 13568 9997 13632
rect 10061 13568 10077 13632
rect 10141 13568 10157 13632
rect 10221 13568 10237 13632
rect 10301 13568 10309 13632
rect 9989 12544 10309 13568
rect 9989 12480 9997 12544
rect 10061 12480 10077 12544
rect 10141 12480 10157 12544
rect 10221 12480 10237 12544
rect 10301 12480 10309 12544
rect 9989 11456 10309 12480
rect 9989 11392 9997 11456
rect 10061 11392 10077 11456
rect 10141 11392 10157 11456
rect 10221 11392 10237 11456
rect 10301 11392 10309 11456
rect 9989 10368 10309 11392
rect 9989 10304 9997 10368
rect 10061 10304 10077 10368
rect 10141 10304 10157 10368
rect 10221 10304 10237 10368
rect 10301 10304 10309 10368
rect 9989 9280 10309 10304
rect 9989 9216 9997 9280
rect 10061 9216 10077 9280
rect 10141 9216 10157 9280
rect 10221 9216 10237 9280
rect 10301 9216 10309 9280
rect 9989 8192 10309 9216
rect 9989 8128 9997 8192
rect 10061 8128 10077 8192
rect 10141 8128 10157 8192
rect 10221 8128 10237 8192
rect 10301 8128 10309 8192
rect 9989 7104 10309 8128
rect 9989 7040 9997 7104
rect 10061 7040 10077 7104
rect 10141 7040 10157 7104
rect 10221 7040 10237 7104
rect 10301 7040 10309 7104
rect 9989 6016 10309 7040
rect 9989 5952 9997 6016
rect 10061 5952 10077 6016
rect 10141 5952 10157 6016
rect 10221 5952 10237 6016
rect 10301 5952 10309 6016
rect 9989 4928 10309 5952
rect 9989 4864 9997 4928
rect 10061 4864 10077 4928
rect 10141 4864 10157 4928
rect 10221 4864 10237 4928
rect 10301 4864 10309 4928
rect 9989 3840 10309 4864
rect 9989 3776 9997 3840
rect 10061 3776 10077 3840
rect 10141 3776 10157 3840
rect 10221 3776 10237 3840
rect 10301 3776 10309 3840
rect 9989 2752 10309 3776
rect 9989 2688 9997 2752
rect 10061 2688 10077 2752
rect 10141 2688 10157 2752
rect 10221 2688 10237 2752
rect 10301 2688 10309 2752
rect 9989 2128 10309 2688
rect 14656 25056 14976 25616
rect 14656 24992 14664 25056
rect 14728 24992 14744 25056
rect 14808 24992 14824 25056
rect 14888 24992 14904 25056
rect 14968 24992 14976 25056
rect 14656 23968 14976 24992
rect 14656 23904 14664 23968
rect 14728 23904 14744 23968
rect 14808 23904 14824 23968
rect 14888 23904 14904 23968
rect 14968 23904 14976 23968
rect 14656 22880 14976 23904
rect 14656 22816 14664 22880
rect 14728 22816 14744 22880
rect 14808 22816 14824 22880
rect 14888 22816 14904 22880
rect 14968 22816 14976 22880
rect 14656 21792 14976 22816
rect 14656 21728 14664 21792
rect 14728 21728 14744 21792
rect 14808 21728 14824 21792
rect 14888 21728 14904 21792
rect 14968 21728 14976 21792
rect 14656 20704 14976 21728
rect 14656 20640 14664 20704
rect 14728 20640 14744 20704
rect 14808 20640 14824 20704
rect 14888 20640 14904 20704
rect 14968 20640 14976 20704
rect 14656 19616 14976 20640
rect 14656 19552 14664 19616
rect 14728 19552 14744 19616
rect 14808 19552 14824 19616
rect 14888 19552 14904 19616
rect 14968 19552 14976 19616
rect 14656 18528 14976 19552
rect 14656 18464 14664 18528
rect 14728 18464 14744 18528
rect 14808 18464 14824 18528
rect 14888 18464 14904 18528
rect 14968 18464 14976 18528
rect 14656 17440 14976 18464
rect 14656 17376 14664 17440
rect 14728 17376 14744 17440
rect 14808 17376 14824 17440
rect 14888 17376 14904 17440
rect 14968 17376 14976 17440
rect 14656 16352 14976 17376
rect 14656 16288 14664 16352
rect 14728 16288 14744 16352
rect 14808 16288 14824 16352
rect 14888 16288 14904 16352
rect 14968 16288 14976 16352
rect 14656 15264 14976 16288
rect 14656 15200 14664 15264
rect 14728 15200 14744 15264
rect 14808 15200 14824 15264
rect 14888 15200 14904 15264
rect 14968 15200 14976 15264
rect 14656 14176 14976 15200
rect 14656 14112 14664 14176
rect 14728 14112 14744 14176
rect 14808 14112 14824 14176
rect 14888 14112 14904 14176
rect 14968 14112 14976 14176
rect 14656 13088 14976 14112
rect 14656 13024 14664 13088
rect 14728 13024 14744 13088
rect 14808 13024 14824 13088
rect 14888 13024 14904 13088
rect 14968 13024 14976 13088
rect 14656 12000 14976 13024
rect 14656 11936 14664 12000
rect 14728 11936 14744 12000
rect 14808 11936 14824 12000
rect 14888 11936 14904 12000
rect 14968 11936 14976 12000
rect 14656 10912 14976 11936
rect 14656 10848 14664 10912
rect 14728 10848 14744 10912
rect 14808 10848 14824 10912
rect 14888 10848 14904 10912
rect 14968 10848 14976 10912
rect 14656 9824 14976 10848
rect 14656 9760 14664 9824
rect 14728 9760 14744 9824
rect 14808 9760 14824 9824
rect 14888 9760 14904 9824
rect 14968 9760 14976 9824
rect 14656 8736 14976 9760
rect 14656 8672 14664 8736
rect 14728 8672 14744 8736
rect 14808 8672 14824 8736
rect 14888 8672 14904 8736
rect 14968 8672 14976 8736
rect 14656 7648 14976 8672
rect 14656 7584 14664 7648
rect 14728 7584 14744 7648
rect 14808 7584 14824 7648
rect 14888 7584 14904 7648
rect 14968 7584 14976 7648
rect 14656 6560 14976 7584
rect 14656 6496 14664 6560
rect 14728 6496 14744 6560
rect 14808 6496 14824 6560
rect 14888 6496 14904 6560
rect 14968 6496 14976 6560
rect 14656 5472 14976 6496
rect 14656 5408 14664 5472
rect 14728 5408 14744 5472
rect 14808 5408 14824 5472
rect 14888 5408 14904 5472
rect 14968 5408 14976 5472
rect 14656 4384 14976 5408
rect 14656 4320 14664 4384
rect 14728 4320 14744 4384
rect 14808 4320 14824 4384
rect 14888 4320 14904 4384
rect 14968 4320 14976 4384
rect 14656 3296 14976 4320
rect 14656 3232 14664 3296
rect 14728 3232 14744 3296
rect 14808 3232 14824 3296
rect 14888 3232 14904 3296
rect 14968 3232 14976 3296
rect 14656 2208 14976 3232
rect 14656 2144 14664 2208
rect 14728 2144 14744 2208
rect 14808 2144 14824 2208
rect 14888 2144 14904 2208
rect 14968 2144 14976 2208
rect 14656 2128 14976 2144
rect 19322 25600 19642 25616
rect 19322 25536 19330 25600
rect 19394 25536 19410 25600
rect 19474 25536 19490 25600
rect 19554 25536 19570 25600
rect 19634 25536 19642 25600
rect 19322 24512 19642 25536
rect 19322 24448 19330 24512
rect 19394 24448 19410 24512
rect 19474 24448 19490 24512
rect 19554 24448 19570 24512
rect 19634 24448 19642 24512
rect 19322 23424 19642 24448
rect 19322 23360 19330 23424
rect 19394 23360 19410 23424
rect 19474 23360 19490 23424
rect 19554 23360 19570 23424
rect 19634 23360 19642 23424
rect 19322 22336 19642 23360
rect 19322 22272 19330 22336
rect 19394 22272 19410 22336
rect 19474 22272 19490 22336
rect 19554 22272 19570 22336
rect 19634 22272 19642 22336
rect 19322 21248 19642 22272
rect 19322 21184 19330 21248
rect 19394 21184 19410 21248
rect 19474 21184 19490 21248
rect 19554 21184 19570 21248
rect 19634 21184 19642 21248
rect 19322 20160 19642 21184
rect 19322 20096 19330 20160
rect 19394 20096 19410 20160
rect 19474 20096 19490 20160
rect 19554 20096 19570 20160
rect 19634 20096 19642 20160
rect 19322 19072 19642 20096
rect 19322 19008 19330 19072
rect 19394 19008 19410 19072
rect 19474 19008 19490 19072
rect 19554 19008 19570 19072
rect 19634 19008 19642 19072
rect 19322 17984 19642 19008
rect 19322 17920 19330 17984
rect 19394 17920 19410 17984
rect 19474 17920 19490 17984
rect 19554 17920 19570 17984
rect 19634 17920 19642 17984
rect 19322 16896 19642 17920
rect 19322 16832 19330 16896
rect 19394 16832 19410 16896
rect 19474 16832 19490 16896
rect 19554 16832 19570 16896
rect 19634 16832 19642 16896
rect 19322 15808 19642 16832
rect 19322 15744 19330 15808
rect 19394 15744 19410 15808
rect 19474 15744 19490 15808
rect 19554 15744 19570 15808
rect 19634 15744 19642 15808
rect 19322 14720 19642 15744
rect 19322 14656 19330 14720
rect 19394 14656 19410 14720
rect 19474 14656 19490 14720
rect 19554 14656 19570 14720
rect 19634 14656 19642 14720
rect 19322 13632 19642 14656
rect 19322 13568 19330 13632
rect 19394 13568 19410 13632
rect 19474 13568 19490 13632
rect 19554 13568 19570 13632
rect 19634 13568 19642 13632
rect 19322 12544 19642 13568
rect 19322 12480 19330 12544
rect 19394 12480 19410 12544
rect 19474 12480 19490 12544
rect 19554 12480 19570 12544
rect 19634 12480 19642 12544
rect 19322 11456 19642 12480
rect 19322 11392 19330 11456
rect 19394 11392 19410 11456
rect 19474 11392 19490 11456
rect 19554 11392 19570 11456
rect 19634 11392 19642 11456
rect 19322 10368 19642 11392
rect 19322 10304 19330 10368
rect 19394 10304 19410 10368
rect 19474 10304 19490 10368
rect 19554 10304 19570 10368
rect 19634 10304 19642 10368
rect 19322 9280 19642 10304
rect 19322 9216 19330 9280
rect 19394 9216 19410 9280
rect 19474 9216 19490 9280
rect 19554 9216 19570 9280
rect 19634 9216 19642 9280
rect 19322 8192 19642 9216
rect 19322 8128 19330 8192
rect 19394 8128 19410 8192
rect 19474 8128 19490 8192
rect 19554 8128 19570 8192
rect 19634 8128 19642 8192
rect 19322 7104 19642 8128
rect 19322 7040 19330 7104
rect 19394 7040 19410 7104
rect 19474 7040 19490 7104
rect 19554 7040 19570 7104
rect 19634 7040 19642 7104
rect 19322 6016 19642 7040
rect 19322 5952 19330 6016
rect 19394 5952 19410 6016
rect 19474 5952 19490 6016
rect 19554 5952 19570 6016
rect 19634 5952 19642 6016
rect 19322 4928 19642 5952
rect 19322 4864 19330 4928
rect 19394 4864 19410 4928
rect 19474 4864 19490 4928
rect 19554 4864 19570 4928
rect 19634 4864 19642 4928
rect 19322 3840 19642 4864
rect 19322 3776 19330 3840
rect 19394 3776 19410 3840
rect 19474 3776 19490 3840
rect 19554 3776 19570 3840
rect 19634 3776 19642 3840
rect 19322 2752 19642 3776
rect 19322 2688 19330 2752
rect 19394 2688 19410 2752
rect 19474 2688 19490 2752
rect 19554 2688 19570 2752
rect 19634 2688 19642 2752
rect 19322 2128 19642 2688
rect 23989 25056 24309 25616
rect 23989 24992 23997 25056
rect 24061 24992 24077 25056
rect 24141 24992 24157 25056
rect 24221 24992 24237 25056
rect 24301 24992 24309 25056
rect 23989 23968 24309 24992
rect 23989 23904 23997 23968
rect 24061 23904 24077 23968
rect 24141 23904 24157 23968
rect 24221 23904 24237 23968
rect 24301 23904 24309 23968
rect 23989 22880 24309 23904
rect 23989 22816 23997 22880
rect 24061 22816 24077 22880
rect 24141 22816 24157 22880
rect 24221 22816 24237 22880
rect 24301 22816 24309 22880
rect 23989 21792 24309 22816
rect 23989 21728 23997 21792
rect 24061 21728 24077 21792
rect 24141 21728 24157 21792
rect 24221 21728 24237 21792
rect 24301 21728 24309 21792
rect 23989 20704 24309 21728
rect 23989 20640 23997 20704
rect 24061 20640 24077 20704
rect 24141 20640 24157 20704
rect 24221 20640 24237 20704
rect 24301 20640 24309 20704
rect 23989 19616 24309 20640
rect 23989 19552 23997 19616
rect 24061 19552 24077 19616
rect 24141 19552 24157 19616
rect 24221 19552 24237 19616
rect 24301 19552 24309 19616
rect 23989 18528 24309 19552
rect 23989 18464 23997 18528
rect 24061 18464 24077 18528
rect 24141 18464 24157 18528
rect 24221 18464 24237 18528
rect 24301 18464 24309 18528
rect 23989 17440 24309 18464
rect 23989 17376 23997 17440
rect 24061 17376 24077 17440
rect 24141 17376 24157 17440
rect 24221 17376 24237 17440
rect 24301 17376 24309 17440
rect 23989 16352 24309 17376
rect 23989 16288 23997 16352
rect 24061 16288 24077 16352
rect 24141 16288 24157 16352
rect 24221 16288 24237 16352
rect 24301 16288 24309 16352
rect 23989 15264 24309 16288
rect 23989 15200 23997 15264
rect 24061 15200 24077 15264
rect 24141 15200 24157 15264
rect 24221 15200 24237 15264
rect 24301 15200 24309 15264
rect 23989 14176 24309 15200
rect 23989 14112 23997 14176
rect 24061 14112 24077 14176
rect 24141 14112 24157 14176
rect 24221 14112 24237 14176
rect 24301 14112 24309 14176
rect 23989 13088 24309 14112
rect 23989 13024 23997 13088
rect 24061 13024 24077 13088
rect 24141 13024 24157 13088
rect 24221 13024 24237 13088
rect 24301 13024 24309 13088
rect 23989 12000 24309 13024
rect 23989 11936 23997 12000
rect 24061 11936 24077 12000
rect 24141 11936 24157 12000
rect 24221 11936 24237 12000
rect 24301 11936 24309 12000
rect 23989 10912 24309 11936
rect 23989 10848 23997 10912
rect 24061 10848 24077 10912
rect 24141 10848 24157 10912
rect 24221 10848 24237 10912
rect 24301 10848 24309 10912
rect 23989 9824 24309 10848
rect 23989 9760 23997 9824
rect 24061 9760 24077 9824
rect 24141 9760 24157 9824
rect 24221 9760 24237 9824
rect 24301 9760 24309 9824
rect 23989 8736 24309 9760
rect 23989 8672 23997 8736
rect 24061 8672 24077 8736
rect 24141 8672 24157 8736
rect 24221 8672 24237 8736
rect 24301 8672 24309 8736
rect 23989 7648 24309 8672
rect 23989 7584 23997 7648
rect 24061 7584 24077 7648
rect 24141 7584 24157 7648
rect 24221 7584 24237 7648
rect 24301 7584 24309 7648
rect 23989 6560 24309 7584
rect 23989 6496 23997 6560
rect 24061 6496 24077 6560
rect 24141 6496 24157 6560
rect 24221 6496 24237 6560
rect 24301 6496 24309 6560
rect 23989 5472 24309 6496
rect 23989 5408 23997 5472
rect 24061 5408 24077 5472
rect 24141 5408 24157 5472
rect 24221 5408 24237 5472
rect 24301 5408 24309 5472
rect 23989 4384 24309 5408
rect 23989 4320 23997 4384
rect 24061 4320 24077 4384
rect 24141 4320 24157 4384
rect 24221 4320 24237 4384
rect 24301 4320 24309 4384
rect 23989 3296 24309 4320
rect 23989 3232 23997 3296
rect 24061 3232 24077 3296
rect 24141 3232 24157 3296
rect 24221 3232 24237 3296
rect 24301 3232 24309 3296
rect 23989 2208 24309 3232
rect 23989 2144 23997 2208
rect 24061 2144 24077 2208
rect 24141 2144 24157 2208
rect 24221 2144 24237 2208
rect 24301 2144 24309 2208
rect 23989 2128 24309 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 816 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 816 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1092 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2196 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2196 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3668 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3300 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 3760 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3300 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4404 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 4864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5968 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5508 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6244 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6520 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6428 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6612 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 7716 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6520 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7624 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9372 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 8820 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9464 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 8728 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 9832 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11672 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 10936 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12224 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12040 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12316 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12132 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13236 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15076 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14524 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15168 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14340 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16272 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15444 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16548 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 17928 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17652 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17376 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18020 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 17744 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 18848 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _35_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20872 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20780 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19124 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20228 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 19952 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _27_
timestamp 1586364061
transform 1 0 22528 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__35__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21424 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_222
timestamp 1586364061
transform 1 0 21240 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_226
timestamp 1586364061
transform 1 0 21608 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_234
timestamp 1586364061
transform 1 0 22344 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21056 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22160 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_244
timestamp 1586364061
transform 1 0 23264 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 22896 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__27__A
timestamp 1586364061
transform 1 0 23080 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23264 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_245
timestamp 1586364061
transform 1 0 23356 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 23724 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23632 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _30_
timestamp 1586364061
transform 1 0 23632 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_257
timestamp 1586364061
transform 1 0 24460 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_252
timestamp 1586364061
transform 1 0 24000 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__28__A
timestamp 1586364061
transform 1 0 24276 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _31_
timestamp 1586364061
transform 1 0 24276 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_264
timestamp 1586364061
transform 1 0 25104 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24644 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__31__A
timestamp 1586364061
transform 1 0 24828 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__29__A
timestamp 1586364061
transform 1 0 25288 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _29_
timestamp 1586364061
transform 1 0 24736 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_276 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26208 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_1_268
timestamp 1586364061
transform 1 0 25472 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26116 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26576 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26576 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_263
timestamp 1586364061
transform 1 0 25012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 816 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3668 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3300 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 3760 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 4864 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 5968 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7072 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9280 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8176 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9372 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10476 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11580 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12684 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 14892 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 13788 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 14984 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16088 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17192 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18296 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20504 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19400 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20596 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21700 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _28_
timestamp 1586364061
transform 1 0 24276 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__30__A
timestamp 1586364061
transform 1 0 23632 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_239
timestamp 1586364061
transform 1 0 22804 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_247
timestamp 1586364061
transform 1 0 23540 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_250
timestamp 1586364061
transform 1 0 23816 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_254
timestamp 1586364061
transform 1 0 24184 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26576 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26116 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_259
timestamp 1586364061
transform 1 0 24644 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_271
timestamp 1586364061
transform 1 0 25748 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26208 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 816 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3300 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4404 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5508 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6244 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6428 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6520 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7624 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 8728 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 9832 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 10936 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12040 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12132 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13236 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14340 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15444 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16548 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17652 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 17744 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 18848 0 1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 20688 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20504 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_208
timestamp 1586364061
transform 1 0 19952 0 1 3808
box -38 -48 590 592
use scs8hd_buf_2  _32_
timestamp 1586364061
transform 1 0 21792 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 21240 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 22344 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_220
timestamp 1586364061
transform 1 0 21056 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_224
timestamp 1586364061
transform 1 0 21424 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_232
timestamp 1586364061
transform 1 0 22160 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_236
timestamp 1586364061
transform 1 0 22528 0 1 3808
box -38 -48 774 592
use scs8hd_buf_2  _26_
timestamp 1586364061
transform 1 0 24276 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23264 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 24092 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_245
timestamp 1586364061
transform 1 0 23356 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26576 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__26__A
timestamp 1586364061
transform 1 0 24828 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_259
timestamp 1586364061
transform 1 0 24644 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_263
timestamp 1586364061
transform 1 0 25012 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_3_275
timestamp 1586364061
transform 1 0 26116 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 816 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2196 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3668 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3300 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 3760 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 4864 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 5968 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7072 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9280 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8176 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9372 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10476 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11580 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12684 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 14892 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 13788 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 14984 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16088 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17192 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18296 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_track_25.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20688 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20504 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19400 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_215
timestamp 1586364061
transform 1 0 20596 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21240 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21608 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21976 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_219
timestamp 1586364061
transform 1 0 20964 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_224
timestamp 1586364061
transform 1 0 21424 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_228
timestamp 1586364061
transform 1 0 21792 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_232
timestamp 1586364061
transform 1 0 22160 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _33_
timestamp 1586364061
transform 1 0 24276 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_244
timestamp 1586364061
transform 1 0 23264 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_252
timestamp 1586364061
transform 1 0 24000 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26576 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26116 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_259
timestamp 1586364061
transform 1 0 24644 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_271
timestamp 1586364061
transform 1 0 25748 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26208 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 816 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3300 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4404 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5508 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6244 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6428 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6520 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7624 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 8728 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 9832 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 10936 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12040 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12132 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13236 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14340 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 16916 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15444 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_171
timestamp 1586364061
transform 1 0 16548 0 1 4896
box -38 -48 406 592
use scs8hd_decap_6  FILLER_5_177
timestamp 1586364061
transform 1 0 17100 0 1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17652 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18020 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_184
timestamp 1586364061
transform 1 0 17744 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_189
timestamp 1586364061
transform 1 0 18204 0 1 4896
box -38 -48 1142 592
use scs8hd_conb_1  _09_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20228 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 19308 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20044 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_203
timestamp 1586364061
transform 1 0 19492 0 1 4896
box -38 -48 590 592
use scs8hd_decap_4  FILLER_5_214
timestamp 1586364061
transform 1 0 20504 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_218
timestamp 1586364061
transform 1 0 20872 0 1 4896
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l2_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21240 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20964 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22252 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_221
timestamp 1586364061
transform 1 0 21148 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_231
timestamp 1586364061
transform 1 0 22068 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_235
timestamp 1586364061
transform 1 0 22436 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23264 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_243
timestamp 1586364061
transform 1 0 23172 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23356 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24460 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26576 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25564 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 816 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 816 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1092 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2196 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3668 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3300 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 3760 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3300 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4404 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 4864 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 5968 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5508 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6244 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6428 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7072 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6520 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7624 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9280 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8176 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9372 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 8728 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 9832 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10476 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11580 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 10936 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12040 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12684 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12132 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13236 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 14892 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 13788 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 14984 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14340 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 16916 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_6_166
timestamp 1586364061
transform 1 0 16088 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_174
timestamp 1586364061
transform 1 0 16824 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15444 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16548 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_184
timestamp 1586364061
transform 1 0 17744 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_179
timestamp 1586364061
transform 1 0 17284 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 17928 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17652 0 1 5984
box -38 -48 130 592
use scs8hd_buf_1  mux_bottom_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18020 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_188
timestamp 1586364061
transform 1 0 18112 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_196
timestamp 1586364061
transform 1 0 18848 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_190
timestamp 1586364061
transform 1 0 18296 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18388 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 18572 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 18940 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18940 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_205
timestamp 1586364061
transform 1 0 19676 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_201
timestamp 1586364061
transform 1 0 19308 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_205
timestamp 1586364061
transform 1 0 19676 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_199
timestamp 1586364061
transform 1 0 19124 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19492 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19952 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 19124 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 19308 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_215
timestamp 1586364061
transform 1 0 20596 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_212
timestamp 1586364061
transform 1 0 20320 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_209
timestamp 1586364061
transform 1 0 20044 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20136 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20504 0 -1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20136 0 1 5984
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20964 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 22068 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_228
timestamp 1586364061
transform 1 0 21792 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_229
timestamp 1586364061
transform 1 0 21884 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_233
timestamp 1586364061
transform 1 0 22252 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23264 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_240
timestamp 1586364061
transform 1 0 22896 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_252
timestamp 1586364061
transform 1 0 24000 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_241
timestamp 1586364061
transform 1 0 22988 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23356 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24460 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26576 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26576 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26116 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_264
timestamp 1586364061
transform 1 0 25104 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 25840 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26208 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25564 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 816 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2196 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3668 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3300 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 3760 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 4864 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 5968 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7072 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9280 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8176 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9372 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10476 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11580 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12684 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 14892 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 13788 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 14984 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16088 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_178
timestamp 1586364061
transform 1 0 17192 0 -1 7072
box -38 -48 590 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 17836 0 -1 7072
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18940 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_1  FILLER_8_184
timestamp 1586364061
transform 1 0 17744 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_189
timestamp 1586364061
transform 1 0 18204 0 -1 7072
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20872 0 -1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20504 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20136 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_206
timestamp 1586364061
transform 1 0 19768 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_212
timestamp 1586364061
transform 1 0 20320 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_215
timestamp 1586364061
transform 1 0 20596 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_237
timestamp 1586364061
transform 1 0 22620 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_249
timestamp 1586364061
transform 1 0 23724 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26576 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26116 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_261
timestamp 1586364061
transform 1 0 24828 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_273
timestamp 1586364061
transform 1 0 25932 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26208 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 816 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1092 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2196 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3300 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4404 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5508 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6244 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6428 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6520 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7624 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 8728 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 9832 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 10936 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12040 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12132 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13236 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14340 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 15720 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 16272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16640 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_159
timestamp 1586364061
transform 1 0 15444 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_166
timestamp 1586364061
transform 1 0 16088 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_170
timestamp 1586364061
transform 1 0 16456 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_174
timestamp 1586364061
transform 1 0 16824 0 1 7072
box -38 -48 774 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 17744 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17652 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 18296 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19032 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17560 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_188
timestamp 1586364061
transform 1 0 18112 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_192
timestamp 1586364061
transform 1 0 18480 0 1 7072
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19584 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19400 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_200
timestamp 1586364061
transform 1 0 19216 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21516 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21884 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22252 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_223
timestamp 1586364061
transform 1 0 21332 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_227
timestamp 1586364061
transform 1 0 21700 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_231
timestamp 1586364061
transform 1 0 22068 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_235
timestamp 1586364061
transform 1 0 22436 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23264 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23172 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23356 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24460 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26576 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25564 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 816 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2196 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3668 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3300 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 3760 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 4864 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 5968 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7072 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9280 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8176 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9372 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10476 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11580 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12684 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 14892 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 13788 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 14984 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16640 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_166
timestamp 1586364061
transform 1 0 16088 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_175
timestamp 1586364061
transform 1 0 16916 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18388 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_187
timestamp 1586364061
transform 1 0 18020 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_6  FILLER_10_193
timestamp 1586364061
transform 1 0 18572 0 -1 8160
box -38 -48 590 592
use scs8hd_conb_1  _11_
timestamp 1586364061
transform 1 0 19216 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20596 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20504 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_199
timestamp 1586364061
transform 1 0 19124 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_203
timestamp 1586364061
transform 1 0 19492 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_211
timestamp 1586364061
transform 1 0 20228 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_224
timestamp 1586364061
transform 1 0 21424 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_236
timestamp 1586364061
transform 1 0 22528 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_248
timestamp 1586364061
transform 1 0 23632 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26576 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26116 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_260
timestamp 1586364061
transform 1 0 24736 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_10_272
timestamp 1586364061
transform 1 0 25840 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26208 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 816 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1092 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2196 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3300 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4404 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5508 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6244 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6428 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6520 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7624 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 8728 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 9832 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 10936 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12040 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12132 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_135
timestamp 1586364061
transform 1 0 13236 0 1 8160
box -38 -48 590 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 13788 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 14340 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_145
timestamp 1586364061
transform 1 0 14156 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_149
timestamp 1586364061
transform 1 0 14524 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 15904 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_161
timestamp 1586364061
transform 1 0 15628 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_166
timestamp 1586364061
transform 1 0 16088 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_11_178
timestamp 1586364061
transform 1 0 17192 0 1 8160
box -38 -48 406 592
use scs8hd_conb_1  _10_
timestamp 1586364061
transform 1 0 18112 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17652 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18940 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18572 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17928 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_182
timestamp 1586364061
transform 1 0 17560 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_184
timestamp 1586364061
transform 1 0 17744 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_191
timestamp 1586364061
transform 1 0 18388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_195
timestamp 1586364061
transform 1 0 18756 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19124 0 1 8160
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_11_218
timestamp 1586364061
transform 1 0 20872 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_230
timestamp 1586364061
transform 1 0 21976 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23264 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_242
timestamp 1586364061
transform 1 0 23080 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23356 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24460 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26576 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25564 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 816 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2196 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3668 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3300 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 3760 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 4864 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 5968 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7072 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9280 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8176 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9372 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10476 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11580 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12684 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 14892 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 13788 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_154
timestamp 1586364061
transform 1 0 14984 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 15904 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_162
timestamp 1586364061
transform 1 0 15720 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_168
timestamp 1586364061
transform 1 0 16272 0 -1 9248
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18388 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_180
timestamp 1586364061
transform 1 0 17376 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_188
timestamp 1586364061
transform 1 0 18112 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20504 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19400 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20780 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_200
timestamp 1586364061
transform 1 0 19216 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_204
timestamp 1586364061
transform 1 0 19584 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_212
timestamp 1586364061
transform 1 0 20320 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_215
timestamp 1586364061
transform 1 0 20596 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_219
timestamp 1586364061
transform 1 0 20964 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_231
timestamp 1586364061
transform 1 0 22068 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_243
timestamp 1586364061
transform 1 0 23172 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_255
timestamp 1586364061
transform 1 0 24276 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26576 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26116 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_267
timestamp 1586364061
transform 1 0 25380 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26208 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 816 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 816 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1092 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2196 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2196 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3668 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3300 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4404 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3300 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 3760 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5508 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6244 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 4864 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 5968 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6428 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6520 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7624 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7072 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9280 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 8728 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 9832 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8176 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9372 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 10936 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10476 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11580 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12040 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12132 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13236 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12684 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14340 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 14892 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_150
timestamp 1586364061
transform 1 0 14616 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_154
timestamp 1586364061
transform 1 0 14984 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 13788 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 14984 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_166
timestamp 1586364061
transform 1 0 16088 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_13_178
timestamp 1586364061
transform 1 0 17192 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16088 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17192 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_188
timestamp 1586364061
transform 1 0 18112 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 17744 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17560 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17928 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17652 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_192
timestamp 1586364061
transform 1 0 18480 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_192
timestamp 1586364061
transform 1 0 18480 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18296 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18664 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18296 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18664 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18848 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18848 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20596 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20504 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20780 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20320 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_215
timestamp 1586364061
transform 1 0 20596 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_205
timestamp 1586364061
transform 1 0 19676 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_211
timestamp 1586364061
transform 1 0 20228 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21148 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21608 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_219
timestamp 1586364061
transform 1 0 20964 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_223
timestamp 1586364061
transform 1 0 21332 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_235
timestamp 1586364061
transform 1 0 22436 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_224
timestamp 1586364061
transform 1 0 21424 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_228
timestamp 1586364061
transform 1 0 21792 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23264 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 23172 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23356 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24460 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_240
timestamp 1586364061
transform 1 0 22896 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_252
timestamp 1586364061
transform 1 0 24000 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26576 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26576 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26116 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25564 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_264
timestamp 1586364061
transform 1 0 25104 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_272
timestamp 1586364061
transform 1 0 25840 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26208 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 816 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1092 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2196 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3300 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4404 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5508 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6244 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6428 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6520 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7624 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 8728 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 9832 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 10936 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12040 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12132 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13236 0 1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 14616 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 15168 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_147
timestamp 1586364061
transform 1 0 14340 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_154
timestamp 1586364061
transform 1 0 14984 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_158
timestamp 1586364061
transform 1 0 15352 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_170
timestamp 1586364061
transform 1 0 16456 0 1 10336
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19032 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17652 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18848 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18480 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_182
timestamp 1586364061
transform 1 0 17560 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_184
timestamp 1586364061
transform 1 0 17744 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_194
timestamp 1586364061
transform 1 0 18664 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_217
timestamp 1586364061
transform 1 0 20780 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21516 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21332 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20964 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_221
timestamp 1586364061
transform 1 0 21148 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_234
timestamp 1586364061
transform 1 0 22344 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23264 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_242
timestamp 1586364061
transform 1 0 23080 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23356 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24460 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26576 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25564 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 816 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2196 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3668 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3300 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 3760 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 4864 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 5968 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7072 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9280 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8176 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9372 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10476 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11580 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12684 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 14892 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14708 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_141
timestamp 1586364061
transform 1 0 13788 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_149
timestamp 1586364061
transform 1 0 14524 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 14984 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16088 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_178
timestamp 1586364061
transform 1 0 17192 0 -1 11424
box -38 -48 590 592
use scs8hd_conb_1  _08_
timestamp 1586364061
transform 1 0 18940 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17744 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18756 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18112 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_186
timestamp 1586364061
transform 1 0 17928 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_190
timestamp 1586364061
transform 1 0 18296 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_194
timestamp 1586364061
transform 1 0 18664 0 -1 11424
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20596 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20504 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19400 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20320 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19768 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_200
timestamp 1586364061
transform 1 0 19216 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_204
timestamp 1586364061
transform 1 0 19584 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_208
timestamp 1586364061
transform 1 0 19952 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_234
timestamp 1586364061
transform 1 0 22344 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_246
timestamp 1586364061
transform 1 0 23448 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26576 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26116 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_258
timestamp 1586364061
transform 1 0 24552 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_270
timestamp 1586364061
transform 1 0 25656 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26024 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26208 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 816 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1092 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2196 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3300 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4404 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5508 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6244 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6428 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6520 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7624 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 8728 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 9832 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 10936 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12040 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12132 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_17_135
timestamp 1586364061
transform 1 0 13236 0 1 11424
box -38 -48 406 592
use scs8hd_conb_1  _12_
timestamp 1586364061
transform 1 0 13696 0 1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 14708 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14524 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14156 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_139
timestamp 1586364061
transform 1 0 13604 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_143
timestamp 1586364061
transform 1 0 13972 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_147
timestamp 1586364061
transform 1 0 14340 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _14_
timestamp 1586364061
transform 1 0 16272 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16732 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17100 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__24__A
timestamp 1586364061
transform 1 0 15720 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_160
timestamp 1586364061
transform 1 0 15536 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_164
timestamp 1586364061
transform 1 0 15904 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_171
timestamp 1586364061
transform 1 0 16548 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 16916 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 17744 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17652 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17468 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18848 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17284 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_193
timestamp 1586364061
transform 1 0 18572 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_198
timestamp 1586364061
transform 1 0 19032 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19400 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19216 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21332 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21700 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 22068 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_221
timestamp 1586364061
transform 1 0 21148 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_225
timestamp 1586364061
transform 1 0 21516 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_229
timestamp 1586364061
transform 1 0 21884 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_233
timestamp 1586364061
transform 1 0 22252 0 1 11424
box -38 -48 774 592
use scs8hd_buf_2  _25_
timestamp 1586364061
transform 1 0 24276 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23264 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_241
timestamp 1586364061
transform 1 0 22988 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_245
timestamp 1586364061
transform 1 0 23356 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_253
timestamp 1586364061
transform 1 0 24092 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26576 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__25__A
timestamp 1586364061
transform 1 0 24828 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_259
timestamp 1586364061
transform 1 0 24644 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_263
timestamp 1586364061
transform 1 0 25012 0 1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_17_275
timestamp 1586364061
transform 1 0 26116 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 816 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3668 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3300 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 3760 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 4864 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 5968 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7072 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9280 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8176 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9372 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10476 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_117
timestamp 1586364061
transform 1 0 11580 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12408 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_125
timestamp 1586364061
transform 1 0 12316 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_128
timestamp 1586364061
transform 1 0 12592 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_136
timestamp 1586364061
transform 1 0 13328 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_141
timestamp 1586364061
transform 1 0 13788 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13604 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  mux_right_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13880 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14156 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14340 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14524 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14708 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 14892 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_154
timestamp 1586364061
transform 1 0 14984 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _24_
timestamp 1586364061
transform 1 0 15168 0 -1 12512
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16272 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15720 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_160
timestamp 1586364061
transform 1 0 15536 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_164
timestamp 1586364061
transform 1 0 15904 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18848 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_187
timestamp 1586364061
transform 1 0 18020 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_195
timestamp 1586364061
transform 1 0 18756 0 -1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20596 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20504 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_205
timestamp 1586364061
transform 1 0 19676 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_213
timestamp 1586364061
transform 1 0 20412 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_224
timestamp 1586364061
transform 1 0 21424 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_236
timestamp 1586364061
transform 1 0 22528 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_248
timestamp 1586364061
transform 1 0 23632 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26576 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26116 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_260
timestamp 1586364061
transform 1 0 24736 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_18_272
timestamp 1586364061
transform 1 0 25840 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26208 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 816 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 816 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1092 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2196 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2196 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3668 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3300 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4404 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3300 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 3760 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5508 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6244 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 4864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 5968 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6428 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6520 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7624 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7072 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9280 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 8728 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 9832 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8176 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9372 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 10936 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10476 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_117
timestamp 1586364061
transform 1 0 11580 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_125
timestamp 1586364061
transform 1 0 12316 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_127
timestamp 1586364061
transform 1 0 12500 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12040 0 1 12512
box -38 -48 130 592
use scs8hd_buf_2  _23_
timestamp 1586364061
transform 1 0 12132 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_135
timestamp 1586364061
transform 1 0 13236 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_131
timestamp 1586364061
transform 1 0 12868 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13052 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13420 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 12684 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12408 0 -1 13600
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 14156 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_148
timestamp 1586364061
transform 1 0 14432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14340 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13604 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_149
timestamp 1586364061
transform 1 0 14524 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_152
timestamp 1586364061
transform 1 0 14800 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14708 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14616 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14984 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 14892 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14984 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15168 0 1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15996 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_175
timestamp 1586364061
transform 1 0 16916 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_163
timestamp 1586364061
transform 1 0 15812 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_167
timestamp 1586364061
transform 1 0 16180 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_179
timestamp 1586364061
transform 1 0 17284 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_188
timestamp 1586364061
transform 1 0 18112 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_184
timestamp 1586364061
transform 1 0 17744 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_182
timestamp 1586364061
transform 1 0 17560 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_179
timestamp 1586364061
transform 1 0 17284 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17376 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17652 0 1 12512
box -38 -48 130 592
use scs8hd_conb_1  _15_
timestamp 1586364061
transform 1 0 17836 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_196
timestamp 1586364061
transform 1 0 18848 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_192
timestamp 1586364061
transform 1 0 18480 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18296 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18664 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19032 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17376 0 -1 13600
box -38 -48 1786 592
use scs8hd_conb_1  _13_
timestamp 1586364061
transform 1 0 20596 0 -1 13600
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19216 0 1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20504 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19308 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_199
timestamp 1586364061
transform 1 0 19124 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_203
timestamp 1586364061
transform 1 0 19492 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_20_211
timestamp 1586364061
transform 1 0 20228 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 20872 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_219
timestamp 1586364061
transform 1 0 20964 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_231
timestamp 1586364061
transform 1 0 22068 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 21976 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_1  mux_right_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23172 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23264 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23540 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_243
timestamp 1586364061
transform 1 0 23172 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23356 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_249
timestamp 1586364061
transform 1 0 23724 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_242
timestamp 1586364061
transform 1 0 23080 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_246
timestamp 1586364061
transform 1 0 23448 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26576 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26576 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26116 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_261
timestamp 1586364061
transform 1 0 24828 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_19_273
timestamp 1586364061
transform 1 0 25932 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_258
timestamp 1586364061
transform 1 0 24552 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_270
timestamp 1586364061
transform 1 0 25656 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26024 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26208 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 816 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1092 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2196 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3300 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4404 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5508 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6244 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6428 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6520 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7624 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 8728 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 9832 0 1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 11028 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_110
timestamp 1586364061
transform 1 0 10936 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_113
timestamp 1586364061
transform 1 0 11212 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12040 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12408 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 11948 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_123
timestamp 1586364061
transform 1 0 12132 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_128
timestamp 1586364061
transform 1 0 12592 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_132
timestamp 1586364061
transform 1 0 12960 0 1 13600
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14248 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14064 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13696 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_142
timestamp 1586364061
transform 1 0 13880 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16180 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17100 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16548 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_165
timestamp 1586364061
transform 1 0 15996 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_169
timestamp 1586364061
transform 1 0 16364 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_173
timestamp 1586364061
transform 1 0 16732 0 1 13600
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18388 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17652 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18204 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17468 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17284 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_184
timestamp 1586364061
transform 1 0 17744 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_188
timestamp 1586364061
transform 1 0 18112 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_210
timestamp 1586364061
transform 1 0 20136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_222
timestamp 1586364061
transform 1 0 21240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_234
timestamp 1586364061
transform 1 0 22344 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23264 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 24276 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_242
timestamp 1586364061
transform 1 0 23080 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_245
timestamp 1586364061
transform 1 0 23356 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_253
timestamp 1586364061
transform 1 0 24092 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24460 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26576 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25564 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 816 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2196 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3668 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3300 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 3760 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 4864 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 5968 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7072 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9280 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8176 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9372 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 11028 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_6  FILLER_22_105
timestamp 1586364061
transform 1 0 10476 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_8  FILLER_22_115
timestamp 1586364061
transform 1 0 11396 0 -1 14688
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12408 0 -1 14688
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_22_123
timestamp 1586364061
transform 1 0 12132 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 14892 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_145
timestamp 1586364061
transform 1 0 14156 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_6  FILLER_22_154
timestamp 1586364061
transform 1 0 14984 0 -1 14688
box -38 -48 590 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15628 0 -1 14688
box -38 -48 866 592
use scs8hd_fill_1  FILLER_22_160
timestamp 1586364061
transform 1 0 15536 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_170
timestamp 1586364061
transform 1 0 16456 0 -1 14688
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17744 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18756 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17560 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_193
timestamp 1586364061
transform 1 0 18572 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_197
timestamp 1586364061
transform 1 0 18940 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  mux_right_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19308 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20504 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_204
timestamp 1586364061
transform 1 0 19584 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_212
timestamp 1586364061
transform 1 0 20320 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20596 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21700 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 24276 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 22804 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_251
timestamp 1586364061
transform 1 0 23908 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26576 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26116 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_259
timestamp 1586364061
transform 1 0 24644 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_271
timestamp 1586364061
transform 1 0 25748 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26208 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 816 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1092 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2196 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3300 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4404 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5508 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6244 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6428 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6520 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7624 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 8728 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_98
timestamp 1586364061
transform 1 0 9832 0 1 14688
box -38 -48 774 592
use scs8hd_buf_2  _21_
timestamp 1586364061
transform 1 0 10660 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__21__A
timestamp 1586364061
transform 1 0 11212 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_106
timestamp 1586364061
transform 1 0 10568 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_111
timestamp 1586364061
transform 1 0 11028 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_115
timestamp 1586364061
transform 1 0 11396 0 1 14688
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12040 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 11948 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12132 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13236 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14340 0 1 14688
box -38 -48 1142 592
use scs8hd_buf_1  mux_right_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16088 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16548 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_159
timestamp 1586364061
transform 1 0 15444 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_165
timestamp 1586364061
transform 1 0 15996 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_169
timestamp 1586364061
transform 1 0 16364 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_173
timestamp 1586364061
transform 1 0 16732 0 1 14688
box -38 -48 774 592
use scs8hd_buf_2  _22_
timestamp 1586364061
transform 1 0 17744 0 1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17652 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__22__A
timestamp 1586364061
transform 1 0 18296 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_181
timestamp 1586364061
transform 1 0 17468 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_188
timestamp 1586364061
transform 1 0 18112 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_192
timestamp 1586364061
transform 1 0 18480 0 1 14688
box -38 -48 774 592
use scs8hd_buf_2  _20_
timestamp 1586364061
transform 1 0 19216 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__20__A
timestamp 1586364061
transform 1 0 19768 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_204
timestamp 1586364061
transform 1 0 19584 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 19952 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21056 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22160 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23264 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23356 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24460 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26576 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25564 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 816 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2196 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3668 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3300 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 3760 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 4864 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 5968 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7072 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9280 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8176 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9372 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10476 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11580 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12684 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 14892 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 13788 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 14984 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16088 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17192 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18296 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20504 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19400 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20596 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21700 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 22804 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 23908 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26576 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26116 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25012 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26208 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 816 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1092 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2196 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3300 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4404 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5508 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6244 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6428 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6520 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7624 0 1 15776
box -38 -48 1142 592
use scs8hd_buf_2  _19_
timestamp 1586364061
transform 1 0 9280 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__18__A
timestamp 1586364061
transform 1 0 9832 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__19__A
timestamp 1586364061
transform 1 0 9096 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_86
timestamp 1586364061
transform 1 0 8728 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9648 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_100
timestamp 1586364061
transform 1 0 10016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_112
timestamp 1586364061
transform 1 0 11120 0 1 15776
box -38 -48 774 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 13420 0 1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12040 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_120
timestamp 1586364061
transform 1 0 11856 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12132 0 1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_25_135
timestamp 1586364061
transform 1 0 13236 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 13972 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_141
timestamp 1586364061
transform 1 0 13788 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_145
timestamp 1586364061
transform 1 0 14156 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_157
timestamp 1586364061
transform 1 0 15260 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_169
timestamp 1586364061
transform 1 0 16364 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17652 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_181
timestamp 1586364061
transform 1 0 17468 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 17744 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 18848 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 19952 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21056 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22160 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23264 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23356 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24460 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26576 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25564 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 816 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 816 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1092 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2196 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3668 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3300 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 3760 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3300 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4404 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 4864 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 5968 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5508 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6244 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _17_
timestamp 1586364061
transform 1 0 7900 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6428 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__16__A
timestamp 1586364061
transform 1 0 7256 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7072 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_62
timestamp 1586364061
transform 1 0 6520 0 1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_72
timestamp 1586364061
transform 1 0 7440 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_76
timestamp 1586364061
transform 1 0 7808 0 1 16864
box -38 -48 130 592
use scs8hd_buf_2  _18_
timestamp 1586364061
transform 1 0 9372 0 -1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9280 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__17__A
timestamp 1586364061
transform 1 0 8452 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8176 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_97
timestamp 1586364061
transform 1 0 9740 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_81
timestamp 1586364061
transform 1 0 8268 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_85
timestamp 1586364061
transform 1 0 8636 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_97
timestamp 1586364061
transform 1 0 9740 0 1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 10476 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_109
timestamp 1586364061
transform 1 0 10844 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_107
timestamp 1586364061
transform 1 0 10660 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_119
timestamp 1586364061
transform 1 0 11764 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12040 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_121
timestamp 1586364061
transform 1 0 11948 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_133
timestamp 1586364061
transform 1 0 13052 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12132 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13236 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 14892 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_145
timestamp 1586364061
transform 1 0 14156 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 14984 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14340 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16088 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17192 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15444 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16548 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17652 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18296 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 17744 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 18848 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20504 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19400 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20596 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 19952 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21700 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21056 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22160 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23264 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 22804 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 23908 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23356 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24460 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26576 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26576 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26116 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25012 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26208 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25564 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 816 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2196 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3668 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3300 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 3760 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 4864 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 5968 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _16_
timestamp 1586364061
transform 1 0 7256 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_68
timestamp 1586364061
transform 1 0 7072 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_74
timestamp 1586364061
transform 1 0 7624 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9280 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_86
timestamp 1586364061
transform 1 0 8728 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9372 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 10476 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_109
timestamp 1586364061
transform 1 0 10844 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_121
timestamp 1586364061
transform 1 0 11948 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_133
timestamp 1586364061
transform 1 0 13052 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 14892 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_145
timestamp 1586364061
transform 1 0 14156 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 14984 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16088 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17192 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18296 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20504 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19400 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20596 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21700 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 22804 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 23908 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26576 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26116 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25012 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26208 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 816 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1092 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2196 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3300 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4404 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5508 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6244 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6428 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 6704 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6520 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_66
timestamp 1586364061
transform 1 0 6888 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_78
timestamp 1586364061
transform 1 0 7992 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_90
timestamp 1586364061
transform 1 0 9096 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_102
timestamp 1586364061
transform 1 0 10200 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_114
timestamp 1586364061
transform 1 0 11304 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12040 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12132 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13236 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14340 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15444 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16548 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17652 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 17744 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 18848 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 19952 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21056 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22160 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23264 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23356 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24460 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26576 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25564 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 816 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2196 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3668 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3300 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 3760 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 4864 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_56
timestamp 1586364061
transform 1 0 5968 0 -1 19040
box -38 -48 590 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 6612 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_62
timestamp 1586364061
transform 1 0 6520 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_67
timestamp 1586364061
transform 1 0 6980 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_79
timestamp 1586364061
transform 1 0 8084 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9280 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9188 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9372 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10476 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11580 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12684 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 14892 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 13788 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 14984 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16088 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17192 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18296 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20504 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19400 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20596 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21700 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 22804 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 23908 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26576 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26116 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25012 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26208 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 816 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1092 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2196 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3300 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_39
timestamp 1586364061
transform 1 0 4404 0 1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 5232 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_47
timestamp 1586364061
transform 1 0 5140 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_50
timestamp 1586364061
transform 1 0 5416 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_58
timestamp 1586364061
transform 1 0 6152 0 1 19040
box -38 -48 314 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 6520 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6428 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 7072 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_66
timestamp 1586364061
transform 1 0 6888 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_70
timestamp 1586364061
transform 1 0 7256 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_82
timestamp 1586364061
transform 1 0 8360 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_94
timestamp 1586364061
transform 1 0 9464 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_106
timestamp 1586364061
transform 1 0 10568 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_31_118
timestamp 1586364061
transform 1 0 11672 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12040 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12132 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13236 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14340 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15444 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16548 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17652 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 17744 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 18848 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 19952 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21056 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22160 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23264 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23356 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24460 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26576 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25564 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 816 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2196 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3668 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3300 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 3760 0 -1 20128
box -38 -48 1142 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 5232 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_32_44
timestamp 1586364061
transform 1 0 4864 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_52
timestamp 1586364061
transform 1 0 5600 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_64
timestamp 1586364061
transform 1 0 6704 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_76
timestamp 1586364061
transform 1 0 7808 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9280 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_88
timestamp 1586364061
transform 1 0 8912 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9372 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10476 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11580 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12684 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 14892 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 13788 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 14984 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16088 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17192 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18296 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20504 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19400 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20596 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21700 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 22804 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 23908 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26576 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26116 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25012 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26208 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 816 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 816 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1092 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2196 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2196 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3668 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3300 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4404 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3300 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 3760 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5508 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6244 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 4864 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 5968 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6428 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6520 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7624 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7072 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9280 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 8728 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 9832 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8176 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9372 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 10936 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10476 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11580 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12040 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12132 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13236 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12684 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 14892 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14340 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 13788 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 14984 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15444 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16548 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16088 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17192 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17652 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 17744 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 18848 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18296 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20504 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 19952 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19400 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20596 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21056 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22160 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21700 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23264 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23356 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24460 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 22804 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 23908 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26576 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26576 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26116 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25564 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25012 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26208 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 816 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1092 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2196 0 1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 3852 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 4404 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 3668 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3300 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_37
timestamp 1586364061
transform 1 0 4220 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_41
timestamp 1586364061
transform 1 0 4588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_53
timestamp 1586364061
transform 1 0 5692 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6428 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6520 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7624 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 8728 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 9832 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 10936 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12040 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12132 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13236 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14340 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15444 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16548 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17652 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 17744 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 18848 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 19952 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21056 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22160 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23264 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23356 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24460 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26576 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25564 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 816 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2196 0 -1 22304
box -38 -48 1142 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 3760 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3668 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3300 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_36
timestamp 1586364061
transform 1 0 4128 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_48
timestamp 1586364061
transform 1 0 5232 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_60
timestamp 1586364061
transform 1 0 6336 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_72
timestamp 1586364061
transform 1 0 7440 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9280 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_84
timestamp 1586364061
transform 1 0 8544 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9372 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10476 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11580 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12684 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 14892 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 13788 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 14984 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16088 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17192 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18296 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20504 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19400 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20596 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21700 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 22804 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 23908 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26576 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26116 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25012 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26208 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 2472 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 816 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 1828 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_3
timestamp 1586364061
transform 1 0 1092 0 1 22304
box -38 -48 774 592
use scs8hd_decap_4  FILLER_37_13
timestamp 1586364061
transform 1 0 2012 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_17
timestamp 1586364061
transform 1 0 2380 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 3024 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_22
timestamp 1586364061
transform 1 0 2840 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_26
timestamp 1586364061
transform 1 0 3208 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_38
timestamp 1586364061
transform 1 0 4312 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_50
timestamp 1586364061
transform 1 0 5416 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_37_58
timestamp 1586364061
transform 1 0 6152 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6428 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6520 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7624 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 8728 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 9832 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 10936 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12040 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12132 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13236 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14340 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15444 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16548 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17652 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 17744 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 18848 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 19952 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21056 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22160 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23264 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23356 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24460 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26576 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25564 0 1 22304
box -38 -48 774 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 1828 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 816 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_3
timestamp 1586364061
transform 1 0 1092 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2196 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3668 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3300 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 3760 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 4864 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 5968 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7072 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9280 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8176 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9372 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10476 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11580 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12684 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 14892 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 13788 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 14984 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16088 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17192 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18296 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20504 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19400 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20596 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21700 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 22804 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 23908 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26576 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26116 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25012 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26208 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 816 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 816 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1092 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2196 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2196 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3668 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4404 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3300 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 3760 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5508 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6244 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 4864 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 5968 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6428 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6520 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7624 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7072 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9280 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 8728 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 9832 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8176 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9372 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 10936 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10476 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11580 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12040 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12132 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13236 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12684 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 14892 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14340 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 13788 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 14984 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15444 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16548 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16088 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17192 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17652 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 17744 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 18848 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18296 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20504 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 19952 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19400 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20596 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21056 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22160 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21700 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23264 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23356 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24460 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 22804 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 23908 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26576 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26576 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26116 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25564 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25012 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26208 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 816 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1092 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2196 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3300 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4404 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5508 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6244 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6428 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6520 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7624 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 8728 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 9832 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 10936 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12040 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12132 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13236 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14340 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15444 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16548 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17652 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 17744 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 18848 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 19952 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21056 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22160 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23264 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23356 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24460 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26576 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25564 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 816 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1092 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2196 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3668 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3300 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 3760 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 4864 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 5968 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6520 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6612 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 7716 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9372 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 8820 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9464 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10568 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11672 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12224 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12316 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13420 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15076 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14524 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15168 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16272 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 17928 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17376 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18020 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 20780 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19124 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20228 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 20872 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 21976 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23632 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23080 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 23724 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26576 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 24828 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 25932 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 6 0 62 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal2 s 13622 27520 13678 28000 6 ccff_head
port 1 nsew default input
rlabel metal2 s 22914 27520 22970 28000 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 27232 280 27712 400 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 27232 7080 27712 7200 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 27232 7760 27712 7880 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 27232 8440 27712 8560 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 27232 9120 27712 9240 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 27232 9800 27712 9920 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 27232 10480 27712 10600 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 27232 11160 27712 11280 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 27232 11840 27712 11960 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 27232 12520 27712 12640 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 27232 13200 27712 13320 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 27232 960 27712 1080 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 27232 1640 27712 1760 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 27232 2320 27712 2440 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 27232 3000 27712 3120 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 27232 3680 27712 3800 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 27232 4360 27712 4480 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 27232 5040 27712 5160 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 27232 5720 27712 5840 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 27232 6400 27712 6520 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 27232 13880 27712 14000 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 27232 20680 27712 20800 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 27232 21360 27712 21480 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 27232 22040 27712 22160 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 27232 22720 27712 22840 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 27232 23400 27712 23520 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 27232 24080 27712 24200 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 27232 24760 27712 24880 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 27232 25440 27712 25560 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 27232 26120 27712 26240 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 27232 26800 27712 26920 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 27232 14560 27712 14680 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 27232 15240 27712 15360 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 27232 15920 27712 16040 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 27232 16600 27712 16720 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 27232 17280 27712 17400 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 27232 17960 27712 18080 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 27232 18640 27712 18760 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 27232 19320 27712 19440 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 27232 20000 27712 20120 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 650 0 706 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 7458 0 7514 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 8102 0 8158 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 8838 0 8894 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 9482 0 9538 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 10218 0 10274 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 10862 0 10918 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 11598 0 11654 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 12242 0 12298 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 12886 0 12942 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 13622 0 13678 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1294 0 1350 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 2030 0 2086 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2674 0 2730 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3410 0 3466 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 4054 0 4110 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4698 0 4754 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 5434 0 5490 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 6078 0 6134 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 6814 0 6870 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 14266 0 14322 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 21074 0 21130 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 21810 0 21866 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 22454 0 22510 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 23190 0 23246 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 23834 0 23890 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 24478 0 24534 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 25214 0 25270 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 25858 0 25914 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 26594 0 26650 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 27238 0 27294 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 15002 0 15058 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 15646 0 15702 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 16290 0 16346 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 17026 0 17082 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 17670 0 17726 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 18406 0 18462 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 19050 0 19106 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 19786 0 19842 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 20430 0 20486 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal2 s 4330 27520 4386 28000 6 prog_clk
port 83 nsew default input
rlabel metal3 s 27232 27480 27712 27600 6 right_top_grid_pin_1_
port 84 nsew default input
rlabel metal4 s 5323 2128 5643 25616 6 vpwr
port 85 nsew default input
rlabel metal4 s 9989 2128 10309 25616 6 vgnd
port 86 nsew default input
<< properties >>
string FIXED_BBOX 1 0 27712 28000
<< end >>
