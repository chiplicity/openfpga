magic
tech EFS8A
magscale 1 2
timestamp 1603801092
<< locali >>
rect 11609 12631 11643 12869
rect 13265 9911 13299 10217
rect 13633 7327 13667 7497
rect 21085 6103 21119 6409
<< viali >>
rect 24581 23817 24615 23851
rect 21729 23749 21763 23783
rect 21244 23613 21278 23647
rect 24188 23613 24222 23647
rect 21315 23477 21349 23511
rect 24259 23477 24293 23511
rect 24581 21641 24615 21675
rect 24188 21437 24222 21471
rect 24259 21301 24293 21335
rect 24188 20961 24222 20995
rect 24259 20757 24293 20791
rect 24213 20553 24247 20587
rect 24188 19873 24222 19907
rect 24259 19669 24293 19703
rect 24172 19261 24206 19295
rect 25041 19261 25075 19295
rect 24259 19193 24293 19227
rect 24673 19125 24707 19159
rect 20508 18785 20542 18819
rect 23176 18785 23210 18819
rect 24188 18785 24222 18819
rect 23247 18649 23281 18683
rect 20579 18581 20613 18615
rect 24259 18581 24293 18615
rect 20441 18377 20475 18411
rect 23477 18241 23511 18275
rect 22164 18173 22198 18207
rect 24188 18173 24222 18207
rect 25168 18173 25202 18207
rect 25593 18173 25627 18207
rect 24581 18105 24615 18139
rect 22235 18037 22269 18071
rect 22649 18037 22683 18071
rect 24259 18037 24293 18071
rect 25041 18037 25075 18071
rect 25271 18037 25305 18071
rect 21545 17833 21579 17867
rect 20533 17697 20567 17731
rect 22649 17697 22683 17731
rect 24188 17697 24222 17731
rect 20717 17493 20751 17527
rect 22281 17493 22315 17527
rect 24259 17493 24293 17527
rect 24213 17289 24247 17323
rect 21269 17153 21303 17187
rect 21637 17153 21671 17187
rect 15749 17085 15783 17119
rect 15933 17085 15967 17119
rect 19521 17085 19555 17119
rect 19705 17085 19739 17119
rect 24724 17085 24758 17119
rect 16577 17017 16611 17051
rect 21361 17017 21395 17051
rect 24811 17017 24845 17051
rect 20073 16949 20107 16983
rect 20625 16949 20659 16983
rect 20993 16949 21027 16983
rect 22281 16949 22315 16983
rect 23661 16949 23695 16983
rect 25133 16949 25167 16983
rect 16025 16745 16059 16779
rect 18417 16745 18451 16779
rect 16669 16677 16703 16711
rect 20809 16677 20843 16711
rect 24903 16677 24937 16711
rect 14921 16609 14955 16643
rect 15565 16609 15599 16643
rect 18233 16609 18267 16643
rect 22557 16609 22591 16643
rect 23788 16609 23822 16643
rect 23891 16609 23925 16643
rect 24816 16609 24850 16643
rect 16577 16541 16611 16575
rect 16853 16541 16887 16575
rect 20717 16541 20751 16575
rect 21361 16541 21395 16575
rect 19521 16405 19555 16439
rect 22465 16405 22499 16439
rect 16577 16201 16611 16235
rect 20441 16201 20475 16235
rect 20717 16201 20751 16235
rect 21453 16201 21487 16235
rect 22557 16201 22591 16235
rect 14553 16065 14587 16099
rect 16945 16065 16979 16099
rect 21637 16065 21671 16099
rect 17405 15997 17439 16031
rect 17681 15997 17715 16031
rect 19521 15997 19555 16031
rect 23017 15997 23051 16031
rect 23293 15997 23327 16031
rect 15657 15929 15691 15963
rect 15749 15929 15783 15963
rect 16301 15929 16335 15963
rect 17589 15929 17623 15963
rect 19429 15929 19463 15963
rect 19883 15929 19917 15963
rect 21729 15929 21763 15963
rect 22281 15929 22315 15963
rect 24213 15929 24247 15963
rect 15105 15861 15139 15895
rect 15473 15861 15507 15895
rect 18693 15861 18727 15895
rect 23477 15861 23511 15895
rect 24765 15861 24799 15895
rect 25317 15861 25351 15895
rect 16209 15657 16243 15691
rect 21637 15657 21671 15691
rect 15651 15589 15685 15623
rect 17221 15589 17255 15623
rect 20803 15589 20837 15623
rect 22281 15589 22315 15623
rect 22373 15589 22407 15623
rect 12897 15521 12931 15555
rect 13044 15521 13078 15555
rect 19061 15521 19095 15555
rect 19245 15521 19279 15555
rect 21361 15521 21395 15555
rect 24397 15521 24431 15555
rect 13265 15453 13299 15487
rect 15289 15453 15323 15487
rect 17129 15453 17163 15487
rect 17405 15453 17439 15487
rect 19521 15453 19555 15487
rect 20441 15453 20475 15487
rect 22557 15453 22591 15487
rect 24489 15453 24523 15487
rect 20257 15385 20291 15419
rect 13173 15317 13207 15351
rect 13541 15317 13575 15351
rect 13909 15317 13943 15351
rect 15013 15317 15047 15351
rect 12253 15113 12287 15147
rect 12989 15113 13023 15147
rect 15657 15113 15691 15147
rect 16301 15113 16335 15147
rect 17037 15113 17071 15147
rect 20073 15113 20107 15147
rect 20533 15113 20567 15147
rect 22281 15113 22315 15147
rect 25225 15113 25259 15147
rect 12621 15045 12655 15079
rect 13909 14977 13943 15011
rect 14737 14977 14771 15011
rect 19245 14977 19279 15011
rect 20809 14977 20843 15011
rect 22557 14977 22591 15011
rect 13449 14909 13483 14943
rect 13725 14909 13759 14943
rect 18601 14909 18635 14943
rect 18969 14909 19003 14943
rect 23017 14909 23051 14943
rect 23293 14909 23327 14943
rect 24832 14909 24866 14943
rect 14185 14841 14219 14875
rect 14645 14841 14679 14875
rect 15099 14841 15133 14875
rect 20901 14841 20935 14875
rect 21453 14841 21487 14875
rect 23201 14841 23235 14875
rect 24305 14841 24339 14875
rect 15933 14773 15967 14807
rect 16485 14773 16519 14807
rect 17957 14773 17991 14807
rect 18325 14773 18359 14807
rect 19521 14773 19555 14807
rect 21729 14773 21763 14807
rect 24903 14773 24937 14807
rect 12989 14569 13023 14603
rect 16485 14569 16519 14603
rect 17865 14569 17899 14603
rect 18601 14569 18635 14603
rect 20257 14569 20291 14603
rect 21361 14569 21395 14603
rect 15013 14501 15047 14535
rect 15565 14501 15599 14535
rect 17497 14501 17531 14535
rect 20803 14501 20837 14535
rect 21637 14501 21671 14535
rect 22373 14501 22407 14535
rect 9677 14433 9711 14467
rect 9861 14433 9895 14467
rect 11793 14433 11827 14467
rect 13449 14433 13483 14467
rect 13725 14433 13759 14467
rect 16669 14433 16703 14467
rect 16853 14433 16887 14467
rect 19061 14433 19095 14467
rect 19337 14433 19371 14467
rect 23845 14433 23879 14467
rect 13909 14365 13943 14399
rect 14921 14365 14955 14399
rect 19521 14365 19555 14399
rect 20441 14365 20475 14399
rect 22281 14365 22315 14399
rect 22925 14365 22959 14399
rect 23753 14365 23787 14399
rect 9953 14229 9987 14263
rect 11977 14229 12011 14263
rect 19797 14229 19831 14263
rect 23201 14229 23235 14263
rect 8941 14025 8975 14059
rect 10137 14025 10171 14059
rect 14093 14025 14127 14059
rect 15657 14025 15691 14059
rect 16393 14025 16427 14059
rect 17405 14025 17439 14059
rect 18877 14025 18911 14059
rect 20257 14025 20291 14059
rect 20625 14025 20659 14059
rect 20901 14025 20935 14059
rect 21453 14025 21487 14059
rect 22649 14025 22683 14059
rect 24213 14025 24247 14059
rect 11057 13957 11091 13991
rect 12437 13957 12471 13991
rect 14553 13957 14587 13991
rect 17037 13957 17071 13991
rect 19245 13957 19279 13991
rect 22189 13957 22223 13991
rect 24949 13957 24983 13991
rect 9861 13889 9895 13923
rect 10505 13889 10539 13923
rect 12253 13889 12287 13923
rect 13817 13889 13851 13923
rect 17957 13889 17991 13923
rect 19337 13889 19371 13923
rect 21637 13889 21671 13923
rect 9217 13821 9251 13855
rect 10873 13821 10907 13855
rect 11333 13821 11367 13855
rect 12529 13821 12563 13855
rect 13081 13821 13115 13855
rect 13449 13821 13483 13855
rect 14829 13821 14863 13855
rect 15105 13821 15139 13855
rect 23017 13821 23051 13855
rect 23201 13821 23235 13855
rect 23753 13821 23787 13855
rect 24765 13821 24799 13855
rect 25317 13821 25351 13855
rect 15381 13753 15415 13787
rect 17681 13753 17715 13787
rect 17773 13753 17807 13787
rect 19699 13753 19733 13787
rect 21729 13753 21763 13787
rect 11701 13685 11735 13719
rect 16485 13685 16519 13719
rect 23293 13685 23327 13719
rect 12437 13481 12471 13515
rect 15013 13481 15047 13515
rect 15473 13481 15507 13515
rect 16485 13481 16519 13515
rect 19153 13481 19187 13515
rect 22281 13481 22315 13515
rect 23477 13481 23511 13515
rect 12805 13413 12839 13447
rect 15927 13413 15961 13447
rect 17221 13413 17255 13447
rect 17405 13413 17439 13447
rect 17497 13413 17531 13447
rect 20625 13413 20659 13447
rect 21177 13413 21211 13447
rect 22557 13413 22591 13447
rect 9401 13345 9435 13379
rect 9953 13345 9987 13379
rect 11885 13345 11919 13379
rect 13081 13345 13115 13379
rect 15565 13345 15599 13379
rect 18877 13345 18911 13379
rect 19061 13345 19095 13379
rect 24213 13345 24247 13379
rect 14185 13277 14219 13311
rect 20533 13277 20567 13311
rect 22465 13277 22499 13311
rect 23109 13277 23143 13311
rect 23937 13277 23971 13311
rect 17957 13209 17991 13243
rect 18785 13209 18819 13243
rect 9493 13141 9527 13175
rect 10505 13141 10539 13175
rect 10781 13141 10815 13175
rect 11701 13141 11735 13175
rect 13817 13141 13851 13175
rect 19705 13141 19739 13175
rect 21453 13141 21487 13175
rect 9217 12937 9251 12971
rect 10137 12937 10171 12971
rect 10597 12937 10631 12971
rect 13633 12937 13667 12971
rect 14093 12937 14127 12971
rect 14277 12937 14311 12971
rect 16945 12937 16979 12971
rect 18969 12937 19003 12971
rect 20441 12937 20475 12971
rect 22465 12937 22499 12971
rect 24213 12937 24247 12971
rect 9493 12869 9527 12903
rect 9769 12869 9803 12903
rect 10459 12869 10493 12903
rect 11333 12869 11367 12903
rect 11609 12869 11643 12903
rect 17313 12869 17347 12903
rect 20993 12869 21027 12903
rect 10689 12801 10723 12835
rect 9309 12733 9343 12767
rect 10321 12665 10355 12699
rect 13964 12801 13998 12835
rect 14185 12801 14219 12835
rect 15749 12801 15783 12835
rect 17681 12801 17715 12835
rect 17957 12801 17991 12835
rect 19797 12801 19831 12835
rect 21085 12801 21119 12835
rect 23569 12801 23603 12835
rect 12161 12733 12195 12767
rect 13817 12733 13851 12767
rect 19153 12733 19187 12767
rect 19705 12733 19739 12767
rect 20864 12733 20898 12767
rect 21453 12733 21487 12767
rect 24765 12733 24799 12767
rect 25317 12733 25351 12767
rect 14829 12665 14863 12699
rect 15289 12665 15323 12699
rect 15657 12665 15691 12699
rect 16111 12665 16145 12699
rect 17773 12665 17807 12699
rect 20717 12665 20751 12699
rect 23293 12665 23327 12699
rect 23385 12665 23419 12699
rect 10965 12597 10999 12631
rect 11609 12597 11643 12631
rect 11701 12597 11735 12631
rect 12253 12597 12287 12631
rect 13081 12597 13115 12631
rect 16669 12597 16703 12631
rect 21729 12597 21763 12631
rect 23017 12597 23051 12631
rect 24949 12597 24983 12631
rect 10597 12393 10631 12427
rect 13081 12393 13115 12427
rect 13817 12393 13851 12427
rect 14185 12393 14219 12427
rect 16117 12393 16151 12427
rect 17313 12393 17347 12427
rect 19705 12393 19739 12427
rect 21085 12393 21119 12427
rect 22281 12393 22315 12427
rect 24995 12393 25029 12427
rect 12529 12325 12563 12359
rect 16485 12325 16519 12359
rect 17037 12325 17071 12359
rect 19429 12325 19463 12359
rect 21682 12325 21716 12359
rect 23477 12325 23511 12359
rect 8113 12257 8147 12291
rect 10045 12257 10079 12291
rect 11057 12257 11091 12291
rect 13173 12257 13207 12291
rect 18325 12257 18359 12291
rect 19061 12257 19095 12291
rect 21361 12257 21395 12291
rect 24892 12257 24926 12291
rect 10965 12189 10999 12223
rect 11425 12189 11459 12223
rect 13541 12189 13575 12223
rect 15289 12189 15323 12223
rect 16393 12189 16427 12223
rect 18693 12189 18727 12223
rect 23385 12189 23419 12223
rect 23661 12189 23695 12223
rect 14553 12121 14587 12155
rect 18463 12121 18497 12155
rect 20717 12121 20751 12155
rect 8297 12053 8331 12087
rect 9953 12053 9987 12087
rect 10229 12053 10263 12087
rect 11222 12053 11256 12087
rect 11333 12053 11367 12087
rect 11517 12053 11551 12087
rect 12161 12053 12195 12087
rect 13338 12053 13372 12087
rect 13449 12053 13483 12087
rect 15841 12053 15875 12087
rect 17773 12053 17807 12087
rect 18233 12053 18267 12087
rect 18601 12053 18635 12087
rect 20257 12053 20291 12087
rect 22557 12053 22591 12087
rect 7745 11849 7779 11883
rect 8665 11849 8699 11883
rect 9401 11849 9435 11883
rect 10137 11849 10171 11883
rect 11241 11849 11275 11883
rect 13265 11849 13299 11883
rect 14277 11849 14311 11883
rect 15197 11849 15231 11883
rect 16485 11849 16519 11883
rect 17313 11849 17347 11883
rect 18858 11849 18892 11883
rect 19797 11849 19831 11883
rect 20257 11849 20291 11883
rect 23017 11849 23051 11883
rect 24765 11849 24799 11883
rect 9125 11781 9159 11815
rect 12253 11781 12287 11815
rect 13725 11781 13759 11815
rect 13955 11781 13989 11815
rect 14093 11781 14127 11815
rect 18969 11781 19003 11815
rect 24305 11781 24339 11815
rect 12345 11713 12379 11747
rect 14185 11713 14219 11747
rect 18141 11713 18175 11747
rect 19061 11713 19095 11747
rect 20809 11713 20843 11747
rect 21177 11713 21211 11747
rect 23385 11713 23419 11747
rect 23661 11713 23695 11747
rect 7193 11645 7227 11679
rect 8205 11645 8239 11679
rect 9217 11645 9251 11679
rect 10229 11645 10263 11679
rect 10781 11645 10815 11679
rect 12124 11645 12158 11679
rect 15381 11645 15415 11679
rect 15841 11645 15875 11679
rect 17716 11645 17750 11679
rect 17819 11645 17853 11679
rect 20416 11645 20450 11679
rect 21361 11645 21395 11679
rect 24857 11645 24891 11679
rect 25409 11645 25443 11679
rect 9677 11577 9711 11611
rect 11977 11577 12011 11611
rect 13817 11577 13851 11611
rect 14921 11577 14955 11611
rect 18693 11577 18727 11611
rect 19429 11577 19463 11611
rect 21682 11577 21716 11611
rect 23477 11577 23511 11611
rect 7377 11509 7411 11543
rect 8389 11509 8423 11543
rect 10505 11509 10539 11543
rect 11701 11509 11735 11543
rect 12621 11509 12655 11543
rect 15473 11509 15507 11543
rect 16761 11509 16795 11543
rect 18509 11509 18543 11543
rect 20487 11509 20521 11543
rect 22281 11509 22315 11543
rect 22649 11509 22683 11543
rect 25041 11509 25075 11543
rect 10045 11305 10079 11339
rect 10965 11305 10999 11339
rect 12161 11305 12195 11339
rect 12437 11305 12471 11339
rect 13633 11305 13667 11339
rect 14001 11305 14035 11339
rect 14461 11305 14495 11339
rect 16485 11305 16519 11339
rect 22281 11305 22315 11339
rect 23477 11305 23511 11339
rect 24121 11305 24155 11339
rect 12621 11237 12655 11271
rect 14829 11237 14863 11271
rect 16301 11237 16335 11271
rect 19705 11237 19739 11271
rect 21913 11237 21947 11271
rect 22649 11237 22683 11271
rect 8113 11169 8147 11203
rect 9861 11169 9895 11203
rect 11057 11169 11091 11203
rect 13265 11169 13299 11203
rect 16669 11169 16703 11203
rect 16853 11169 16887 11203
rect 18141 11169 18175 11203
rect 18693 11169 18727 11203
rect 20441 11169 20475 11203
rect 20901 11169 20935 11203
rect 21453 11169 21487 11203
rect 24305 11169 24339 11203
rect 24489 11169 24523 11203
rect 10597 11101 10631 11135
rect 11425 11101 11459 11135
rect 11517 11101 11551 11135
rect 15197 11101 15231 11135
rect 17405 11101 17439 11135
rect 19061 11101 19095 11135
rect 20993 11101 21027 11135
rect 22557 11101 22591 11135
rect 23017 11101 23051 11135
rect 8297 11033 8331 11067
rect 9769 11033 9803 11067
rect 11222 11033 11256 11067
rect 15105 11033 15139 11067
rect 17865 11033 17899 11067
rect 19153 11033 19187 11067
rect 11333 10965 11367 10999
rect 14967 10965 15001 10999
rect 15289 10965 15323 10999
rect 18509 10965 18543 10999
rect 18831 10965 18865 10999
rect 18969 10965 19003 10999
rect 8113 10761 8147 10795
rect 9861 10761 9895 10795
rect 11333 10761 11367 10795
rect 11701 10761 11735 10795
rect 13081 10761 13115 10795
rect 13449 10761 13483 10795
rect 13817 10761 13851 10795
rect 14166 10761 14200 10795
rect 16577 10761 16611 10795
rect 19291 10761 19325 10795
rect 20165 10761 20199 10795
rect 22281 10761 22315 10795
rect 24765 10761 24799 10795
rect 8481 10693 8515 10727
rect 9217 10693 9251 10727
rect 14277 10693 14311 10727
rect 19429 10693 19463 10727
rect 22925 10693 22959 10727
rect 24397 10693 24431 10727
rect 12069 10625 12103 10659
rect 14369 10625 14403 10659
rect 15013 10625 15047 10659
rect 18693 10625 18727 10659
rect 19521 10625 19555 10659
rect 20625 10625 20659 10659
rect 21269 10625 21303 10659
rect 8297 10557 8331 10591
rect 9309 10557 9343 10591
rect 10321 10557 10355 10591
rect 10781 10557 10815 10591
rect 14001 10557 14035 10591
rect 15657 10557 15691 10591
rect 17589 10557 17623 10591
rect 18049 10557 18083 10591
rect 20717 10557 20751 10591
rect 21177 10557 21211 10591
rect 21729 10557 21763 10591
rect 23201 10557 23235 10591
rect 24949 10557 24983 10591
rect 25501 10557 25535 10591
rect 8849 10489 8883 10523
rect 11057 10489 11091 10523
rect 12161 10489 12195 10523
rect 12713 10489 12747 10523
rect 15565 10489 15599 10523
rect 17313 10489 17347 10523
rect 18325 10489 18359 10523
rect 19153 10489 19187 10523
rect 19889 10489 19923 10523
rect 22557 10489 22591 10523
rect 23522 10489 23556 10523
rect 9493 10421 9527 10455
rect 14645 10421 14679 10455
rect 15381 10421 15415 10455
rect 16945 10421 16979 10455
rect 24121 10421 24155 10455
rect 25133 10421 25167 10455
rect 9861 10217 9895 10251
rect 11241 10217 11275 10251
rect 11517 10217 11551 10251
rect 13081 10217 13115 10251
rect 13265 10217 13299 10251
rect 14185 10217 14219 10251
rect 14553 10217 14587 10251
rect 16209 10217 16243 10251
rect 17589 10217 17623 10251
rect 19153 10217 19187 10251
rect 19521 10217 19555 10251
rect 19889 10217 19923 10251
rect 20625 10217 20659 10251
rect 21913 10217 21947 10251
rect 22557 10217 22591 10251
rect 10683 10149 10717 10183
rect 12253 10149 12287 10183
rect 9309 10081 9343 10115
rect 10321 10081 10355 10115
rect 12161 10013 12195 10047
rect 12713 9945 12747 9979
rect 16755 10149 16789 10183
rect 21355 10149 21389 10183
rect 24213 10149 24247 10183
rect 13633 10081 13667 10115
rect 14829 10081 14863 10115
rect 15289 10081 15323 10115
rect 16393 10081 16427 10115
rect 18141 10081 18175 10115
rect 18288 10081 18322 10115
rect 20993 10081 21027 10115
rect 23084 10081 23118 10115
rect 15565 10013 15599 10047
rect 18509 10013 18543 10047
rect 24121 10013 24155 10047
rect 24765 10013 24799 10047
rect 13541 9945 13575 9979
rect 9493 9877 9527 9911
rect 10137 9877 10171 9911
rect 11977 9877 12011 9911
rect 13265 9877 13299 9911
rect 13817 9877 13851 9911
rect 15841 9877 15875 9911
rect 17313 9877 17347 9911
rect 17957 9877 17991 9911
rect 18417 9877 18451 9911
rect 18601 9877 18635 9911
rect 23155 9877 23189 9911
rect 9033 9673 9067 9707
rect 14921 9673 14955 9707
rect 15197 9673 15231 9707
rect 17313 9673 17347 9707
rect 18693 9673 18727 9707
rect 18969 9673 19003 9707
rect 19318 9673 19352 9707
rect 20165 9673 20199 9707
rect 11333 9605 11367 9639
rect 11793 9605 11827 9639
rect 12989 9605 13023 9639
rect 16025 9605 16059 9639
rect 20809 9605 20843 9639
rect 21085 9605 21119 9639
rect 22465 9605 22499 9639
rect 10137 9537 10171 9571
rect 11057 9537 11091 9571
rect 15473 9537 15507 9571
rect 17681 9537 17715 9571
rect 19521 9537 19555 9571
rect 21269 9537 21303 9571
rect 22833 9537 22867 9571
rect 25501 9537 25535 9571
rect 9176 9469 9210 9503
rect 9585 9469 9619 9503
rect 13357 9469 13391 9503
rect 13725 9469 13759 9503
rect 13909 9469 13943 9503
rect 14277 9469 14311 9503
rect 19383 9469 19417 9503
rect 22189 9469 22223 9503
rect 24857 9469 24891 9503
rect 9263 9401 9297 9435
rect 10413 9401 10447 9435
rect 10505 9401 10539 9435
rect 12621 9401 12655 9435
rect 15565 9401 15599 9435
rect 17037 9401 17071 9435
rect 17773 9401 17807 9435
rect 18325 9401 18359 9435
rect 19153 9401 19187 9435
rect 21590 9401 21624 9435
rect 24213 9401 24247 9435
rect 24305 9401 24339 9435
rect 25133 9401 25167 9435
rect 11977 9333 12011 9367
rect 14553 9333 14587 9367
rect 16485 9333 16519 9367
rect 19797 9333 19831 9367
rect 23477 9333 23511 9367
rect 24029 9333 24063 9367
rect 10965 9129 10999 9163
rect 12069 9129 12103 9163
rect 12437 9129 12471 9163
rect 12805 9129 12839 9163
rect 14645 9129 14679 9163
rect 16485 9129 16519 9163
rect 18601 9129 18635 9163
rect 19153 9129 19187 9163
rect 19475 9129 19509 9163
rect 24121 9129 24155 9163
rect 11470 9061 11504 9095
rect 13081 9061 13115 9095
rect 16853 9061 16887 9095
rect 17681 9061 17715 9095
rect 19797 9061 19831 9095
rect 21453 9061 21487 9095
rect 22005 9061 22039 9095
rect 22741 9061 22775 9095
rect 22925 9061 22959 9095
rect 23017 9061 23051 9095
rect 24397 9061 24431 9095
rect 10229 8993 10263 9027
rect 10321 8993 10355 9027
rect 10597 8993 10631 9027
rect 11149 8993 11183 9027
rect 14829 8993 14863 9027
rect 15657 8993 15691 9027
rect 19404 8993 19438 9027
rect 24489 8993 24523 9027
rect 12989 8925 13023 8959
rect 13357 8925 13391 8959
rect 15565 8925 15599 8959
rect 17589 8925 17623 8959
rect 17865 8925 17899 8959
rect 21361 8925 21395 8959
rect 23201 8925 23235 8959
rect 15657 8857 15691 8891
rect 17405 8857 17439 8891
rect 13909 8789 13943 8823
rect 20901 8789 20935 8823
rect 9493 8585 9527 8619
rect 11241 8585 11275 8619
rect 13449 8585 13483 8619
rect 15013 8585 15047 8619
rect 16945 8585 16979 8619
rect 19245 8585 19279 8619
rect 20717 8585 20751 8619
rect 21913 8585 21947 8619
rect 22649 8585 22683 8619
rect 23017 8585 23051 8619
rect 24397 8585 24431 8619
rect 24949 8585 24983 8619
rect 9769 8517 9803 8551
rect 11793 8517 11827 8551
rect 14277 8517 14311 8551
rect 10505 8449 10539 8483
rect 12713 8449 12747 8483
rect 12989 8449 13023 8483
rect 15473 8449 15507 8483
rect 17405 8449 17439 8483
rect 17589 8449 17623 8483
rect 23569 8449 23603 8483
rect 9953 8381 9987 8415
rect 10413 8381 10447 8415
rect 12069 8381 12103 8415
rect 13541 8381 13575 8415
rect 14001 8381 14035 8415
rect 14369 8381 14403 8415
rect 16393 8381 16427 8415
rect 18233 8381 18267 8415
rect 19337 8381 19371 8415
rect 19797 8381 19831 8415
rect 20901 8381 20935 8415
rect 21361 8381 21395 8415
rect 24765 8381 24799 8415
rect 25317 8381 25351 8415
rect 8941 8313 8975 8347
rect 15381 8313 15415 8347
rect 15835 8313 15869 8347
rect 18877 8313 18911 8347
rect 20073 8313 20107 8347
rect 23293 8313 23327 8347
rect 23385 8313 23419 8347
rect 21177 8245 21211 8279
rect 10045 8041 10079 8075
rect 10597 8041 10631 8075
rect 11333 8041 11367 8075
rect 12069 8041 12103 8075
rect 12989 8041 13023 8075
rect 14185 8041 14219 8075
rect 14645 8041 14679 8075
rect 15749 8041 15783 8075
rect 16393 8041 16427 8075
rect 17773 8041 17807 8075
rect 18417 8041 18451 8075
rect 19797 8041 19831 8075
rect 21637 8041 21671 8075
rect 23293 8041 23327 8075
rect 15191 7973 15225 8007
rect 17174 7973 17208 8007
rect 20803 7973 20837 8007
rect 22373 7973 22407 8007
rect 8205 7905 8239 7939
rect 10321 7905 10355 7939
rect 10873 7905 10907 7939
rect 12228 7905 12262 7939
rect 13265 7905 13299 7939
rect 14829 7905 14863 7939
rect 16853 7905 16887 7939
rect 18969 7905 19003 7939
rect 19245 7905 19279 7939
rect 23845 7905 23879 7939
rect 8297 7837 8331 7871
rect 9309 7837 9343 7871
rect 13909 7837 13943 7871
rect 16025 7837 16059 7871
rect 19521 7837 19555 7871
rect 20441 7837 20475 7871
rect 22281 7837 22315 7871
rect 22557 7837 22591 7871
rect 23569 7837 23603 7871
rect 23753 7837 23787 7871
rect 12299 7769 12333 7803
rect 18141 7701 18175 7735
rect 21361 7701 21395 7735
rect 7653 7497 7687 7531
rect 10229 7497 10263 7531
rect 11425 7497 11459 7531
rect 13081 7497 13115 7531
rect 13633 7497 13667 7531
rect 13725 7497 13759 7531
rect 15381 7497 15415 7531
rect 15749 7497 15783 7531
rect 17221 7497 17255 7531
rect 19061 7497 19095 7531
rect 19521 7497 19555 7531
rect 20717 7497 20751 7531
rect 20993 7497 21027 7531
rect 22465 7497 22499 7531
rect 7745 7361 7779 7395
rect 8665 7361 8699 7395
rect 9861 7361 9895 7395
rect 13449 7361 13483 7395
rect 14645 7429 14679 7463
rect 17865 7361 17899 7395
rect 18417 7361 18451 7395
rect 20165 7361 20199 7395
rect 21177 7361 21211 7395
rect 23293 7361 23327 7395
rect 23569 7361 23603 7395
rect 9033 7293 9067 7327
rect 9309 7293 9343 7327
rect 10321 7293 10355 7327
rect 10873 7293 10907 7327
rect 12253 7293 12287 7327
rect 12529 7293 12563 7327
rect 13633 7293 13667 7327
rect 13909 7293 13943 7327
rect 14369 7293 14403 7327
rect 14737 7293 14771 7327
rect 15933 7293 15967 7327
rect 19613 7293 19647 7327
rect 20073 7293 20107 7327
rect 22097 7293 22131 7327
rect 24765 7293 24799 7327
rect 25317 7293 25351 7327
rect 9493 7225 9527 7259
rect 11057 7225 11091 7259
rect 16945 7225 16979 7259
rect 18141 7225 18175 7259
rect 18233 7225 18267 7259
rect 21498 7225 21532 7259
rect 23017 7225 23051 7259
rect 23385 7225 23419 7259
rect 11701 7157 11735 7191
rect 12069 7157 12103 7191
rect 16117 7157 16151 7191
rect 24213 7157 24247 7191
rect 24949 7157 24983 7191
rect 12621 6953 12655 6987
rect 14277 6953 14311 6987
rect 15289 6953 15323 6987
rect 19061 6953 19095 6987
rect 19705 6953 19739 6987
rect 20901 6953 20935 6987
rect 21269 6953 21303 6987
rect 22465 6953 22499 6987
rect 10223 6885 10257 6919
rect 13357 6885 13391 6919
rect 18141 6885 18175 6919
rect 21637 6885 21671 6919
rect 22189 6885 22223 6919
rect 23385 6885 23419 6919
rect 8113 6817 8147 6851
rect 8849 6817 8883 6851
rect 9861 6817 9895 6851
rect 11057 6817 11091 6851
rect 11701 6817 11735 6851
rect 12161 6817 12195 6851
rect 14896 6817 14930 6851
rect 16393 6817 16427 6851
rect 20476 6817 20510 6851
rect 20579 6817 20613 6851
rect 24765 6817 24799 6851
rect 12345 6749 12379 6783
rect 13265 6749 13299 6783
rect 13909 6749 13943 6783
rect 16577 6749 16611 6783
rect 18049 6749 18083 6783
rect 18417 6749 18451 6783
rect 21545 6749 21579 6783
rect 23293 6749 23327 6783
rect 23569 6749 23603 6783
rect 10781 6613 10815 6647
rect 14967 6613 15001 6647
rect 15749 6613 15783 6647
rect 24949 6613 24983 6647
rect 6503 6409 6537 6443
rect 9677 6409 9711 6443
rect 10045 6409 10079 6443
rect 11701 6409 11735 6443
rect 13541 6409 13575 6443
rect 18601 6409 18635 6443
rect 19613 6409 19647 6443
rect 21085 6409 21119 6443
rect 21177 6409 21211 6443
rect 23017 6409 23051 6443
rect 24581 6409 24615 6443
rect 15105 6341 15139 6375
rect 8113 6273 8147 6307
rect 11977 6273 12011 6307
rect 13265 6273 13299 6307
rect 14185 6273 14219 6307
rect 16025 6273 16059 6307
rect 16301 6273 16335 6307
rect 17681 6273 17715 6307
rect 18141 6273 18175 6307
rect 6411 6205 6445 6239
rect 6825 6205 6859 6239
rect 7612 6205 7646 6239
rect 8481 6205 8515 6239
rect 9217 6205 9251 6239
rect 10137 6205 10171 6239
rect 19797 6205 19831 6239
rect 20257 6205 20291 6239
rect 20901 6205 20935 6239
rect 7699 6137 7733 6171
rect 10458 6137 10492 6171
rect 12339 6137 12373 6171
rect 14093 6137 14127 6171
rect 14547 6137 14581 6171
rect 16117 6137 16151 6171
rect 17773 6137 17807 6171
rect 20533 6137 20567 6171
rect 22649 6273 22683 6307
rect 21361 6205 21395 6239
rect 23201 6205 23235 6239
rect 23661 6205 23695 6239
rect 24765 6205 24799 6239
rect 25317 6205 25351 6239
rect 21723 6137 21757 6171
rect 8849 6069 8883 6103
rect 11057 6069 11091 6103
rect 11425 6069 11459 6103
rect 12897 6069 12931 6103
rect 15473 6069 15507 6103
rect 15841 6069 15875 6103
rect 17405 6069 17439 6103
rect 21085 6069 21119 6103
rect 22281 6069 22315 6103
rect 23293 6069 23327 6103
rect 24949 6069 24983 6103
rect 10505 5865 10539 5899
rect 10873 5865 10907 5899
rect 12621 5865 12655 5899
rect 14277 5865 14311 5899
rect 16025 5865 16059 5899
rect 17681 5865 17715 5899
rect 18049 5865 18083 5899
rect 19245 5865 19279 5899
rect 20533 5865 20567 5899
rect 21545 5865 21579 5899
rect 9677 5797 9711 5831
rect 11419 5797 11453 5831
rect 12253 5797 12287 5831
rect 13081 5797 13115 5831
rect 15191 5797 15225 5831
rect 16761 5797 16795 5831
rect 19889 5797 19923 5831
rect 20257 5797 20291 5831
rect 21821 5797 21855 5831
rect 22326 5797 22360 5831
rect 23201 5797 23235 5831
rect 23937 5797 23971 5831
rect 6584 5729 6618 5763
rect 8205 5729 8239 5763
rect 11057 5729 11091 5763
rect 14829 5729 14863 5763
rect 18417 5729 18451 5763
rect 18601 5729 18635 5763
rect 20441 5729 20475 5763
rect 20901 5729 20935 5763
rect 23569 5729 23603 5763
rect 8297 5661 8331 5695
rect 9585 5661 9619 5695
rect 9861 5661 9895 5695
rect 12989 5661 13023 5695
rect 13357 5661 13391 5695
rect 16669 5661 16703 5695
rect 16945 5661 16979 5695
rect 18693 5661 18727 5695
rect 22005 5661 22039 5695
rect 23845 5661 23879 5695
rect 6687 5593 6721 5627
rect 24397 5593 24431 5627
rect 11977 5525 12011 5559
rect 15749 5525 15783 5559
rect 22925 5525 22959 5559
rect 6181 5321 6215 5355
rect 7377 5321 7411 5355
rect 8849 5321 8883 5355
rect 10045 5321 10079 5355
rect 11701 5321 11735 5355
rect 14185 5321 14219 5355
rect 16945 5321 16979 5355
rect 17865 5321 17899 5355
rect 20073 5321 20107 5355
rect 20533 5321 20567 5355
rect 24489 5321 24523 5355
rect 10413 5253 10447 5287
rect 16577 5253 16611 5287
rect 19797 5253 19831 5287
rect 24857 5253 24891 5287
rect 6457 5185 6491 5219
rect 9769 5185 9803 5219
rect 12529 5185 12563 5219
rect 15749 5185 15783 5219
rect 17313 5185 17347 5219
rect 18325 5185 18359 5219
rect 20625 5185 20659 5219
rect 22373 5185 22407 5219
rect 23569 5185 23603 5219
rect 7009 5117 7043 5151
rect 8113 5117 8147 5151
rect 10924 5117 10958 5151
rect 14553 5117 14587 5151
rect 15289 5117 15323 5151
rect 16393 5117 16427 5151
rect 19245 5117 19279 5151
rect 25041 5117 25075 5151
rect 25593 5117 25627 5151
rect 8205 5049 8239 5083
rect 9125 5049 9159 5083
rect 9217 5049 9251 5083
rect 11011 5049 11045 5083
rect 12437 5049 12471 5083
rect 12891 5049 12925 5083
rect 14645 5049 14679 5083
rect 18233 5049 18267 5083
rect 18687 5049 18721 5083
rect 20946 5049 20980 5083
rect 22005 5049 22039 5083
rect 23661 5049 23695 5083
rect 24213 5049 24247 5083
rect 8481 4981 8515 5015
rect 11425 4981 11459 5015
rect 13449 4981 13483 5015
rect 13725 4981 13759 5015
rect 16209 4981 16243 5015
rect 21545 4981 21579 5015
rect 23017 4981 23051 5015
rect 25225 4981 25259 5015
rect 5675 4777 5709 4811
rect 10321 4777 10355 4811
rect 11793 4777 11827 4811
rect 12529 4777 12563 4811
rect 12989 4777 13023 4811
rect 18233 4777 18267 4811
rect 21361 4777 21395 4811
rect 22097 4777 22131 4811
rect 23385 4777 23419 4811
rect 10867 4709 10901 4743
rect 13357 4709 13391 4743
rect 16571 4709 16605 4743
rect 18963 4709 18997 4743
rect 20803 4709 20837 4743
rect 23661 4709 23695 4743
rect 4592 4641 4626 4675
rect 5604 4641 5638 4675
rect 8205 4641 8239 4675
rect 9493 4641 9527 4675
rect 10505 4641 10539 4675
rect 15105 4641 15139 4675
rect 16209 4641 16243 4675
rect 18601 4641 18635 4675
rect 20441 4641 20475 4675
rect 22189 4641 22223 4675
rect 22741 4641 22775 4675
rect 6549 4573 6583 4607
rect 8297 4573 8331 4607
rect 13265 4573 13299 4607
rect 13909 4573 13943 4607
rect 23569 4573 23603 4607
rect 24213 4573 24247 4607
rect 4663 4505 4697 4539
rect 22373 4505 22407 4539
rect 11425 4437 11459 4471
rect 15289 4437 15323 4471
rect 17129 4437 17163 4471
rect 17589 4437 17623 4471
rect 19521 4437 19555 4471
rect 11333 4233 11367 4267
rect 13449 4233 13483 4267
rect 16761 4233 16795 4267
rect 18601 4233 18635 4267
rect 20901 4233 20935 4267
rect 21361 4233 21395 4267
rect 24213 4233 24247 4267
rect 20625 4165 20659 4199
rect 7653 4097 7687 4131
rect 10413 4097 10447 4131
rect 12437 4097 12471 4131
rect 13081 4097 13115 4131
rect 14001 4097 14035 4131
rect 14277 4097 14311 4131
rect 15565 4097 15599 4131
rect 17957 4097 17991 4131
rect 18969 4097 19003 4131
rect 19889 4097 19923 4131
rect 21545 4097 21579 4131
rect 22557 4097 22591 4131
rect 23017 4097 23051 4131
rect 23569 4097 23603 4131
rect 3304 4029 3338 4063
rect 4316 4029 4350 4063
rect 5328 4029 5362 4063
rect 6089 4029 6123 4063
rect 7745 4029 7779 4063
rect 8665 4029 8699 4063
rect 9125 4029 9159 4063
rect 15749 4029 15783 4063
rect 24765 4029 24799 4063
rect 25317 4029 25351 4063
rect 5169 3961 5203 3995
rect 10229 3961 10263 3995
rect 10505 3961 10539 3995
rect 11057 3961 11091 3995
rect 12161 3961 12195 3995
rect 12529 3961 12563 3995
rect 14093 3961 14127 3995
rect 16393 3961 16427 3995
rect 17313 3961 17347 3995
rect 17681 3961 17715 3995
rect 17773 3961 17807 3995
rect 19613 3961 19647 3995
rect 19705 3961 19739 3995
rect 21637 3961 21671 3995
rect 22189 3961 22223 3995
rect 23293 3961 23327 3995
rect 23385 3961 23419 3995
rect 3375 3893 3409 3927
rect 3789 3893 3823 3927
rect 4387 3893 4421 3927
rect 4801 3893 4835 3927
rect 5399 3893 5433 3927
rect 5721 3893 5755 3927
rect 6733 3893 6767 3927
rect 9033 3893 9067 3927
rect 13725 3893 13759 3927
rect 14921 3893 14955 3927
rect 19429 3893 19463 3927
rect 24949 3893 24983 3927
rect 4019 3689 4053 3723
rect 6043 3689 6077 3723
rect 8067 3689 8101 3723
rect 10689 3689 10723 3723
rect 12437 3689 12471 3723
rect 14185 3689 14219 3723
rect 15289 3689 15323 3723
rect 16853 3689 16887 3723
rect 21453 3689 21487 3723
rect 9861 3621 9895 3655
rect 11425 3621 11459 3655
rect 16025 3621 16059 3655
rect 17589 3621 17623 3655
rect 20257 3621 20291 3655
rect 20533 3621 20567 3655
rect 20625 3621 20659 3655
rect 22189 3621 22223 3655
rect 23753 3621 23787 3655
rect 3948 3553 3982 3587
rect 4960 3553 4994 3587
rect 5972 3553 6006 3587
rect 7996 3553 8030 3587
rect 13541 3553 13575 3587
rect 14896 3553 14930 3587
rect 18969 3553 19003 3587
rect 6917 3485 6951 3519
rect 9769 3485 9803 3519
rect 10229 3485 10263 3519
rect 11149 3485 11183 3519
rect 11333 3485 11367 3519
rect 11977 3485 12011 3519
rect 12713 3485 12747 3519
rect 15933 3485 15967 3519
rect 16209 3485 16243 3519
rect 17313 3485 17347 3519
rect 17497 3485 17531 3519
rect 20809 3485 20843 3519
rect 22097 3485 22131 3519
rect 22373 3485 22407 3519
rect 23661 3485 23695 3519
rect 23937 3485 23971 3519
rect 18049 3417 18083 3451
rect 19521 3417 19555 3451
rect 5031 3349 5065 3383
rect 9493 3349 9527 3383
rect 13633 3349 13667 3383
rect 14967 3349 15001 3383
rect 18417 3349 18451 3383
rect 19153 3349 19187 3383
rect 23201 3349 23235 3383
rect 2777 3145 2811 3179
rect 3375 3145 3409 3179
rect 3789 3145 3823 3179
rect 4065 3145 4099 3179
rect 4387 3145 4421 3179
rect 5077 3145 5111 3179
rect 5813 3145 5847 3179
rect 6089 3145 6123 3179
rect 9217 3145 9251 3179
rect 10137 3145 10171 3179
rect 11793 3145 11827 3179
rect 13173 3145 13207 3179
rect 13633 3145 13667 3179
rect 15749 3145 15783 3179
rect 17037 3145 17071 3179
rect 20349 3145 20383 3179
rect 23017 3145 23051 3179
rect 24581 3145 24615 3179
rect 24949 3145 24983 3179
rect 9447 3077 9481 3111
rect 22373 3077 22407 3111
rect 24213 3077 24247 3111
rect 8849 3009 8883 3043
rect 10413 3009 10447 3043
rect 11057 3009 11091 3043
rect 12069 3009 12103 3043
rect 12345 3009 12379 3043
rect 13817 3009 13851 3043
rect 14277 3009 14311 3043
rect 17681 3009 17715 3043
rect 18049 3009 18083 3043
rect 19705 3009 19739 3043
rect 21545 3009 21579 3043
rect 2276 2941 2310 2975
rect 3304 2941 3338 2975
rect 4284 2941 4318 2975
rect 4709 2941 4743 2975
rect 5312 2941 5346 2975
rect 7193 2941 7227 2975
rect 7320 2941 7354 2975
rect 8343 2941 8377 2975
rect 8435 2941 8469 2975
rect 9376 2941 9410 2975
rect 15473 2941 15507 2975
rect 16485 2941 16519 2975
rect 23293 2941 23327 2975
rect 24765 2941 24799 2975
rect 25317 2941 25351 2975
rect 2363 2873 2397 2907
rect 5399 2873 5433 2907
rect 9861 2873 9895 2907
rect 10505 2873 10539 2907
rect 12161 2873 12195 2907
rect 13909 2873 13943 2907
rect 14921 2873 14955 2907
rect 16669 2873 16703 2907
rect 17313 2873 17347 2907
rect 17773 2873 17807 2907
rect 18785 2873 18819 2907
rect 19337 2873 19371 2907
rect 19429 2873 19463 2907
rect 20901 2873 20935 2907
rect 20993 2873 21027 2907
rect 23201 2873 23235 2907
rect 7423 2805 7457 2839
rect 8021 2805 8055 2839
rect 11333 2805 11367 2839
rect 19153 2805 19187 2839
rect 20717 2805 20751 2839
rect 22097 2805 22131 2839
rect 1627 2601 1661 2635
rect 4479 2601 4513 2635
rect 7331 2601 7365 2635
rect 7745 2601 7779 2635
rect 8343 2601 8377 2635
rect 9631 2601 9665 2635
rect 13265 2601 13299 2635
rect 14829 2601 14863 2635
rect 16117 2601 16151 2635
rect 23385 2601 23419 2635
rect 25271 2601 25305 2635
rect 9125 2533 9159 2567
rect 11977 2533 12011 2567
rect 12345 2533 12379 2567
rect 15013 2533 15047 2567
rect 18325 2533 18359 2567
rect 18601 2533 18635 2567
rect 20717 2533 20751 2567
rect 23569 2533 23603 2567
rect 1556 2465 1590 2499
rect 2568 2465 2602 2499
rect 4376 2465 4410 2499
rect 4801 2465 4835 2499
rect 7260 2465 7294 2499
rect 8272 2465 8306 2499
rect 9560 2465 9594 2499
rect 10689 2465 10723 2499
rect 13817 2465 13851 2499
rect 14369 2465 14403 2499
rect 15105 2465 15139 2499
rect 16669 2465 16703 2499
rect 17221 2465 17255 2499
rect 20533 2465 20567 2499
rect 20809 2465 20843 2499
rect 22281 2465 22315 2499
rect 22833 2465 22867 2499
rect 23661 2465 23695 2499
rect 25168 2465 25202 2499
rect 25593 2465 25627 2499
rect 5353 2397 5387 2431
rect 10413 2397 10447 2431
rect 10505 2397 10539 2431
rect 11517 2397 11551 2431
rect 12253 2397 12287 2431
rect 12529 2397 12563 2431
rect 18509 2397 18543 2431
rect 16853 2329 16887 2363
rect 19061 2329 19095 2363
rect 2041 2261 2075 2295
rect 2639 2261 2673 2295
rect 3053 2261 3087 2295
rect 8757 2261 8791 2295
rect 10045 2261 10079 2295
rect 14001 2261 14035 2295
rect 17589 2261 17623 2295
rect 19429 2261 19463 2295
rect 20073 2261 20107 2295
rect 22465 2261 22499 2295
<< metal1 >>
rect 3682 27412 3688 27464
rect 3740 27452 3746 27464
rect 4786 27452 4792 27464
rect 3740 27424 4792 27452
rect 3740 27412 3746 27424
rect 4786 27412 4792 27424
rect 4844 27412 4850 27464
rect 632 25594 26392 25616
rect 632 25542 9843 25594
rect 9895 25542 9907 25594
rect 9959 25542 9971 25594
rect 10023 25542 10035 25594
rect 10087 25542 19176 25594
rect 19228 25542 19240 25594
rect 19292 25542 19304 25594
rect 19356 25542 19368 25594
rect 19420 25542 26392 25594
rect 632 25520 26392 25542
rect 632 25050 26392 25072
rect 632 24998 5176 25050
rect 5228 24998 5240 25050
rect 5292 24998 5304 25050
rect 5356 24998 5368 25050
rect 5420 24998 14510 25050
rect 14562 24998 14574 25050
rect 14626 24998 14638 25050
rect 14690 24998 14702 25050
rect 14754 24998 23843 25050
rect 23895 24998 23907 25050
rect 23959 24998 23971 25050
rect 24023 24998 24035 25050
rect 24087 24998 26392 25050
rect 632 24976 26392 24998
rect 632 24506 26392 24528
rect 632 24454 9843 24506
rect 9895 24454 9907 24506
rect 9959 24454 9971 24506
rect 10023 24454 10035 24506
rect 10087 24454 19176 24506
rect 19228 24454 19240 24506
rect 19292 24454 19304 24506
rect 19356 24454 19368 24506
rect 19420 24454 26392 24506
rect 632 24432 26392 24454
rect 632 23962 26392 23984
rect 632 23910 5176 23962
rect 5228 23910 5240 23962
rect 5292 23910 5304 23962
rect 5356 23910 5368 23962
rect 5420 23910 14510 23962
rect 14562 23910 14574 23962
rect 14626 23910 14638 23962
rect 14690 23910 14702 23962
rect 14754 23910 23843 23962
rect 23895 23910 23907 23962
rect 23959 23910 23971 23962
rect 24023 23910 24035 23962
rect 24087 23910 26392 23962
rect 632 23888 26392 23910
rect 24290 23808 24296 23860
rect 24348 23848 24354 23860
rect 24569 23851 24627 23857
rect 24569 23848 24581 23851
rect 24348 23820 24581 23848
rect 24348 23808 24354 23820
rect 24569 23817 24581 23820
rect 24615 23817 24627 23851
rect 24569 23811 24627 23817
rect 21717 23783 21775 23789
rect 21717 23749 21729 23783
rect 21763 23780 21775 23783
rect 22910 23780 22916 23792
rect 21763 23752 22916 23780
rect 21763 23749 21775 23752
rect 21717 23743 21775 23749
rect 21232 23647 21290 23653
rect 21232 23613 21244 23647
rect 21278 23644 21290 23647
rect 21732 23644 21760 23743
rect 22910 23740 22916 23752
rect 22968 23740 22974 23792
rect 21278 23616 21760 23644
rect 24176 23647 24234 23653
rect 21278 23613 21290 23616
rect 21232 23607 21290 23613
rect 24176 23613 24188 23647
rect 24222 23644 24234 23647
rect 24290 23644 24296 23656
rect 24222 23616 24296 23644
rect 24222 23613 24234 23616
rect 24176 23607 24234 23613
rect 24290 23604 24296 23616
rect 24348 23604 24354 23656
rect 20334 23468 20340 23520
rect 20392 23508 20398 23520
rect 21303 23511 21361 23517
rect 21303 23508 21315 23511
rect 20392 23480 21315 23508
rect 20392 23468 20398 23480
rect 21303 23477 21315 23480
rect 21349 23477 21361 23511
rect 21303 23471 21361 23477
rect 23002 23468 23008 23520
rect 23060 23508 23066 23520
rect 24247 23511 24305 23517
rect 24247 23508 24259 23511
rect 23060 23480 24259 23508
rect 23060 23468 23066 23480
rect 24247 23477 24259 23480
rect 24293 23477 24305 23511
rect 24247 23471 24305 23477
rect 632 23418 26392 23440
rect 632 23366 9843 23418
rect 9895 23366 9907 23418
rect 9959 23366 9971 23418
rect 10023 23366 10035 23418
rect 10087 23366 19176 23418
rect 19228 23366 19240 23418
rect 19292 23366 19304 23418
rect 19356 23366 19368 23418
rect 19420 23366 26392 23418
rect 632 23344 26392 23366
rect 632 22874 26392 22896
rect 632 22822 5176 22874
rect 5228 22822 5240 22874
rect 5292 22822 5304 22874
rect 5356 22822 5368 22874
rect 5420 22822 14510 22874
rect 14562 22822 14574 22874
rect 14626 22822 14638 22874
rect 14690 22822 14702 22874
rect 14754 22822 23843 22874
rect 23895 22822 23907 22874
rect 23959 22822 23971 22874
rect 24023 22822 24035 22874
rect 24087 22822 26392 22874
rect 632 22800 26392 22822
rect 632 22330 26392 22352
rect 632 22278 9843 22330
rect 9895 22278 9907 22330
rect 9959 22278 9971 22330
rect 10023 22278 10035 22330
rect 10087 22278 19176 22330
rect 19228 22278 19240 22330
rect 19292 22278 19304 22330
rect 19356 22278 19368 22330
rect 19420 22278 26392 22330
rect 632 22256 26392 22278
rect 632 21786 26392 21808
rect 632 21734 5176 21786
rect 5228 21734 5240 21786
rect 5292 21734 5304 21786
rect 5356 21734 5368 21786
rect 5420 21734 14510 21786
rect 14562 21734 14574 21786
rect 14626 21734 14638 21786
rect 14690 21734 14702 21786
rect 14754 21734 23843 21786
rect 23895 21734 23907 21786
rect 23959 21734 23971 21786
rect 24023 21734 24035 21786
rect 24087 21734 26392 21786
rect 632 21712 26392 21734
rect 24290 21632 24296 21684
rect 24348 21672 24354 21684
rect 24569 21675 24627 21681
rect 24569 21672 24581 21675
rect 24348 21644 24581 21672
rect 24348 21632 24354 21644
rect 24569 21641 24581 21644
rect 24615 21641 24627 21675
rect 24569 21635 24627 21641
rect 24176 21471 24234 21477
rect 24176 21437 24188 21471
rect 24222 21468 24234 21471
rect 24290 21468 24296 21480
rect 24222 21440 24296 21468
rect 24222 21437 24234 21440
rect 24176 21431 24234 21437
rect 24290 21428 24296 21440
rect 24348 21428 24354 21480
rect 22358 21292 22364 21344
rect 22416 21332 22422 21344
rect 24247 21335 24305 21341
rect 24247 21332 24259 21335
rect 22416 21304 24259 21332
rect 22416 21292 22422 21304
rect 24247 21301 24259 21304
rect 24293 21301 24305 21335
rect 24247 21295 24305 21301
rect 632 21242 26392 21264
rect 632 21190 9843 21242
rect 9895 21190 9907 21242
rect 9959 21190 9971 21242
rect 10023 21190 10035 21242
rect 10087 21190 19176 21242
rect 19228 21190 19240 21242
rect 19292 21190 19304 21242
rect 19356 21190 19368 21242
rect 19420 21190 26392 21242
rect 632 21168 26392 21190
rect 24198 21001 24204 21004
rect 24176 20995 24204 21001
rect 24176 20961 24188 20995
rect 24176 20955 24204 20961
rect 24198 20952 24204 20955
rect 24256 20952 24262 21004
rect 23278 20748 23284 20800
rect 23336 20788 23342 20800
rect 24247 20791 24305 20797
rect 24247 20788 24259 20791
rect 23336 20760 24259 20788
rect 23336 20748 23342 20760
rect 24247 20757 24259 20760
rect 24293 20757 24305 20791
rect 24247 20751 24305 20757
rect 632 20698 26392 20720
rect 632 20646 5176 20698
rect 5228 20646 5240 20698
rect 5292 20646 5304 20698
rect 5356 20646 5368 20698
rect 5420 20646 14510 20698
rect 14562 20646 14574 20698
rect 14626 20646 14638 20698
rect 14690 20646 14702 20698
rect 14754 20646 23843 20698
rect 23895 20646 23907 20698
rect 23959 20646 23971 20698
rect 24023 20646 24035 20698
rect 24087 20646 26392 20698
rect 632 20624 26392 20646
rect 24198 20584 24204 20596
rect 24159 20556 24204 20584
rect 24198 20544 24204 20556
rect 24256 20544 24262 20596
rect 632 20154 26392 20176
rect 632 20102 9843 20154
rect 9895 20102 9907 20154
rect 9959 20102 9971 20154
rect 10023 20102 10035 20154
rect 10087 20102 19176 20154
rect 19228 20102 19240 20154
rect 19292 20102 19304 20154
rect 19356 20102 19368 20154
rect 19420 20102 26392 20154
rect 632 20080 26392 20102
rect 24176 19907 24234 19913
rect 24176 19873 24188 19907
rect 24222 19904 24234 19907
rect 25026 19904 25032 19916
rect 24222 19876 25032 19904
rect 24222 19873 24234 19876
rect 24176 19867 24234 19873
rect 25026 19864 25032 19876
rect 25084 19864 25090 19916
rect 23002 19660 23008 19712
rect 23060 19700 23066 19712
rect 24247 19703 24305 19709
rect 24247 19700 24259 19703
rect 23060 19672 24259 19700
rect 23060 19660 23066 19672
rect 24247 19669 24259 19672
rect 24293 19669 24305 19703
rect 24247 19663 24305 19669
rect 632 19610 26392 19632
rect 632 19558 5176 19610
rect 5228 19558 5240 19610
rect 5292 19558 5304 19610
rect 5356 19558 5368 19610
rect 5420 19558 14510 19610
rect 14562 19558 14574 19610
rect 14626 19558 14638 19610
rect 14690 19558 14702 19610
rect 14754 19558 23843 19610
rect 23895 19558 23907 19610
rect 23959 19558 23971 19610
rect 24023 19558 24035 19610
rect 24087 19558 26392 19610
rect 632 19536 26392 19558
rect 24160 19295 24218 19301
rect 24160 19261 24172 19295
rect 24206 19292 24218 19295
rect 25026 19292 25032 19304
rect 24206 19264 24704 19292
rect 24987 19264 25032 19292
rect 24206 19261 24218 19264
rect 24160 19255 24218 19261
rect 23002 19184 23008 19236
rect 23060 19224 23066 19236
rect 24247 19227 24305 19233
rect 24247 19224 24259 19227
rect 23060 19196 24259 19224
rect 23060 19184 23066 19196
rect 24247 19193 24259 19196
rect 24293 19193 24305 19227
rect 24247 19187 24305 19193
rect 24676 19165 24704 19264
rect 25026 19252 25032 19264
rect 25084 19252 25090 19304
rect 24661 19159 24719 19165
rect 24661 19125 24673 19159
rect 24707 19156 24719 19159
rect 25486 19156 25492 19168
rect 24707 19128 25492 19156
rect 24707 19125 24719 19128
rect 24661 19119 24719 19125
rect 25486 19116 25492 19128
rect 25544 19116 25550 19168
rect 632 19066 26392 19088
rect 632 19014 9843 19066
rect 9895 19014 9907 19066
rect 9959 19014 9971 19066
rect 10023 19014 10035 19066
rect 10087 19014 19176 19066
rect 19228 19014 19240 19066
rect 19292 19014 19304 19066
rect 19356 19014 19368 19066
rect 19420 19014 26392 19066
rect 632 18992 26392 19014
rect 20518 18825 20524 18828
rect 20496 18819 20524 18825
rect 20496 18785 20508 18819
rect 20496 18779 20524 18785
rect 20518 18776 20524 18779
rect 20576 18776 20582 18828
rect 23164 18819 23222 18825
rect 23164 18785 23176 18819
rect 23210 18816 23222 18819
rect 23462 18816 23468 18828
rect 23210 18788 23468 18816
rect 23210 18785 23222 18788
rect 23164 18779 23222 18785
rect 23462 18776 23468 18788
rect 23520 18776 23526 18828
rect 24176 18819 24234 18825
rect 24176 18785 24188 18819
rect 24222 18816 24234 18819
rect 25026 18816 25032 18828
rect 24222 18788 25032 18816
rect 24222 18785 24234 18788
rect 24176 18779 24234 18785
rect 25026 18776 25032 18788
rect 25084 18776 25090 18828
rect 23002 18640 23008 18692
rect 23060 18680 23066 18692
rect 23235 18683 23293 18689
rect 23235 18680 23247 18683
rect 23060 18652 23247 18680
rect 23060 18640 23066 18652
rect 23235 18649 23247 18652
rect 23281 18649 23293 18683
rect 23235 18643 23293 18649
rect 20518 18572 20524 18624
rect 20576 18621 20582 18624
rect 20576 18615 20625 18621
rect 20576 18581 20579 18615
rect 20613 18581 20625 18615
rect 20576 18575 20625 18581
rect 20576 18572 20582 18575
rect 23094 18572 23100 18624
rect 23152 18612 23158 18624
rect 24247 18615 24305 18621
rect 24247 18612 24259 18615
rect 23152 18584 24259 18612
rect 23152 18572 23158 18584
rect 24247 18581 24259 18584
rect 24293 18581 24305 18615
rect 24247 18575 24305 18581
rect 632 18522 26392 18544
rect 632 18470 5176 18522
rect 5228 18470 5240 18522
rect 5292 18470 5304 18522
rect 5356 18470 5368 18522
rect 5420 18470 14510 18522
rect 14562 18470 14574 18522
rect 14626 18470 14638 18522
rect 14690 18470 14702 18522
rect 14754 18470 23843 18522
rect 23895 18470 23907 18522
rect 23959 18470 23971 18522
rect 24023 18470 24035 18522
rect 24087 18470 26392 18522
rect 632 18448 26392 18470
rect 20426 18408 20432 18420
rect 20387 18380 20432 18408
rect 20426 18368 20432 18380
rect 20484 18368 20490 18420
rect 23462 18272 23468 18284
rect 23375 18244 23468 18272
rect 23462 18232 23468 18244
rect 23520 18272 23526 18284
rect 24290 18272 24296 18284
rect 23520 18244 24296 18272
rect 23520 18232 23526 18244
rect 24290 18232 24296 18244
rect 24348 18232 24354 18284
rect 22152 18207 22210 18213
rect 22152 18173 22164 18207
rect 22198 18204 22210 18207
rect 24176 18207 24234 18213
rect 22198 18176 22680 18204
rect 22198 18173 22210 18176
rect 22152 18167 22210 18173
rect 22652 18080 22680 18176
rect 24176 18173 24188 18207
rect 24222 18204 24234 18207
rect 24222 18173 24244 18204
rect 24176 18167 24244 18173
rect 23646 18096 23652 18148
rect 23704 18136 23710 18148
rect 24216 18136 24244 18167
rect 25118 18164 25124 18216
rect 25176 18213 25182 18216
rect 25176 18207 25214 18213
rect 25202 18204 25214 18207
rect 25581 18207 25639 18213
rect 25581 18204 25593 18207
rect 25202 18176 25593 18204
rect 25202 18173 25214 18176
rect 25176 18167 25214 18173
rect 25581 18173 25593 18176
rect 25627 18173 25639 18207
rect 25581 18167 25639 18173
rect 25176 18164 25182 18167
rect 24569 18139 24627 18145
rect 24569 18136 24581 18139
rect 23704 18108 24581 18136
rect 23704 18096 23710 18108
rect 24569 18105 24581 18108
rect 24615 18105 24627 18139
rect 24569 18099 24627 18105
rect 22082 18028 22088 18080
rect 22140 18068 22146 18080
rect 22223 18071 22281 18077
rect 22223 18068 22235 18071
rect 22140 18040 22235 18068
rect 22140 18028 22146 18040
rect 22223 18037 22235 18040
rect 22269 18037 22281 18071
rect 22634 18068 22640 18080
rect 22595 18040 22640 18068
rect 22223 18031 22281 18037
rect 22634 18028 22640 18040
rect 22692 18028 22698 18080
rect 23462 18028 23468 18080
rect 23520 18068 23526 18080
rect 24247 18071 24305 18077
rect 24247 18068 24259 18071
rect 23520 18040 24259 18068
rect 23520 18028 23526 18040
rect 24247 18037 24259 18040
rect 24293 18037 24305 18071
rect 25026 18068 25032 18080
rect 24987 18040 25032 18068
rect 24247 18031 24305 18037
rect 25026 18028 25032 18040
rect 25084 18028 25090 18080
rect 25210 18028 25216 18080
rect 25268 18077 25274 18080
rect 25268 18071 25317 18077
rect 25268 18037 25271 18071
rect 25305 18037 25317 18071
rect 25268 18031 25317 18037
rect 25268 18028 25274 18031
rect 632 17978 26392 18000
rect 632 17926 9843 17978
rect 9895 17926 9907 17978
rect 9959 17926 9971 17978
rect 10023 17926 10035 17978
rect 10087 17926 19176 17978
rect 19228 17926 19240 17978
rect 19292 17926 19304 17978
rect 19356 17926 19368 17978
rect 19420 17926 26392 17978
rect 632 17904 26392 17926
rect 21530 17864 21536 17876
rect 21491 17836 21536 17864
rect 21530 17824 21536 17836
rect 21588 17824 21594 17876
rect 20426 17688 20432 17740
rect 20484 17728 20490 17740
rect 20521 17731 20579 17737
rect 20521 17728 20533 17731
rect 20484 17700 20533 17728
rect 20484 17688 20490 17700
rect 20521 17697 20533 17700
rect 20567 17697 20579 17731
rect 20521 17691 20579 17697
rect 22637 17731 22695 17737
rect 22637 17697 22649 17731
rect 22683 17728 22695 17731
rect 22726 17728 22732 17740
rect 22683 17700 22732 17728
rect 22683 17697 22695 17700
rect 22637 17691 22695 17697
rect 22726 17688 22732 17700
rect 22784 17688 22790 17740
rect 24198 17737 24204 17740
rect 24176 17731 24204 17737
rect 24176 17697 24188 17731
rect 24176 17691 24204 17697
rect 24198 17688 24204 17691
rect 24256 17688 24262 17740
rect 20702 17524 20708 17536
rect 20663 17496 20708 17524
rect 20702 17484 20708 17496
rect 20760 17484 20766 17536
rect 22174 17484 22180 17536
rect 22232 17524 22238 17536
rect 22269 17527 22327 17533
rect 22269 17524 22281 17527
rect 22232 17496 22281 17524
rect 22232 17484 22238 17496
rect 22269 17493 22281 17496
rect 22315 17493 22327 17527
rect 22269 17487 22327 17493
rect 23002 17484 23008 17536
rect 23060 17524 23066 17536
rect 24247 17527 24305 17533
rect 24247 17524 24259 17527
rect 23060 17496 24259 17524
rect 23060 17484 23066 17496
rect 24247 17493 24259 17496
rect 24293 17493 24305 17527
rect 24247 17487 24305 17493
rect 632 17434 26392 17456
rect 632 17382 5176 17434
rect 5228 17382 5240 17434
rect 5292 17382 5304 17434
rect 5356 17382 5368 17434
rect 5420 17382 14510 17434
rect 14562 17382 14574 17434
rect 14626 17382 14638 17434
rect 14690 17382 14702 17434
rect 14754 17382 23843 17434
rect 23895 17382 23907 17434
rect 23959 17382 23971 17434
rect 24023 17382 24035 17434
rect 24087 17382 26392 17434
rect 632 17360 26392 17382
rect 24198 17320 24204 17332
rect 24159 17292 24204 17320
rect 24198 17280 24204 17292
rect 24256 17280 24262 17332
rect 21530 17252 21536 17264
rect 21272 17224 21536 17252
rect 21272 17193 21300 17224
rect 21530 17212 21536 17224
rect 21588 17212 21594 17264
rect 21257 17187 21315 17193
rect 21257 17153 21269 17187
rect 21303 17153 21315 17187
rect 21257 17147 21315 17153
rect 21622 17144 21628 17196
rect 21680 17184 21686 17196
rect 21680 17156 21725 17184
rect 21680 17144 21686 17156
rect 15737 17119 15795 17125
rect 15737 17085 15749 17119
rect 15783 17116 15795 17119
rect 15921 17119 15979 17125
rect 15921 17116 15933 17119
rect 15783 17088 15933 17116
rect 15783 17085 15795 17088
rect 15737 17079 15795 17085
rect 15921 17085 15933 17088
rect 15967 17116 15979 17119
rect 16194 17116 16200 17128
rect 15967 17088 16200 17116
rect 15967 17085 15979 17088
rect 15921 17079 15979 17085
rect 16194 17076 16200 17088
rect 16252 17076 16258 17128
rect 19509 17119 19567 17125
rect 19509 17085 19521 17119
rect 19555 17116 19567 17119
rect 19693 17119 19751 17125
rect 19693 17116 19705 17119
rect 19555 17088 19705 17116
rect 19555 17085 19567 17088
rect 19509 17079 19567 17085
rect 19693 17085 19705 17088
rect 19739 17116 19751 17119
rect 19966 17116 19972 17128
rect 19739 17088 19972 17116
rect 19739 17085 19751 17088
rect 19693 17079 19751 17085
rect 19966 17076 19972 17088
rect 20024 17076 20030 17128
rect 24712 17119 24770 17125
rect 24712 17085 24724 17119
rect 24758 17116 24770 17119
rect 24758 17088 24923 17116
rect 24758 17085 24770 17088
rect 24712 17079 24770 17085
rect 16562 17048 16568 17060
rect 16523 17020 16568 17048
rect 16562 17008 16568 17020
rect 16620 17008 16626 17060
rect 21349 17051 21407 17057
rect 21349 17017 21361 17051
rect 21395 17017 21407 17051
rect 21349 17011 21407 17017
rect 20061 16983 20119 16989
rect 20061 16949 20073 16983
rect 20107 16980 20119 16983
rect 20150 16980 20156 16992
rect 20107 16952 20156 16980
rect 20107 16949 20119 16952
rect 20061 16943 20119 16949
rect 20150 16940 20156 16952
rect 20208 16940 20214 16992
rect 20426 16940 20432 16992
rect 20484 16980 20490 16992
rect 20613 16983 20671 16989
rect 20613 16980 20625 16983
rect 20484 16952 20625 16980
rect 20484 16940 20490 16952
rect 20613 16949 20625 16952
rect 20659 16980 20671 16983
rect 20981 16983 21039 16989
rect 20981 16980 20993 16983
rect 20659 16952 20993 16980
rect 20659 16949 20671 16952
rect 20613 16943 20671 16949
rect 20981 16949 20993 16952
rect 21027 16980 21039 16983
rect 21364 16980 21392 17011
rect 24382 17008 24388 17060
rect 24440 17048 24446 17060
rect 24799 17051 24857 17057
rect 24799 17048 24811 17051
rect 24440 17020 24811 17048
rect 24440 17008 24446 17020
rect 24799 17017 24811 17020
rect 24845 17017 24857 17051
rect 24799 17011 24857 17017
rect 21027 16952 21392 16980
rect 22269 16983 22327 16989
rect 21027 16949 21039 16952
rect 20981 16943 21039 16949
rect 22269 16949 22281 16983
rect 22315 16980 22327 16983
rect 22726 16980 22732 16992
rect 22315 16952 22732 16980
rect 22315 16949 22327 16952
rect 22269 16943 22327 16949
rect 22726 16940 22732 16952
rect 22784 16940 22790 16992
rect 23370 16940 23376 16992
rect 23428 16980 23434 16992
rect 23649 16983 23707 16989
rect 23649 16980 23661 16983
rect 23428 16952 23661 16980
rect 23428 16940 23434 16952
rect 23649 16949 23661 16952
rect 23695 16949 23707 16983
rect 23649 16943 23707 16949
rect 24290 16940 24296 16992
rect 24348 16980 24354 16992
rect 24895 16980 24923 17088
rect 25121 16983 25179 16989
rect 25121 16980 25133 16983
rect 24348 16952 25133 16980
rect 24348 16940 24354 16952
rect 25121 16949 25133 16952
rect 25167 16949 25179 16983
rect 25121 16943 25179 16949
rect 632 16890 26392 16912
rect 632 16838 9843 16890
rect 9895 16838 9907 16890
rect 9959 16838 9971 16890
rect 10023 16838 10035 16890
rect 10087 16838 19176 16890
rect 19228 16838 19240 16890
rect 19292 16838 19304 16890
rect 19356 16838 19368 16890
rect 19420 16838 26392 16890
rect 632 16816 26392 16838
rect 15642 16736 15648 16788
rect 15700 16776 15706 16788
rect 16010 16776 16016 16788
rect 15700 16748 16016 16776
rect 15700 16736 15706 16748
rect 16010 16736 16016 16748
rect 16068 16736 16074 16788
rect 18405 16779 18463 16785
rect 18405 16745 18417 16779
rect 18451 16776 18463 16779
rect 18678 16776 18684 16788
rect 18451 16748 18684 16776
rect 18451 16745 18463 16748
rect 18405 16739 18463 16745
rect 18678 16736 18684 16748
rect 18736 16736 18742 16788
rect 16562 16668 16568 16720
rect 16620 16708 16626 16720
rect 16657 16711 16715 16717
rect 16657 16708 16669 16711
rect 16620 16680 16669 16708
rect 16620 16668 16626 16680
rect 16657 16677 16669 16680
rect 16703 16677 16715 16711
rect 16657 16671 16715 16677
rect 20702 16668 20708 16720
rect 20760 16708 20766 16720
rect 20797 16711 20855 16717
rect 20797 16708 20809 16711
rect 20760 16680 20809 16708
rect 20760 16668 20766 16680
rect 20797 16677 20809 16680
rect 20843 16677 20855 16711
rect 20797 16671 20855 16677
rect 24382 16668 24388 16720
rect 24440 16708 24446 16720
rect 24891 16711 24949 16717
rect 24891 16708 24903 16711
rect 24440 16680 24903 16708
rect 24440 16668 24446 16680
rect 24891 16677 24903 16680
rect 24937 16677 24949 16711
rect 24891 16671 24949 16677
rect 14906 16640 14912 16652
rect 14867 16612 14912 16640
rect 14906 16600 14912 16612
rect 14964 16600 14970 16652
rect 15553 16643 15611 16649
rect 15553 16609 15565 16643
rect 15599 16640 15611 16643
rect 15734 16640 15740 16652
rect 15599 16612 15740 16640
rect 15599 16609 15611 16612
rect 15553 16603 15611 16609
rect 15734 16600 15740 16612
rect 15792 16600 15798 16652
rect 18218 16640 18224 16652
rect 18179 16612 18224 16640
rect 18218 16600 18224 16612
rect 18276 16600 18282 16652
rect 22542 16640 22548 16652
rect 22503 16612 22548 16640
rect 22542 16600 22548 16612
rect 22600 16600 22606 16652
rect 23738 16600 23744 16652
rect 23796 16649 23802 16652
rect 23796 16643 23834 16649
rect 23822 16609 23834 16643
rect 23796 16603 23834 16609
rect 23879 16643 23937 16649
rect 23879 16609 23891 16643
rect 23925 16640 23937 16643
rect 24198 16640 24204 16652
rect 23925 16612 24204 16640
rect 23925 16609 23937 16612
rect 23879 16603 23937 16609
rect 23796 16600 23802 16603
rect 24198 16600 24204 16612
rect 24256 16600 24262 16652
rect 24804 16643 24862 16649
rect 24804 16609 24816 16643
rect 24850 16640 24862 16643
rect 25394 16640 25400 16652
rect 24850 16612 25400 16640
rect 24850 16609 24862 16612
rect 24804 16603 24862 16609
rect 25394 16600 25400 16612
rect 25452 16600 25458 16652
rect 16565 16575 16623 16581
rect 16565 16541 16577 16575
rect 16611 16572 16623 16575
rect 16654 16572 16660 16584
rect 16611 16544 16660 16572
rect 16611 16541 16623 16544
rect 16565 16535 16623 16541
rect 16654 16532 16660 16544
rect 16712 16532 16718 16584
rect 16838 16572 16844 16584
rect 16799 16544 16844 16572
rect 16838 16532 16844 16544
rect 16896 16532 16902 16584
rect 20242 16532 20248 16584
rect 20300 16572 20306 16584
rect 20705 16575 20763 16581
rect 20705 16572 20717 16575
rect 20300 16544 20717 16572
rect 20300 16532 20306 16544
rect 20705 16541 20717 16544
rect 20751 16541 20763 16575
rect 20705 16535 20763 16541
rect 21349 16575 21407 16581
rect 21349 16541 21361 16575
rect 21395 16572 21407 16575
rect 21438 16572 21444 16584
rect 21395 16544 21444 16572
rect 21395 16541 21407 16544
rect 21349 16535 21407 16541
rect 21438 16532 21444 16544
rect 21496 16572 21502 16584
rect 21622 16572 21628 16584
rect 21496 16544 21628 16572
rect 21496 16532 21502 16544
rect 21622 16532 21628 16544
rect 21680 16532 21686 16584
rect 19506 16436 19512 16448
rect 19467 16408 19512 16436
rect 19506 16396 19512 16408
rect 19564 16396 19570 16448
rect 22450 16436 22456 16448
rect 22411 16408 22456 16436
rect 22450 16396 22456 16408
rect 22508 16396 22514 16448
rect 632 16346 26392 16368
rect 632 16294 5176 16346
rect 5228 16294 5240 16346
rect 5292 16294 5304 16346
rect 5356 16294 5368 16346
rect 5420 16294 14510 16346
rect 14562 16294 14574 16346
rect 14626 16294 14638 16346
rect 14690 16294 14702 16346
rect 14754 16294 23843 16346
rect 23895 16294 23907 16346
rect 23959 16294 23971 16346
rect 24023 16294 24035 16346
rect 24087 16294 26392 16346
rect 632 16272 26392 16294
rect 16562 16232 16568 16244
rect 16523 16204 16568 16232
rect 16562 16192 16568 16204
rect 16620 16192 16626 16244
rect 20426 16232 20432 16244
rect 20387 16204 20432 16232
rect 20426 16192 20432 16204
rect 20484 16192 20490 16244
rect 20702 16232 20708 16244
rect 20663 16204 20708 16232
rect 20702 16192 20708 16204
rect 20760 16192 20766 16244
rect 21441 16235 21499 16241
rect 21441 16201 21453 16235
rect 21487 16232 21499 16235
rect 21714 16232 21720 16244
rect 21487 16204 21720 16232
rect 21487 16201 21499 16204
rect 21441 16195 21499 16201
rect 21714 16192 21720 16204
rect 21772 16232 21778 16244
rect 22542 16232 22548 16244
rect 21772 16204 22548 16232
rect 21772 16192 21778 16204
rect 22542 16192 22548 16204
rect 22600 16192 22606 16244
rect 14541 16099 14599 16105
rect 14541 16065 14553 16099
rect 14587 16096 14599 16099
rect 16654 16096 16660 16108
rect 14587 16068 16660 16096
rect 14587 16065 14599 16068
rect 14541 16059 14599 16065
rect 16654 16056 16660 16068
rect 16712 16096 16718 16108
rect 16933 16099 16991 16105
rect 16933 16096 16945 16099
rect 16712 16068 16945 16096
rect 16712 16056 16718 16068
rect 16933 16065 16945 16068
rect 16979 16065 16991 16099
rect 16933 16059 16991 16065
rect 21438 16056 21444 16108
rect 21496 16096 21502 16108
rect 21625 16099 21683 16105
rect 21625 16096 21637 16099
rect 21496 16068 21637 16096
rect 21496 16056 21502 16068
rect 21625 16065 21637 16068
rect 21671 16065 21683 16099
rect 21625 16059 21683 16065
rect 17390 16028 17396 16040
rect 17303 16000 17396 16028
rect 17390 15988 17396 16000
rect 17448 16028 17454 16040
rect 17669 16031 17727 16037
rect 17669 16028 17681 16031
rect 17448 16000 17681 16028
rect 17448 15988 17454 16000
rect 17669 15997 17681 16000
rect 17715 15997 17727 16031
rect 19506 16028 19512 16040
rect 19467 16000 19512 16028
rect 17669 15991 17727 15997
rect 19506 15988 19512 16000
rect 19564 15988 19570 16040
rect 23005 16031 23063 16037
rect 23005 15997 23017 16031
rect 23051 16028 23063 16031
rect 23278 16028 23284 16040
rect 23051 16000 23284 16028
rect 23051 15997 23063 16000
rect 23005 15991 23063 15997
rect 23278 15988 23284 16000
rect 23336 15988 23342 16040
rect 15642 15960 15648 15972
rect 15603 15932 15648 15960
rect 15642 15920 15648 15932
rect 15700 15920 15706 15972
rect 15734 15920 15740 15972
rect 15792 15960 15798 15972
rect 16289 15963 16347 15969
rect 15792 15932 15837 15960
rect 15792 15920 15798 15932
rect 16289 15929 16301 15963
rect 16335 15960 16347 15963
rect 17114 15960 17120 15972
rect 16335 15932 17120 15960
rect 16335 15929 16347 15932
rect 16289 15923 16347 15929
rect 17114 15920 17120 15932
rect 17172 15920 17178 15972
rect 17577 15963 17635 15969
rect 17577 15929 17589 15963
rect 17623 15929 17635 15963
rect 17577 15923 17635 15929
rect 19417 15963 19475 15969
rect 19417 15929 19429 15963
rect 19463 15960 19475 15963
rect 19871 15963 19929 15969
rect 19871 15960 19883 15963
rect 19463 15932 19883 15960
rect 19463 15929 19475 15932
rect 19417 15923 19475 15929
rect 19871 15929 19883 15932
rect 19917 15960 19929 15963
rect 20886 15960 20892 15972
rect 19917 15932 20892 15960
rect 19917 15929 19929 15932
rect 19871 15923 19929 15929
rect 15093 15895 15151 15901
rect 15093 15861 15105 15895
rect 15139 15892 15151 15895
rect 15461 15895 15519 15901
rect 15461 15892 15473 15895
rect 15139 15864 15473 15892
rect 15139 15861 15151 15864
rect 15093 15855 15151 15861
rect 15461 15861 15473 15864
rect 15507 15892 15519 15895
rect 15752 15892 15780 15920
rect 15507 15864 15780 15892
rect 15507 15861 15519 15864
rect 15461 15855 15519 15861
rect 16746 15852 16752 15904
rect 16804 15892 16810 15904
rect 17592 15892 17620 15923
rect 20886 15920 20892 15932
rect 20944 15920 20950 15972
rect 21714 15960 21720 15972
rect 21675 15932 21720 15960
rect 21714 15920 21720 15932
rect 21772 15920 21778 15972
rect 22269 15963 22327 15969
rect 22269 15929 22281 15963
rect 22315 15960 22327 15963
rect 22542 15960 22548 15972
rect 22315 15932 22548 15960
rect 22315 15929 22327 15932
rect 22269 15923 22327 15929
rect 22542 15920 22548 15932
rect 22600 15960 22606 15972
rect 23738 15960 23744 15972
rect 22600 15932 23744 15960
rect 22600 15920 22606 15932
rect 23738 15920 23744 15932
rect 23796 15960 23802 15972
rect 24201 15963 24259 15969
rect 24201 15960 24213 15963
rect 23796 15932 24213 15960
rect 23796 15920 23802 15932
rect 24201 15929 24213 15932
rect 24247 15929 24259 15963
rect 24201 15923 24259 15929
rect 16804 15864 17620 15892
rect 16804 15852 16810 15864
rect 18218 15852 18224 15904
rect 18276 15892 18282 15904
rect 18681 15895 18739 15901
rect 18681 15892 18693 15895
rect 18276 15864 18693 15892
rect 18276 15852 18282 15864
rect 18681 15861 18693 15864
rect 18727 15892 18739 15895
rect 18770 15892 18776 15904
rect 18727 15864 18776 15892
rect 18727 15861 18739 15864
rect 18681 15855 18739 15861
rect 18770 15852 18776 15864
rect 18828 15852 18834 15904
rect 23465 15895 23523 15901
rect 23465 15861 23477 15895
rect 23511 15892 23523 15895
rect 23554 15892 23560 15904
rect 23511 15864 23560 15892
rect 23511 15861 23523 15864
rect 23465 15855 23523 15861
rect 23554 15852 23560 15864
rect 23612 15852 23618 15904
rect 24750 15892 24756 15904
rect 24711 15864 24756 15892
rect 24750 15852 24756 15864
rect 24808 15852 24814 15904
rect 25305 15895 25363 15901
rect 25305 15861 25317 15895
rect 25351 15892 25363 15895
rect 25394 15892 25400 15904
rect 25351 15864 25400 15892
rect 25351 15861 25363 15864
rect 25305 15855 25363 15861
rect 25394 15852 25400 15864
rect 25452 15852 25458 15904
rect 632 15802 26392 15824
rect 632 15750 9843 15802
rect 9895 15750 9907 15802
rect 9959 15750 9971 15802
rect 10023 15750 10035 15802
rect 10087 15750 19176 15802
rect 19228 15750 19240 15802
rect 19292 15750 19304 15802
rect 19356 15750 19368 15802
rect 19420 15750 26392 15802
rect 632 15728 26392 15750
rect 16194 15688 16200 15700
rect 16155 15660 16200 15688
rect 16194 15648 16200 15660
rect 16252 15688 16258 15700
rect 17022 15688 17028 15700
rect 16252 15660 17028 15688
rect 16252 15648 16258 15660
rect 17022 15648 17028 15660
rect 17080 15688 17086 15700
rect 17080 15660 17252 15688
rect 17080 15648 17086 15660
rect 15639 15623 15697 15629
rect 15639 15589 15651 15623
rect 15685 15620 15697 15623
rect 15918 15620 15924 15632
rect 15685 15592 15924 15620
rect 15685 15589 15697 15592
rect 15639 15583 15697 15589
rect 15918 15580 15924 15592
rect 15976 15580 15982 15632
rect 17224 15629 17252 15660
rect 21438 15648 21444 15700
rect 21496 15688 21502 15700
rect 21625 15691 21683 15697
rect 21625 15688 21637 15691
rect 21496 15660 21637 15688
rect 21496 15648 21502 15660
rect 21625 15657 21637 15660
rect 21671 15657 21683 15691
rect 21625 15651 21683 15657
rect 17209 15623 17267 15629
rect 17209 15589 17221 15623
rect 17255 15589 17267 15623
rect 17209 15583 17267 15589
rect 20791 15623 20849 15629
rect 20791 15589 20803 15623
rect 20837 15620 20849 15623
rect 20886 15620 20892 15632
rect 20837 15592 20892 15620
rect 20837 15589 20849 15592
rect 20791 15583 20849 15589
rect 20886 15580 20892 15592
rect 20944 15580 20950 15632
rect 22266 15620 22272 15632
rect 22227 15592 22272 15620
rect 22266 15580 22272 15592
rect 22324 15580 22330 15632
rect 22361 15623 22419 15629
rect 22361 15589 22373 15623
rect 22407 15620 22419 15623
rect 22450 15620 22456 15632
rect 22407 15592 22456 15620
rect 22407 15589 22419 15592
rect 22361 15583 22419 15589
rect 22450 15580 22456 15592
rect 22508 15580 22514 15632
rect 12882 15552 12888 15564
rect 12843 15524 12888 15552
rect 12882 15512 12888 15524
rect 12940 15512 12946 15564
rect 13066 15561 13072 15564
rect 13032 15555 13072 15561
rect 13032 15521 13044 15555
rect 13032 15515 13072 15521
rect 13066 15512 13072 15515
rect 13124 15512 13130 15564
rect 19046 15552 19052 15564
rect 19007 15524 19052 15552
rect 19046 15512 19052 15524
rect 19104 15512 19110 15564
rect 19138 15512 19144 15564
rect 19196 15552 19202 15564
rect 19233 15555 19291 15561
rect 19233 15552 19245 15555
rect 19196 15524 19245 15552
rect 19196 15512 19202 15524
rect 19233 15521 19245 15524
rect 19279 15521 19291 15555
rect 19233 15515 19291 15521
rect 21349 15555 21407 15561
rect 21349 15521 21361 15555
rect 21395 15552 21407 15555
rect 21714 15552 21720 15564
rect 21395 15524 21720 15552
rect 21395 15521 21407 15524
rect 21349 15515 21407 15521
rect 21714 15512 21720 15524
rect 21772 15512 21778 15564
rect 24385 15555 24443 15561
rect 24385 15521 24397 15555
rect 24431 15552 24443 15555
rect 24566 15552 24572 15564
rect 24431 15524 24572 15552
rect 24431 15521 24443 15524
rect 24385 15515 24443 15521
rect 24566 15512 24572 15524
rect 24624 15512 24630 15564
rect 12606 15444 12612 15496
rect 12664 15484 12670 15496
rect 13253 15487 13311 15493
rect 13253 15484 13265 15487
rect 12664 15456 13265 15484
rect 12664 15444 12670 15456
rect 13253 15453 13265 15456
rect 13299 15484 13311 15487
rect 13618 15484 13624 15496
rect 13299 15456 13624 15484
rect 13299 15453 13311 15456
rect 13253 15447 13311 15453
rect 13618 15444 13624 15456
rect 13676 15484 13682 15496
rect 14814 15484 14820 15496
rect 13676 15456 14820 15484
rect 13676 15444 13682 15456
rect 14814 15444 14820 15456
rect 14872 15444 14878 15496
rect 15277 15487 15335 15493
rect 15277 15453 15289 15487
rect 15323 15484 15335 15487
rect 15366 15484 15372 15496
rect 15323 15456 15372 15484
rect 15323 15453 15335 15456
rect 15277 15447 15335 15453
rect 15366 15444 15372 15456
rect 15424 15484 15430 15496
rect 16010 15484 16016 15496
rect 15424 15456 16016 15484
rect 15424 15444 15430 15456
rect 16010 15444 16016 15456
rect 16068 15444 16074 15496
rect 17114 15484 17120 15496
rect 17075 15456 17120 15484
rect 17114 15444 17120 15456
rect 17172 15444 17178 15496
rect 17393 15487 17451 15493
rect 17393 15453 17405 15487
rect 17439 15453 17451 15487
rect 17393 15447 17451 15453
rect 19509 15487 19567 15493
rect 19509 15453 19521 15487
rect 19555 15484 19567 15487
rect 20058 15484 20064 15496
rect 19555 15456 20064 15484
rect 19555 15453 19567 15456
rect 19509 15447 19567 15453
rect 11778 15376 11784 15428
rect 11836 15416 11842 15428
rect 12146 15416 12152 15428
rect 11836 15388 12152 15416
rect 11836 15376 11842 15388
rect 12146 15376 12152 15388
rect 12204 15416 12210 15428
rect 12204 15388 13204 15416
rect 12204 15376 12210 15388
rect 13176 15360 13204 15388
rect 16838 15376 16844 15428
rect 16896 15416 16902 15428
rect 17408 15416 17436 15447
rect 20058 15444 20064 15456
rect 20116 15484 20122 15496
rect 20429 15487 20487 15493
rect 20429 15484 20441 15487
rect 20116 15456 20441 15484
rect 20116 15444 20122 15456
rect 20429 15453 20441 15456
rect 20475 15453 20487 15487
rect 22542 15484 22548 15496
rect 22503 15456 22548 15484
rect 20429 15447 20487 15453
rect 22542 15444 22548 15456
rect 22600 15444 22606 15496
rect 24477 15487 24535 15493
rect 24477 15453 24489 15487
rect 24523 15484 24535 15487
rect 24842 15484 24848 15496
rect 24523 15456 24848 15484
rect 24523 15453 24535 15456
rect 24477 15447 24535 15453
rect 24842 15444 24848 15456
rect 24900 15444 24906 15496
rect 20242 15416 20248 15428
rect 16896 15388 17436 15416
rect 20203 15388 20248 15416
rect 16896 15376 16902 15388
rect 20242 15376 20248 15388
rect 20300 15376 20306 15428
rect 13158 15348 13164 15360
rect 13119 15320 13164 15348
rect 13158 15308 13164 15320
rect 13216 15308 13222 15360
rect 13526 15348 13532 15360
rect 13487 15320 13532 15348
rect 13526 15308 13532 15320
rect 13584 15308 13590 15360
rect 13710 15308 13716 15360
rect 13768 15348 13774 15360
rect 13897 15351 13955 15357
rect 13897 15348 13909 15351
rect 13768 15320 13909 15348
rect 13768 15308 13774 15320
rect 13897 15317 13909 15320
rect 13943 15317 13955 15351
rect 14998 15348 15004 15360
rect 14959 15320 15004 15348
rect 13897 15311 13955 15317
rect 14998 15308 15004 15320
rect 15056 15308 15062 15360
rect 632 15258 26392 15280
rect 632 15206 5176 15258
rect 5228 15206 5240 15258
rect 5292 15206 5304 15258
rect 5356 15206 5368 15258
rect 5420 15206 14510 15258
rect 14562 15206 14574 15258
rect 14626 15206 14638 15258
rect 14690 15206 14702 15258
rect 14754 15206 23843 15258
rect 23895 15206 23907 15258
rect 23959 15206 23971 15258
rect 24023 15206 24035 15258
rect 24087 15206 26392 15258
rect 632 15184 26392 15206
rect 12241 15147 12299 15153
rect 12241 15113 12253 15147
rect 12287 15144 12299 15147
rect 12514 15144 12520 15156
rect 12287 15116 12520 15144
rect 12287 15113 12299 15116
rect 12241 15107 12299 15113
rect 12514 15104 12520 15116
rect 12572 15144 12578 15156
rect 12882 15144 12888 15156
rect 12572 15116 12888 15144
rect 12572 15104 12578 15116
rect 12882 15104 12888 15116
rect 12940 15104 12946 15156
rect 12977 15147 13035 15153
rect 12977 15113 12989 15147
rect 13023 15144 13035 15147
rect 13158 15144 13164 15156
rect 13023 15116 13164 15144
rect 13023 15113 13035 15116
rect 12977 15107 13035 15113
rect 13158 15104 13164 15116
rect 13216 15104 13222 15156
rect 15645 15147 15703 15153
rect 15645 15113 15657 15147
rect 15691 15144 15703 15147
rect 15734 15144 15740 15156
rect 15691 15116 15740 15144
rect 15691 15113 15703 15116
rect 15645 15107 15703 15113
rect 15734 15104 15740 15116
rect 15792 15104 15798 15156
rect 16102 15104 16108 15156
rect 16160 15144 16166 15156
rect 16289 15147 16347 15153
rect 16289 15144 16301 15147
rect 16160 15116 16301 15144
rect 16160 15104 16166 15116
rect 16289 15113 16301 15116
rect 16335 15113 16347 15147
rect 17022 15144 17028 15156
rect 16983 15116 17028 15144
rect 16289 15107 16347 15113
rect 17022 15104 17028 15116
rect 17080 15104 17086 15156
rect 20058 15144 20064 15156
rect 20019 15116 20064 15144
rect 20058 15104 20064 15116
rect 20116 15104 20122 15156
rect 20521 15147 20579 15153
rect 20521 15113 20533 15147
rect 20567 15144 20579 15147
rect 20886 15144 20892 15156
rect 20567 15116 20892 15144
rect 20567 15113 20579 15116
rect 20521 15107 20579 15113
rect 20886 15104 20892 15116
rect 20944 15104 20950 15156
rect 22269 15147 22327 15153
rect 22269 15113 22281 15147
rect 22315 15144 22327 15147
rect 22450 15144 22456 15156
rect 22315 15116 22456 15144
rect 22315 15113 22327 15116
rect 22269 15107 22327 15113
rect 22450 15104 22456 15116
rect 22508 15104 22514 15156
rect 24934 15104 24940 15156
rect 24992 15144 24998 15156
rect 25213 15147 25271 15153
rect 25213 15144 25225 15147
rect 24992 15116 25225 15144
rect 24992 15104 24998 15116
rect 25213 15113 25225 15116
rect 25259 15113 25271 15147
rect 25213 15107 25271 15113
rect 12606 15076 12612 15088
rect 12567 15048 12612 15076
rect 12606 15036 12612 15048
rect 12664 15036 12670 15088
rect 13897 15011 13955 15017
rect 13897 14977 13909 15011
rect 13943 15008 13955 15011
rect 14725 15011 14783 15017
rect 14725 15008 14737 15011
rect 13943 14980 14737 15008
rect 13943 14977 13955 14980
rect 13897 14971 13955 14977
rect 14725 14977 14737 14980
rect 14771 15008 14783 15011
rect 14998 15008 15004 15020
rect 14771 14980 15004 15008
rect 14771 14977 14783 14980
rect 14725 14971 14783 14977
rect 14998 14968 15004 14980
rect 15056 14968 15062 15020
rect 19233 15011 19291 15017
rect 19233 14977 19245 15011
rect 19279 15008 19291 15011
rect 19506 15008 19512 15020
rect 19279 14980 19512 15008
rect 19279 14977 19291 14980
rect 19233 14971 19291 14977
rect 19506 14968 19512 14980
rect 19564 14968 19570 15020
rect 20334 14968 20340 15020
rect 20392 15008 20398 15020
rect 20797 15011 20855 15017
rect 20797 15008 20809 15011
rect 20392 14980 20809 15008
rect 20392 14968 20398 14980
rect 20797 14977 20809 14980
rect 20843 14977 20855 15011
rect 20797 14971 20855 14977
rect 22266 14968 22272 15020
rect 22324 15008 22330 15020
rect 22545 15011 22603 15017
rect 22545 15008 22557 15011
rect 22324 14980 22557 15008
rect 22324 14968 22330 14980
rect 22545 14977 22557 14980
rect 22591 14977 22603 15011
rect 22545 14971 22603 14977
rect 13434 14940 13440 14952
rect 13395 14912 13440 14940
rect 13434 14900 13440 14912
rect 13492 14900 13498 14952
rect 13710 14940 13716 14952
rect 13671 14912 13716 14940
rect 13710 14900 13716 14912
rect 13768 14900 13774 14952
rect 18586 14940 18592 14952
rect 18547 14912 18592 14940
rect 18586 14900 18592 14912
rect 18644 14900 18650 14952
rect 18957 14943 19015 14949
rect 18957 14909 18969 14943
rect 19003 14940 19015 14943
rect 19138 14940 19144 14952
rect 19003 14912 19144 14940
rect 19003 14909 19015 14912
rect 18957 14903 19015 14909
rect 13452 14872 13480 14900
rect 14173 14875 14231 14881
rect 14173 14872 14185 14875
rect 13452 14844 14185 14872
rect 14173 14841 14185 14844
rect 14219 14841 14231 14875
rect 14173 14835 14231 14841
rect 14633 14875 14691 14881
rect 14633 14841 14645 14875
rect 14679 14872 14691 14875
rect 15087 14875 15145 14881
rect 15087 14872 15099 14875
rect 14679 14844 15099 14872
rect 14679 14841 14691 14844
rect 14633 14835 14691 14841
rect 15087 14841 15099 14844
rect 15133 14872 15145 14875
rect 18972 14872 19000 14903
rect 19138 14900 19144 14912
rect 19196 14900 19202 14952
rect 23002 14940 23008 14952
rect 22915 14912 23008 14940
rect 23002 14900 23008 14912
rect 23060 14940 23066 14952
rect 23281 14943 23339 14949
rect 23281 14940 23293 14943
rect 23060 14912 23293 14940
rect 23060 14900 23066 14912
rect 23281 14909 23293 14912
rect 23327 14909 23339 14943
rect 23281 14903 23339 14909
rect 24820 14943 24878 14949
rect 24820 14909 24832 14943
rect 24866 14940 24878 14943
rect 24934 14940 24940 14952
rect 24866 14912 24940 14940
rect 24866 14909 24878 14912
rect 24820 14903 24878 14909
rect 24934 14900 24940 14912
rect 24992 14900 24998 14952
rect 15133 14844 15964 14872
rect 15133 14841 15145 14844
rect 15087 14835 15145 14841
rect 15936 14816 15964 14844
rect 18328 14844 19000 14872
rect 15918 14804 15924 14816
rect 15879 14776 15924 14804
rect 15918 14764 15924 14776
rect 15976 14764 15982 14816
rect 16473 14807 16531 14813
rect 16473 14773 16485 14807
rect 16519 14804 16531 14807
rect 16930 14804 16936 14816
rect 16519 14776 16936 14804
rect 16519 14773 16531 14776
rect 16473 14767 16531 14773
rect 16930 14764 16936 14776
rect 16988 14764 16994 14816
rect 17942 14804 17948 14816
rect 17903 14776 17948 14804
rect 17942 14764 17948 14776
rect 18000 14804 18006 14816
rect 18328 14813 18356 14844
rect 19966 14832 19972 14884
rect 20024 14872 20030 14884
rect 20242 14872 20248 14884
rect 20024 14844 20248 14872
rect 20024 14832 20030 14844
rect 20242 14832 20248 14844
rect 20300 14872 20306 14884
rect 20889 14875 20947 14881
rect 20889 14872 20901 14875
rect 20300 14844 20901 14872
rect 20300 14832 20306 14844
rect 20889 14841 20901 14844
rect 20935 14841 20947 14875
rect 20889 14835 20947 14841
rect 21441 14875 21499 14881
rect 21441 14841 21453 14875
rect 21487 14872 21499 14875
rect 21622 14872 21628 14884
rect 21487 14844 21628 14872
rect 21487 14841 21499 14844
rect 21441 14835 21499 14841
rect 18313 14807 18371 14813
rect 18313 14804 18325 14807
rect 18000 14776 18325 14804
rect 18000 14764 18006 14776
rect 18313 14773 18325 14776
rect 18359 14773 18371 14807
rect 18313 14767 18371 14773
rect 19046 14764 19052 14816
rect 19104 14804 19110 14816
rect 19509 14807 19567 14813
rect 19509 14804 19521 14807
rect 19104 14776 19521 14804
rect 19104 14764 19110 14776
rect 19509 14773 19521 14776
rect 19555 14773 19567 14807
rect 20904 14804 20932 14835
rect 21622 14832 21628 14844
rect 21680 14832 21686 14884
rect 23186 14872 23192 14884
rect 23147 14844 23192 14872
rect 23186 14832 23192 14844
rect 23244 14832 23250 14884
rect 24293 14875 24351 14881
rect 24293 14841 24305 14875
rect 24339 14872 24351 14875
rect 24566 14872 24572 14884
rect 24339 14844 24572 14872
rect 24339 14841 24351 14844
rect 24293 14835 24351 14841
rect 24566 14832 24572 14844
rect 24624 14832 24630 14884
rect 21717 14807 21775 14813
rect 21717 14804 21729 14807
rect 20904 14776 21729 14804
rect 19509 14767 19567 14773
rect 21717 14773 21729 14776
rect 21763 14773 21775 14807
rect 21717 14767 21775 14773
rect 24474 14764 24480 14816
rect 24532 14804 24538 14816
rect 24891 14807 24949 14813
rect 24891 14804 24903 14807
rect 24532 14776 24903 14804
rect 24532 14764 24538 14776
rect 24891 14773 24903 14776
rect 24937 14773 24949 14807
rect 24891 14767 24949 14773
rect 632 14714 26392 14736
rect 632 14662 9843 14714
rect 9895 14662 9907 14714
rect 9959 14662 9971 14714
rect 10023 14662 10035 14714
rect 10087 14662 19176 14714
rect 19228 14662 19240 14714
rect 19292 14662 19304 14714
rect 19356 14662 19368 14714
rect 19420 14662 26392 14714
rect 632 14640 26392 14662
rect 12977 14603 13035 14609
rect 12977 14569 12989 14603
rect 13023 14600 13035 14603
rect 13066 14600 13072 14612
rect 13023 14572 13072 14600
rect 13023 14569 13035 14572
rect 12977 14563 13035 14569
rect 13066 14560 13072 14572
rect 13124 14560 13130 14612
rect 16010 14560 16016 14612
rect 16068 14600 16074 14612
rect 16473 14603 16531 14609
rect 16473 14600 16485 14603
rect 16068 14572 16485 14600
rect 16068 14560 16074 14572
rect 16473 14569 16485 14572
rect 16519 14569 16531 14603
rect 17850 14600 17856 14612
rect 17811 14572 17856 14600
rect 16473 14563 16531 14569
rect 17850 14560 17856 14572
rect 17908 14560 17914 14612
rect 18586 14600 18592 14612
rect 18547 14572 18592 14600
rect 18586 14560 18592 14572
rect 18644 14560 18650 14612
rect 20245 14603 20303 14609
rect 20245 14569 20257 14603
rect 20291 14600 20303 14603
rect 20334 14600 20340 14612
rect 20291 14572 20340 14600
rect 20291 14569 20303 14572
rect 20245 14563 20303 14569
rect 20334 14560 20340 14572
rect 20392 14560 20398 14612
rect 21349 14603 21407 14609
rect 21349 14569 21361 14603
rect 21395 14600 21407 14603
rect 21438 14600 21444 14612
rect 21395 14572 21444 14600
rect 21395 14569 21407 14572
rect 21349 14563 21407 14569
rect 21438 14560 21444 14572
rect 21496 14600 21502 14612
rect 23002 14600 23008 14612
rect 21496 14572 23008 14600
rect 21496 14560 21502 14572
rect 23002 14560 23008 14572
rect 23060 14560 23066 14612
rect 9570 14492 9576 14544
rect 9628 14532 9634 14544
rect 9628 14504 9892 14532
rect 9628 14492 9634 14504
rect 9662 14464 9668 14476
rect 9623 14436 9668 14464
rect 9662 14424 9668 14436
rect 9720 14424 9726 14476
rect 9864 14473 9892 14504
rect 14906 14492 14912 14544
rect 14964 14532 14970 14544
rect 15001 14535 15059 14541
rect 15001 14532 15013 14535
rect 14964 14504 15013 14532
rect 14964 14492 14970 14504
rect 15001 14501 15013 14504
rect 15047 14501 15059 14535
rect 15001 14495 15059 14501
rect 15553 14535 15611 14541
rect 15553 14501 15565 14535
rect 15599 14532 15611 14535
rect 17114 14532 17120 14544
rect 15599 14504 17120 14532
rect 15599 14501 15611 14504
rect 15553 14495 15611 14501
rect 17114 14492 17120 14504
rect 17172 14532 17178 14544
rect 17485 14535 17543 14541
rect 17485 14532 17497 14535
rect 17172 14504 17497 14532
rect 17172 14492 17178 14504
rect 17485 14501 17497 14504
rect 17531 14501 17543 14535
rect 17485 14495 17543 14501
rect 20610 14492 20616 14544
rect 20668 14532 20674 14544
rect 20791 14535 20849 14541
rect 20791 14532 20803 14535
rect 20668 14504 20803 14532
rect 20668 14492 20674 14504
rect 20791 14501 20803 14504
rect 20837 14532 20849 14535
rect 20886 14532 20892 14544
rect 20837 14504 20892 14532
rect 20837 14501 20849 14504
rect 20791 14495 20849 14501
rect 20886 14492 20892 14504
rect 20944 14492 20950 14544
rect 21622 14492 21628 14544
rect 21680 14532 21686 14544
rect 22361 14535 22419 14541
rect 21680 14504 21725 14532
rect 21680 14492 21686 14504
rect 22361 14501 22373 14535
rect 22407 14532 22419 14535
rect 22634 14532 22640 14544
rect 22407 14504 22640 14532
rect 22407 14501 22419 14504
rect 22361 14495 22419 14501
rect 22634 14492 22640 14504
rect 22692 14532 22698 14544
rect 23186 14532 23192 14544
rect 22692 14504 23192 14532
rect 22692 14492 22698 14504
rect 23186 14492 23192 14504
rect 23244 14492 23250 14544
rect 9849 14467 9907 14473
rect 9849 14433 9861 14467
rect 9895 14433 9907 14467
rect 9849 14427 9907 14433
rect 11781 14467 11839 14473
rect 11781 14433 11793 14467
rect 11827 14464 11839 14467
rect 11870 14464 11876 14476
rect 11827 14436 11876 14464
rect 11827 14433 11839 14436
rect 11781 14427 11839 14433
rect 11870 14424 11876 14436
rect 11928 14424 11934 14476
rect 13434 14464 13440 14476
rect 13395 14436 13440 14464
rect 13434 14424 13440 14436
rect 13492 14424 13498 14476
rect 13713 14467 13771 14473
rect 13713 14433 13725 14467
rect 13759 14464 13771 14467
rect 13802 14464 13808 14476
rect 13759 14436 13808 14464
rect 13759 14433 13771 14436
rect 13713 14427 13771 14433
rect 13802 14424 13808 14436
rect 13860 14424 13866 14476
rect 16654 14464 16660 14476
rect 16615 14436 16660 14464
rect 16654 14424 16660 14436
rect 16712 14424 16718 14476
rect 16838 14464 16844 14476
rect 16799 14436 16844 14464
rect 16838 14424 16844 14436
rect 16896 14424 16902 14476
rect 19046 14464 19052 14476
rect 19007 14436 19052 14464
rect 19046 14424 19052 14436
rect 19104 14424 19110 14476
rect 19325 14467 19383 14473
rect 19325 14433 19337 14467
rect 19371 14464 19383 14467
rect 19690 14464 19696 14476
rect 19371 14436 19696 14464
rect 19371 14433 19383 14436
rect 19325 14427 19383 14433
rect 19690 14424 19696 14436
rect 19748 14424 19754 14476
rect 23646 14424 23652 14476
rect 23704 14464 23710 14476
rect 23833 14467 23891 14473
rect 23833 14464 23845 14467
rect 23704 14436 23845 14464
rect 23704 14424 23710 14436
rect 23833 14433 23845 14436
rect 23879 14433 23891 14467
rect 23833 14427 23891 14433
rect 13897 14399 13955 14405
rect 13897 14365 13909 14399
rect 13943 14396 13955 14399
rect 14354 14396 14360 14408
rect 13943 14368 14360 14396
rect 13943 14365 13955 14368
rect 13897 14359 13955 14365
rect 14354 14356 14360 14368
rect 14412 14356 14418 14408
rect 14906 14396 14912 14408
rect 14867 14368 14912 14396
rect 14906 14356 14912 14368
rect 14964 14356 14970 14408
rect 19509 14399 19567 14405
rect 19509 14365 19521 14399
rect 19555 14396 19567 14399
rect 20429 14399 20487 14405
rect 20429 14396 20441 14399
rect 19555 14368 20441 14396
rect 19555 14365 19567 14368
rect 19509 14359 19567 14365
rect 20429 14365 20441 14368
rect 20475 14396 20487 14399
rect 20886 14396 20892 14408
rect 20475 14368 20892 14396
rect 20475 14365 20487 14368
rect 20429 14359 20487 14365
rect 20886 14356 20892 14368
rect 20944 14356 20950 14408
rect 22266 14396 22272 14408
rect 22227 14368 22272 14396
rect 22266 14356 22272 14368
rect 22324 14356 22330 14408
rect 22910 14396 22916 14408
rect 22871 14368 22916 14396
rect 22910 14356 22916 14368
rect 22968 14356 22974 14408
rect 23002 14356 23008 14408
rect 23060 14396 23066 14408
rect 23741 14399 23799 14405
rect 23741 14396 23753 14399
rect 23060 14368 23753 14396
rect 23060 14356 23066 14368
rect 23741 14365 23753 14368
rect 23787 14365 23799 14399
rect 23741 14359 23799 14365
rect 9294 14220 9300 14272
rect 9352 14260 9358 14272
rect 9941 14263 9999 14269
rect 9941 14260 9953 14263
rect 9352 14232 9953 14260
rect 9352 14220 9358 14232
rect 9941 14229 9953 14232
rect 9987 14229 9999 14263
rect 9941 14223 9999 14229
rect 11965 14263 12023 14269
rect 11965 14229 11977 14263
rect 12011 14260 12023 14263
rect 12330 14260 12336 14272
rect 12011 14232 12336 14260
rect 12011 14229 12023 14232
rect 11965 14223 12023 14229
rect 12330 14220 12336 14232
rect 12388 14220 12394 14272
rect 19782 14260 19788 14272
rect 19743 14232 19788 14260
rect 19782 14220 19788 14232
rect 19840 14220 19846 14272
rect 23186 14260 23192 14272
rect 23147 14232 23192 14260
rect 23186 14220 23192 14232
rect 23244 14220 23250 14272
rect 632 14170 26392 14192
rect 632 14118 5176 14170
rect 5228 14118 5240 14170
rect 5292 14118 5304 14170
rect 5356 14118 5368 14170
rect 5420 14118 14510 14170
rect 14562 14118 14574 14170
rect 14626 14118 14638 14170
rect 14690 14118 14702 14170
rect 14754 14118 23843 14170
rect 23895 14118 23907 14170
rect 23959 14118 23971 14170
rect 24023 14118 24035 14170
rect 24087 14118 26392 14170
rect 632 14096 26392 14118
rect 8926 14056 8932 14068
rect 8887 14028 8932 14056
rect 8926 14016 8932 14028
rect 8984 14016 8990 14068
rect 9570 14016 9576 14068
rect 9628 14056 9634 14068
rect 10125 14059 10183 14065
rect 10125 14056 10137 14059
rect 9628 14028 10137 14056
rect 9628 14016 9634 14028
rect 10125 14025 10137 14028
rect 10171 14025 10183 14059
rect 10125 14019 10183 14025
rect 13710 14016 13716 14068
rect 13768 14056 13774 14068
rect 14081 14059 14139 14065
rect 14081 14056 14093 14059
rect 13768 14028 14093 14056
rect 13768 14016 13774 14028
rect 14081 14025 14093 14028
rect 14127 14025 14139 14059
rect 14081 14019 14139 14025
rect 11045 13991 11103 13997
rect 11045 13957 11057 13991
rect 11091 13988 11103 13991
rect 11778 13988 11784 14000
rect 11091 13960 11784 13988
rect 11091 13957 11103 13960
rect 11045 13951 11103 13957
rect 11778 13948 11784 13960
rect 11836 13948 11842 14000
rect 12425 13991 12483 13997
rect 12425 13988 12437 13991
rect 11980 13960 12437 13988
rect 9662 13880 9668 13932
rect 9720 13920 9726 13932
rect 9849 13923 9907 13929
rect 9849 13920 9861 13923
rect 9720 13892 9861 13920
rect 9720 13880 9726 13892
rect 9849 13889 9861 13892
rect 9895 13920 9907 13923
rect 10493 13923 10551 13929
rect 10493 13920 10505 13923
rect 9895 13892 10505 13920
rect 9895 13889 9907 13892
rect 9849 13883 9907 13889
rect 10493 13889 10505 13892
rect 10539 13889 10551 13923
rect 10493 13883 10551 13889
rect 8926 13812 8932 13864
rect 8984 13852 8990 13864
rect 9205 13855 9263 13861
rect 9205 13852 9217 13855
rect 8984 13824 9217 13852
rect 8984 13812 8990 13824
rect 9205 13821 9217 13824
rect 9251 13852 9263 13855
rect 9386 13852 9392 13864
rect 9251 13824 9392 13852
rect 9251 13821 9263 13824
rect 9205 13815 9263 13821
rect 9386 13812 9392 13824
rect 9444 13812 9450 13864
rect 10582 13812 10588 13864
rect 10640 13852 10646 13864
rect 10861 13855 10919 13861
rect 10861 13852 10873 13855
rect 10640 13824 10873 13852
rect 10640 13812 10646 13824
rect 10861 13821 10873 13824
rect 10907 13852 10919 13855
rect 11321 13855 11379 13861
rect 11321 13852 11333 13855
rect 10907 13824 11333 13852
rect 10907 13821 10919 13824
rect 10861 13815 10919 13821
rect 11321 13821 11333 13824
rect 11367 13821 11379 13855
rect 11980 13852 12008 13960
rect 12425 13957 12437 13960
rect 12471 13957 12483 13991
rect 12425 13951 12483 13957
rect 12241 13923 12299 13929
rect 12241 13889 12253 13923
rect 12287 13920 12299 13923
rect 13802 13920 13808 13932
rect 12287 13892 13112 13920
rect 13763 13892 13808 13920
rect 12287 13889 12299 13892
rect 12241 13883 12299 13889
rect 13084 13864 13112 13892
rect 13802 13880 13808 13892
rect 13860 13880 13866 13932
rect 14096 13920 14124 14019
rect 14998 14016 15004 14068
rect 15056 14056 15062 14068
rect 15645 14059 15703 14065
rect 15645 14056 15657 14059
rect 15056 14028 15657 14056
rect 15056 14016 15062 14028
rect 15645 14025 15657 14028
rect 15691 14025 15703 14059
rect 16378 14056 16384 14068
rect 16291 14028 16384 14056
rect 15645 14019 15703 14025
rect 16378 14016 16384 14028
rect 16436 14056 16442 14068
rect 16838 14056 16844 14068
rect 16436 14028 16844 14056
rect 16436 14016 16442 14028
rect 16838 14016 16844 14028
rect 16896 14016 16902 14068
rect 17390 14056 17396 14068
rect 17351 14028 17396 14056
rect 17390 14016 17396 14028
rect 17448 14016 17454 14068
rect 18865 14059 18923 14065
rect 18865 14025 18877 14059
rect 18911 14056 18923 14059
rect 19046 14056 19052 14068
rect 18911 14028 19052 14056
rect 18911 14025 18923 14028
rect 18865 14019 18923 14025
rect 14541 13991 14599 13997
rect 14541 13957 14553 13991
rect 14587 13988 14599 13991
rect 14814 13988 14820 14000
rect 14587 13960 14820 13988
rect 14587 13957 14599 13960
rect 14541 13951 14599 13957
rect 14814 13948 14820 13960
rect 14872 13988 14878 14000
rect 16654 13988 16660 14000
rect 14872 13960 16660 13988
rect 14872 13948 14878 13960
rect 16654 13948 16660 13960
rect 16712 13988 16718 14000
rect 17025 13991 17083 13997
rect 17025 13988 17037 13991
rect 16712 13960 17037 13988
rect 16712 13948 16718 13960
rect 17025 13957 17037 13960
rect 17071 13988 17083 13991
rect 18880 13988 18908 14019
rect 19046 14016 19052 14028
rect 19104 14016 19110 14068
rect 20242 14056 20248 14068
rect 20203 14028 20248 14056
rect 20242 14016 20248 14028
rect 20300 14016 20306 14068
rect 20610 14056 20616 14068
rect 20571 14028 20616 14056
rect 20610 14016 20616 14028
rect 20668 14016 20674 14068
rect 20886 14056 20892 14068
rect 20847 14028 20892 14056
rect 20886 14016 20892 14028
rect 20944 14016 20950 14068
rect 21438 14056 21444 14068
rect 21399 14028 21444 14056
rect 21438 14016 21444 14028
rect 21496 14016 21502 14068
rect 22634 14056 22640 14068
rect 22595 14028 22640 14056
rect 22634 14016 22640 14028
rect 22692 14016 22698 14068
rect 22910 14016 22916 14068
rect 22968 14016 22974 14068
rect 23646 14016 23652 14068
rect 23704 14056 23710 14068
rect 24201 14059 24259 14065
rect 24201 14056 24213 14059
rect 23704 14028 24213 14056
rect 23704 14016 23710 14028
rect 24201 14025 24213 14028
rect 24247 14025 24259 14059
rect 24201 14019 24259 14025
rect 17071 13960 18908 13988
rect 19233 13991 19291 13997
rect 17071 13957 17083 13960
rect 17025 13951 17083 13957
rect 19233 13957 19245 13991
rect 19279 13988 19291 13991
rect 20628 13988 20656 14016
rect 19279 13960 20656 13988
rect 22177 13991 22235 13997
rect 19279 13957 19291 13960
rect 19233 13951 19291 13957
rect 14262 13920 14268 13932
rect 14096 13892 14268 13920
rect 14262 13880 14268 13892
rect 14320 13920 14326 13932
rect 17942 13920 17948 13932
rect 14320 13892 15136 13920
rect 17903 13892 17948 13920
rect 14320 13880 14326 13892
rect 12514 13852 12520 13864
rect 11321 13815 11379 13821
rect 11428 13824 12008 13852
rect 12475 13824 12520 13852
rect 11428 13796 11456 13824
rect 12514 13812 12520 13824
rect 12572 13812 12578 13864
rect 13066 13852 13072 13864
rect 13027 13824 13072 13852
rect 13066 13812 13072 13824
rect 13124 13812 13130 13864
rect 13434 13852 13440 13864
rect 13395 13824 13440 13852
rect 13434 13812 13440 13824
rect 13492 13812 13498 13864
rect 14814 13852 14820 13864
rect 14775 13824 14820 13852
rect 14814 13812 14820 13824
rect 14872 13812 14878 13864
rect 15108 13861 15136 13892
rect 17942 13880 17948 13892
rect 18000 13880 18006 13932
rect 19325 13923 19383 13929
rect 19325 13889 19337 13923
rect 19371 13920 19383 13923
rect 19782 13920 19788 13932
rect 19371 13892 19788 13920
rect 19371 13889 19383 13892
rect 19325 13883 19383 13889
rect 19782 13880 19788 13892
rect 19840 13880 19846 13932
rect 15093 13855 15151 13861
rect 15093 13821 15105 13855
rect 15139 13821 15151 13855
rect 15093 13815 15151 13821
rect 11410 13744 11416 13796
rect 11468 13744 11474 13796
rect 15366 13784 15372 13796
rect 15327 13756 15372 13784
rect 15366 13744 15372 13756
rect 15424 13744 15430 13796
rect 17666 13784 17672 13796
rect 17627 13756 17672 13784
rect 17666 13744 17672 13756
rect 17724 13744 17730 13796
rect 17761 13787 17819 13793
rect 17761 13753 17773 13787
rect 17807 13753 17819 13787
rect 17761 13747 17819 13753
rect 19687 13787 19745 13793
rect 19687 13753 19699 13787
rect 19733 13784 19745 13787
rect 19886 13784 19914 13960
rect 22177 13957 22189 13991
rect 22223 13988 22235 13991
rect 22928 13988 22956 14016
rect 22223 13960 22956 13988
rect 24937 13991 24995 13997
rect 22223 13957 22235 13960
rect 22177 13951 22235 13957
rect 24937 13957 24949 13991
rect 24983 13988 24995 13991
rect 25302 13988 25308 14000
rect 24983 13960 25308 13988
rect 24983 13957 24995 13960
rect 24937 13951 24995 13957
rect 25302 13948 25308 13960
rect 25360 13948 25366 14000
rect 21162 13880 21168 13932
rect 21220 13920 21226 13932
rect 21622 13920 21628 13932
rect 21220 13892 21628 13920
rect 21220 13880 21226 13892
rect 21622 13880 21628 13892
rect 21680 13920 21686 13932
rect 21680 13892 21773 13920
rect 21680 13880 21686 13892
rect 21438 13812 21444 13864
rect 21496 13812 21502 13864
rect 23002 13852 23008 13864
rect 22963 13824 23008 13852
rect 23002 13812 23008 13824
rect 23060 13852 23066 13864
rect 23189 13855 23247 13861
rect 23189 13852 23201 13855
rect 23060 13824 23201 13852
rect 23060 13812 23066 13824
rect 23189 13821 23201 13824
rect 23235 13821 23247 13855
rect 23189 13815 23247 13821
rect 23278 13812 23284 13864
rect 23336 13852 23342 13864
rect 23741 13855 23799 13861
rect 23741 13852 23753 13855
rect 23336 13824 23753 13852
rect 23336 13812 23342 13824
rect 23741 13821 23753 13824
rect 23787 13852 23799 13855
rect 24014 13852 24020 13864
rect 23787 13824 24020 13852
rect 23787 13821 23799 13824
rect 23741 13815 23799 13821
rect 24014 13812 24020 13824
rect 24072 13812 24078 13864
rect 24382 13812 24388 13864
rect 24440 13852 24446 13864
rect 24753 13855 24811 13861
rect 24753 13852 24765 13855
rect 24440 13824 24765 13852
rect 24440 13812 24446 13824
rect 24753 13821 24765 13824
rect 24799 13852 24811 13855
rect 25305 13855 25363 13861
rect 25305 13852 25317 13855
rect 24799 13824 25317 13852
rect 24799 13821 24811 13824
rect 24753 13815 24811 13821
rect 25305 13821 25317 13824
rect 25351 13821 25363 13855
rect 25305 13815 25363 13821
rect 19733 13756 19914 13784
rect 21456 13784 21484 13812
rect 21717 13787 21775 13793
rect 21717 13784 21729 13787
rect 21456 13756 21729 13784
rect 19733 13753 19745 13756
rect 19687 13747 19745 13753
rect 21717 13753 21729 13756
rect 21763 13753 21775 13787
rect 21717 13747 21775 13753
rect 10674 13676 10680 13728
rect 10732 13716 10738 13728
rect 11689 13719 11747 13725
rect 11689 13716 11701 13719
rect 10732 13688 11701 13716
rect 10732 13676 10738 13688
rect 11689 13685 11701 13688
rect 11735 13716 11747 13719
rect 11870 13716 11876 13728
rect 11735 13688 11876 13716
rect 11735 13685 11747 13688
rect 11689 13679 11747 13685
rect 11870 13676 11876 13688
rect 11928 13676 11934 13728
rect 16470 13716 16476 13728
rect 16431 13688 16476 13716
rect 16470 13676 16476 13688
rect 16528 13676 16534 13728
rect 17390 13676 17396 13728
rect 17448 13716 17454 13728
rect 17776 13716 17804 13747
rect 17448 13688 17804 13716
rect 17448 13676 17454 13688
rect 23186 13676 23192 13728
rect 23244 13716 23250 13728
rect 23281 13719 23339 13725
rect 23281 13716 23293 13719
rect 23244 13688 23293 13716
rect 23244 13676 23250 13688
rect 23281 13685 23293 13688
rect 23327 13685 23339 13719
rect 23281 13679 23339 13685
rect 632 13626 26392 13648
rect 632 13574 9843 13626
rect 9895 13574 9907 13626
rect 9959 13574 9971 13626
rect 10023 13574 10035 13626
rect 10087 13574 19176 13626
rect 19228 13574 19240 13626
rect 19292 13574 19304 13626
rect 19356 13574 19368 13626
rect 19420 13574 26392 13626
rect 632 13552 26392 13574
rect 12425 13515 12483 13521
rect 12425 13481 12437 13515
rect 12471 13512 12483 13515
rect 12514 13512 12520 13524
rect 12471 13484 12520 13512
rect 12471 13481 12483 13484
rect 12425 13475 12483 13481
rect 12514 13472 12520 13484
rect 12572 13512 12578 13524
rect 12572 13484 12836 13512
rect 12572 13472 12578 13484
rect 12808 13453 12836 13484
rect 14906 13472 14912 13524
rect 14964 13512 14970 13524
rect 15001 13515 15059 13521
rect 15001 13512 15013 13515
rect 14964 13484 15013 13512
rect 14964 13472 14970 13484
rect 15001 13481 15013 13484
rect 15047 13512 15059 13515
rect 15090 13512 15096 13524
rect 15047 13484 15096 13512
rect 15047 13481 15059 13484
rect 15001 13475 15059 13481
rect 15090 13472 15096 13484
rect 15148 13472 15154 13524
rect 15461 13515 15519 13521
rect 15461 13481 15473 13515
rect 15507 13512 15519 13515
rect 16010 13512 16016 13524
rect 15507 13484 16016 13512
rect 15507 13481 15519 13484
rect 15461 13475 15519 13481
rect 16010 13472 16016 13484
rect 16068 13472 16074 13524
rect 16473 13515 16531 13521
rect 16473 13481 16485 13515
rect 16519 13512 16531 13515
rect 17298 13512 17304 13524
rect 16519 13484 17304 13512
rect 16519 13481 16531 13484
rect 16473 13475 16531 13481
rect 17298 13472 17304 13484
rect 17356 13472 17362 13524
rect 17942 13512 17948 13524
rect 17408 13484 17948 13512
rect 15918 13453 15924 13456
rect 12793 13447 12851 13453
rect 12793 13413 12805 13447
rect 12839 13413 12851 13447
rect 15915 13444 15924 13453
rect 15831 13416 15924 13444
rect 12793 13407 12851 13413
rect 15915 13407 15924 13416
rect 15976 13444 15982 13456
rect 16286 13444 16292 13456
rect 15976 13416 16292 13444
rect 15918 13404 15924 13407
rect 15976 13404 15982 13416
rect 16286 13404 16292 13416
rect 16344 13404 16350 13456
rect 17022 13404 17028 13456
rect 17080 13444 17086 13456
rect 17408 13453 17436 13484
rect 17942 13472 17948 13484
rect 18000 13472 18006 13524
rect 18862 13472 18868 13524
rect 18920 13512 18926 13524
rect 19141 13515 19199 13521
rect 19141 13512 19153 13515
rect 18920 13484 19153 13512
rect 18920 13472 18926 13484
rect 19141 13481 19153 13484
rect 19187 13481 19199 13515
rect 22266 13512 22272 13524
rect 22227 13484 22272 13512
rect 19141 13475 19199 13481
rect 22266 13472 22272 13484
rect 22324 13472 22330 13524
rect 23278 13472 23284 13524
rect 23336 13512 23342 13524
rect 23465 13515 23523 13521
rect 23465 13512 23477 13515
rect 23336 13484 23477 13512
rect 23336 13472 23342 13484
rect 23465 13481 23477 13484
rect 23511 13512 23523 13515
rect 24290 13512 24296 13524
rect 23511 13484 24296 13512
rect 23511 13481 23523 13484
rect 23465 13475 23523 13481
rect 24290 13472 24296 13484
rect 24348 13472 24354 13524
rect 17209 13447 17267 13453
rect 17209 13444 17221 13447
rect 17080 13416 17221 13444
rect 17080 13404 17086 13416
rect 17209 13413 17221 13416
rect 17255 13444 17267 13447
rect 17393 13447 17451 13453
rect 17393 13444 17405 13447
rect 17255 13416 17405 13444
rect 17255 13413 17267 13416
rect 17209 13407 17267 13413
rect 17393 13413 17405 13416
rect 17439 13413 17451 13447
rect 17393 13407 17451 13413
rect 17485 13447 17543 13453
rect 17485 13413 17497 13447
rect 17531 13444 17543 13447
rect 17574 13444 17580 13456
rect 17531 13416 17580 13444
rect 17531 13413 17543 13416
rect 17485 13407 17543 13413
rect 17574 13404 17580 13416
rect 17632 13404 17638 13456
rect 19598 13444 19604 13456
rect 18880 13416 19604 13444
rect 9386 13376 9392 13388
rect 9347 13348 9392 13376
rect 9386 13336 9392 13348
rect 9444 13336 9450 13388
rect 9570 13336 9576 13388
rect 9628 13376 9634 13388
rect 9941 13379 9999 13385
rect 9941 13376 9953 13379
rect 9628 13348 9953 13376
rect 9628 13336 9634 13348
rect 9941 13345 9953 13348
rect 9987 13345 9999 13379
rect 11870 13376 11876 13388
rect 11831 13348 11876 13376
rect 9941 13339 9999 13345
rect 11870 13336 11876 13348
rect 11928 13336 11934 13388
rect 13066 13376 13072 13388
rect 13027 13348 13072 13376
rect 13066 13336 13072 13348
rect 13124 13336 13130 13388
rect 14354 13336 14360 13388
rect 14412 13376 14418 13388
rect 15553 13379 15611 13385
rect 15553 13376 15565 13379
rect 14412 13348 15565 13376
rect 14412 13336 14418 13348
rect 15553 13345 15565 13348
rect 15599 13376 15611 13379
rect 16102 13376 16108 13388
rect 15599 13348 16108 13376
rect 15599 13345 15611 13348
rect 15553 13339 15611 13345
rect 16102 13336 16108 13348
rect 16160 13336 16166 13388
rect 18880 13385 18908 13416
rect 19598 13404 19604 13416
rect 19656 13404 19662 13456
rect 20150 13404 20156 13456
rect 20208 13444 20214 13456
rect 20613 13447 20671 13453
rect 20613 13444 20625 13447
rect 20208 13416 20625 13444
rect 20208 13404 20214 13416
rect 20613 13413 20625 13416
rect 20659 13413 20671 13447
rect 21162 13444 21168 13456
rect 21123 13416 21168 13444
rect 20613 13407 20671 13413
rect 21162 13404 21168 13416
rect 21220 13404 21226 13456
rect 22450 13404 22456 13456
rect 22508 13444 22514 13456
rect 22545 13447 22603 13453
rect 22545 13444 22557 13447
rect 22508 13416 22557 13444
rect 22508 13404 22514 13416
rect 22545 13413 22557 13416
rect 22591 13444 22603 13447
rect 22910 13444 22916 13456
rect 22591 13416 22916 13444
rect 22591 13413 22603 13416
rect 22545 13407 22603 13413
rect 22910 13404 22916 13416
rect 22968 13404 22974 13456
rect 18865 13379 18923 13385
rect 18865 13345 18877 13379
rect 18911 13345 18923 13379
rect 18865 13339 18923 13345
rect 18954 13336 18960 13388
rect 19012 13376 19018 13388
rect 19049 13379 19107 13385
rect 19049 13376 19061 13379
rect 19012 13348 19061 13376
rect 19012 13336 19018 13348
rect 19049 13345 19061 13348
rect 19095 13345 19107 13379
rect 24198 13376 24204 13388
rect 24159 13348 24204 13376
rect 19049 13339 19107 13345
rect 24198 13336 24204 13348
rect 24256 13336 24262 13388
rect 11778 13268 11784 13320
rect 11836 13308 11842 13320
rect 14078 13308 14084 13320
rect 11836 13280 14084 13308
rect 11836 13268 11842 13280
rect 14078 13268 14084 13280
rect 14136 13308 14142 13320
rect 14173 13311 14231 13317
rect 14173 13308 14185 13311
rect 14136 13280 14185 13308
rect 14136 13268 14142 13280
rect 14173 13277 14185 13280
rect 14219 13277 14231 13311
rect 14173 13271 14231 13277
rect 20334 13268 20340 13320
rect 20392 13308 20398 13320
rect 20521 13311 20579 13317
rect 20521 13308 20533 13311
rect 20392 13280 20533 13308
rect 20392 13268 20398 13280
rect 20521 13277 20533 13280
rect 20567 13277 20579 13311
rect 20521 13271 20579 13277
rect 22453 13311 22511 13317
rect 22453 13277 22465 13311
rect 22499 13308 22511 13311
rect 22542 13308 22548 13320
rect 22499 13280 22548 13308
rect 22499 13277 22511 13280
rect 22453 13271 22511 13277
rect 22542 13268 22548 13280
rect 22600 13268 22606 13320
rect 23094 13308 23100 13320
rect 23055 13280 23100 13308
rect 23094 13268 23100 13280
rect 23152 13268 23158 13320
rect 23738 13268 23744 13320
rect 23796 13308 23802 13320
rect 23925 13311 23983 13317
rect 23925 13308 23937 13311
rect 23796 13280 23937 13308
rect 23796 13268 23802 13280
rect 23925 13277 23937 13280
rect 23971 13277 23983 13311
rect 23925 13271 23983 13277
rect 17942 13240 17948 13252
rect 17903 13212 17948 13240
rect 17942 13200 17948 13212
rect 18000 13200 18006 13252
rect 18773 13243 18831 13249
rect 18773 13209 18785 13243
rect 18819 13240 18831 13243
rect 18819 13212 19736 13240
rect 18819 13209 18831 13212
rect 18773 13203 18831 13209
rect 19708 13184 19736 13212
rect 9202 13132 9208 13184
rect 9260 13172 9266 13184
rect 9481 13175 9539 13181
rect 9481 13172 9493 13175
rect 9260 13144 9493 13172
rect 9260 13132 9266 13144
rect 9481 13141 9493 13144
rect 9527 13141 9539 13175
rect 10490 13172 10496 13184
rect 10451 13144 10496 13172
rect 9481 13135 9539 13141
rect 10490 13132 10496 13144
rect 10548 13132 10554 13184
rect 10674 13132 10680 13184
rect 10732 13172 10738 13184
rect 10769 13175 10827 13181
rect 10769 13172 10781 13175
rect 10732 13144 10781 13172
rect 10732 13132 10738 13144
rect 10769 13141 10781 13144
rect 10815 13141 10827 13175
rect 11686 13172 11692 13184
rect 11647 13144 11692 13172
rect 10769 13135 10827 13141
rect 11686 13132 11692 13144
rect 11744 13132 11750 13184
rect 11778 13132 11784 13184
rect 11836 13172 11842 13184
rect 13802 13172 13808 13184
rect 11836 13144 13808 13172
rect 11836 13132 11842 13144
rect 13802 13132 13808 13144
rect 13860 13132 13866 13184
rect 19690 13172 19696 13184
rect 19651 13144 19696 13172
rect 19690 13132 19696 13144
rect 19748 13132 19754 13184
rect 21070 13132 21076 13184
rect 21128 13172 21134 13184
rect 21441 13175 21499 13181
rect 21441 13172 21453 13175
rect 21128 13144 21453 13172
rect 21128 13132 21134 13144
rect 21441 13141 21453 13144
rect 21487 13141 21499 13175
rect 21441 13135 21499 13141
rect 632 13082 26392 13104
rect 632 13030 5176 13082
rect 5228 13030 5240 13082
rect 5292 13030 5304 13082
rect 5356 13030 5368 13082
rect 5420 13030 14510 13082
rect 14562 13030 14574 13082
rect 14626 13030 14638 13082
rect 14690 13030 14702 13082
rect 14754 13030 23843 13082
rect 23895 13030 23907 13082
rect 23959 13030 23971 13082
rect 24023 13030 24035 13082
rect 24087 13030 26392 13082
rect 632 13008 26392 13030
rect 9205 12971 9263 12977
rect 9205 12937 9217 12971
rect 9251 12968 9263 12971
rect 9294 12968 9300 12980
rect 9251 12940 9300 12968
rect 9251 12937 9263 12940
rect 9205 12931 9263 12937
rect 9294 12928 9300 12940
rect 9352 12928 9358 12980
rect 9386 12928 9392 12980
rect 9444 12968 9450 12980
rect 10125 12971 10183 12977
rect 10125 12968 10137 12971
rect 9444 12940 10137 12968
rect 9444 12928 9450 12940
rect 10125 12937 10137 12940
rect 10171 12937 10183 12971
rect 10582 12968 10588 12980
rect 10543 12940 10588 12968
rect 10125 12931 10183 12937
rect 10582 12928 10588 12940
rect 10640 12928 10646 12980
rect 11410 12968 11416 12980
rect 11323 12940 11416 12968
rect 9478 12900 9484 12912
rect 9439 12872 9484 12900
rect 9478 12860 9484 12872
rect 9536 12860 9542 12912
rect 9570 12860 9576 12912
rect 9628 12900 9634 12912
rect 9757 12903 9815 12909
rect 9757 12900 9769 12903
rect 9628 12872 9769 12900
rect 9628 12860 9634 12872
rect 9757 12869 9769 12872
rect 9803 12869 9815 12903
rect 9757 12863 9815 12869
rect 10214 12860 10220 12912
rect 10272 12900 10278 12912
rect 11336 12909 11364 12940
rect 11410 12928 11416 12940
rect 11468 12968 11474 12980
rect 12054 12968 12060 12980
rect 11468 12940 12060 12968
rect 11468 12928 11474 12940
rect 12054 12928 12060 12940
rect 12112 12928 12118 12980
rect 13618 12968 13624 12980
rect 13579 12940 13624 12968
rect 13618 12928 13624 12940
rect 13676 12928 13682 12980
rect 14078 12968 14084 12980
rect 14039 12940 14084 12968
rect 14078 12928 14084 12940
rect 14136 12928 14142 12980
rect 14262 12968 14268 12980
rect 14223 12940 14268 12968
rect 14262 12928 14268 12940
rect 14320 12928 14326 12980
rect 16930 12968 16936 12980
rect 16891 12940 16936 12968
rect 16930 12928 16936 12940
rect 16988 12928 16994 12980
rect 18954 12968 18960 12980
rect 18915 12940 18960 12968
rect 18954 12928 18960 12940
rect 19012 12928 19018 12980
rect 20150 12928 20156 12980
rect 20208 12968 20214 12980
rect 20429 12971 20487 12977
rect 20429 12968 20441 12971
rect 20208 12940 20441 12968
rect 20208 12928 20214 12940
rect 20429 12937 20441 12940
rect 20475 12937 20487 12971
rect 22450 12968 22456 12980
rect 22411 12940 22456 12968
rect 20429 12931 20487 12937
rect 22450 12928 22456 12940
rect 22508 12928 22514 12980
rect 24198 12968 24204 12980
rect 24159 12940 24204 12968
rect 24198 12928 24204 12940
rect 24256 12928 24262 12980
rect 10447 12903 10505 12909
rect 10447 12900 10459 12903
rect 10272 12872 10459 12900
rect 10272 12860 10278 12872
rect 10447 12869 10459 12872
rect 10493 12900 10505 12903
rect 11321 12903 11379 12909
rect 11321 12900 11333 12903
rect 10493 12872 11333 12900
rect 10493 12869 10505 12872
rect 10447 12863 10505 12869
rect 11321 12869 11333 12872
rect 11367 12869 11379 12903
rect 11321 12863 11379 12869
rect 11597 12903 11655 12909
rect 11597 12869 11609 12903
rect 11643 12900 11655 12903
rect 12146 12900 12152 12912
rect 11643 12872 12152 12900
rect 11643 12869 11655 12872
rect 11597 12863 11655 12869
rect 12146 12860 12152 12872
rect 12204 12860 12210 12912
rect 13636 12900 13664 12928
rect 13636 12872 14216 12900
rect 10674 12832 10680 12844
rect 10635 12804 10680 12832
rect 10674 12792 10680 12804
rect 10732 12792 10738 12844
rect 9294 12764 9300 12776
rect 9255 12736 9300 12764
rect 9294 12724 9300 12736
rect 9352 12724 9358 12776
rect 12164 12773 12192 12860
rect 14188 12841 14216 12872
rect 13952 12835 14010 12841
rect 13952 12832 13964 12835
rect 13636 12804 13964 12832
rect 12149 12767 12207 12773
rect 12149 12733 12161 12767
rect 12195 12733 12207 12767
rect 12149 12727 12207 12733
rect 9202 12656 9208 12708
rect 9260 12696 9266 12708
rect 10309 12699 10367 12705
rect 10309 12696 10321 12699
rect 9260 12668 10321 12696
rect 9260 12656 9266 12668
rect 10309 12665 10321 12668
rect 10355 12696 10367 12699
rect 10490 12696 10496 12708
rect 10355 12668 10496 12696
rect 10355 12665 10367 12668
rect 10309 12659 10367 12665
rect 10490 12656 10496 12668
rect 10548 12656 10554 12708
rect 13342 12656 13348 12708
rect 13400 12696 13406 12708
rect 13636 12696 13664 12804
rect 13952 12801 13964 12804
rect 13998 12801 14010 12835
rect 13952 12795 14010 12801
rect 14173 12835 14231 12841
rect 14173 12801 14185 12835
rect 14219 12801 14231 12835
rect 14173 12795 14231 12801
rect 15737 12835 15795 12841
rect 15737 12801 15749 12835
rect 15783 12832 15795 12835
rect 16010 12832 16016 12844
rect 15783 12804 16016 12832
rect 15783 12801 15795 12804
rect 15737 12795 15795 12801
rect 16010 12792 16016 12804
rect 16068 12792 16074 12844
rect 16948 12832 16976 12928
rect 17298 12900 17304 12912
rect 17259 12872 17304 12900
rect 17298 12860 17304 12872
rect 17356 12860 17362 12912
rect 20702 12860 20708 12912
rect 20760 12900 20766 12912
rect 20981 12903 21039 12909
rect 20981 12900 20993 12903
rect 20760 12872 20993 12900
rect 20760 12860 20766 12872
rect 20981 12869 20993 12872
rect 21027 12869 21039 12903
rect 20981 12863 21039 12869
rect 17669 12835 17727 12841
rect 17669 12832 17681 12835
rect 16948 12804 17681 12832
rect 17669 12801 17681 12804
rect 17715 12801 17727 12835
rect 17942 12832 17948 12844
rect 17903 12804 17948 12832
rect 17669 12795 17727 12801
rect 17942 12792 17948 12804
rect 18000 12792 18006 12844
rect 19782 12832 19788 12844
rect 19743 12804 19788 12832
rect 19782 12792 19788 12804
rect 19840 12792 19846 12844
rect 20242 12792 20248 12844
rect 20300 12832 20306 12844
rect 21070 12832 21076 12844
rect 20300 12804 21076 12832
rect 20300 12792 20306 12804
rect 21070 12792 21076 12804
rect 21128 12792 21134 12844
rect 23094 12792 23100 12844
rect 23152 12832 23158 12844
rect 23557 12835 23615 12841
rect 23557 12832 23569 12835
rect 23152 12804 23569 12832
rect 23152 12792 23158 12804
rect 23557 12801 23569 12804
rect 23603 12801 23615 12835
rect 23557 12795 23615 12801
rect 13802 12764 13808 12776
rect 13763 12736 13808 12764
rect 13802 12724 13808 12736
rect 13860 12764 13866 12776
rect 14354 12764 14360 12776
rect 13860 12736 14360 12764
rect 13860 12724 13866 12736
rect 14354 12724 14360 12736
rect 14412 12724 14418 12776
rect 18494 12724 18500 12776
rect 18552 12764 18558 12776
rect 19141 12767 19199 12773
rect 19141 12764 19153 12767
rect 18552 12736 19153 12764
rect 18552 12724 18558 12736
rect 19141 12733 19153 12736
rect 19187 12764 19199 12767
rect 19506 12764 19512 12776
rect 19187 12736 19512 12764
rect 19187 12733 19199 12736
rect 19141 12727 19199 12733
rect 19506 12724 19512 12736
rect 19564 12724 19570 12776
rect 19690 12764 19696 12776
rect 19651 12736 19696 12764
rect 19690 12724 19696 12736
rect 19748 12724 19754 12776
rect 20886 12773 20892 12776
rect 20852 12767 20892 12773
rect 20852 12733 20864 12767
rect 20852 12727 20892 12733
rect 20886 12724 20892 12727
rect 20944 12724 20950 12776
rect 21438 12764 21444 12776
rect 21399 12736 21444 12764
rect 21438 12724 21444 12736
rect 21496 12724 21502 12776
rect 22634 12724 22640 12776
rect 22692 12764 22698 12776
rect 23002 12764 23008 12776
rect 22692 12736 23008 12764
rect 22692 12724 22698 12736
rect 23002 12724 23008 12736
rect 23060 12724 23066 12776
rect 24753 12767 24811 12773
rect 24753 12733 24765 12767
rect 24799 12764 24811 12767
rect 25026 12764 25032 12776
rect 24799 12736 25032 12764
rect 24799 12733 24811 12736
rect 24753 12727 24811 12733
rect 25026 12724 25032 12736
rect 25084 12764 25090 12776
rect 25305 12767 25363 12773
rect 25305 12764 25317 12767
rect 25084 12736 25317 12764
rect 25084 12724 25090 12736
rect 25305 12733 25317 12736
rect 25351 12733 25363 12767
rect 25305 12727 25363 12733
rect 14817 12699 14875 12705
rect 14817 12696 14829 12699
rect 13400 12668 14829 12696
rect 13400 12656 13406 12668
rect 14817 12665 14829 12668
rect 14863 12696 14875 12699
rect 14906 12696 14912 12708
rect 14863 12668 14912 12696
rect 14863 12665 14875 12668
rect 14817 12659 14875 12665
rect 14906 12656 14912 12668
rect 14964 12656 14970 12708
rect 15277 12699 15335 12705
rect 15277 12665 15289 12699
rect 15323 12696 15335 12699
rect 15645 12699 15703 12705
rect 15645 12696 15657 12699
rect 15323 12668 15657 12696
rect 15323 12665 15335 12668
rect 15277 12659 15335 12665
rect 15645 12665 15657 12668
rect 15691 12696 15703 12699
rect 16099 12699 16157 12705
rect 16099 12696 16111 12699
rect 15691 12668 16111 12696
rect 15691 12665 15703 12668
rect 15645 12659 15703 12665
rect 16099 12665 16111 12668
rect 16145 12696 16157 12699
rect 16286 12696 16292 12708
rect 16145 12668 16292 12696
rect 16145 12665 16157 12668
rect 16099 12659 16157 12665
rect 16286 12656 16292 12668
rect 16344 12656 16350 12708
rect 17298 12656 17304 12708
rect 17356 12696 17362 12708
rect 17761 12699 17819 12705
rect 17761 12696 17773 12699
rect 17356 12668 17773 12696
rect 17356 12656 17362 12668
rect 17761 12665 17773 12668
rect 17807 12665 17819 12699
rect 17761 12659 17819 12665
rect 20426 12656 20432 12708
rect 20484 12696 20490 12708
rect 20705 12699 20763 12705
rect 20705 12696 20717 12699
rect 20484 12668 20717 12696
rect 20484 12656 20490 12668
rect 20705 12665 20717 12668
rect 20751 12665 20763 12699
rect 20705 12659 20763 12665
rect 10858 12588 10864 12640
rect 10916 12628 10922 12640
rect 10953 12631 11011 12637
rect 10953 12628 10965 12631
rect 10916 12600 10965 12628
rect 10916 12588 10922 12600
rect 10953 12597 10965 12600
rect 10999 12597 11011 12631
rect 10953 12591 11011 12597
rect 11318 12588 11324 12640
rect 11376 12628 11382 12640
rect 11597 12631 11655 12637
rect 11597 12628 11609 12631
rect 11376 12600 11609 12628
rect 11376 12588 11382 12600
rect 11597 12597 11609 12600
rect 11643 12628 11655 12631
rect 11689 12631 11747 12637
rect 11689 12628 11701 12631
rect 11643 12600 11701 12628
rect 11643 12597 11655 12600
rect 11597 12591 11655 12597
rect 11689 12597 11701 12600
rect 11735 12597 11747 12631
rect 12238 12628 12244 12640
rect 12199 12600 12244 12628
rect 11689 12591 11747 12597
rect 12238 12588 12244 12600
rect 12296 12588 12302 12640
rect 13066 12628 13072 12640
rect 13027 12600 13072 12628
rect 13066 12588 13072 12600
rect 13124 12588 13130 12640
rect 16654 12628 16660 12640
rect 16615 12600 16660 12628
rect 16654 12588 16660 12600
rect 16712 12628 16718 12640
rect 17574 12628 17580 12640
rect 16712 12600 17580 12628
rect 16712 12588 16718 12600
rect 17574 12588 17580 12600
rect 17632 12588 17638 12640
rect 20720 12628 20748 12659
rect 22910 12656 22916 12708
rect 22968 12696 22974 12708
rect 23278 12696 23284 12708
rect 22968 12668 23048 12696
rect 23239 12668 23284 12696
rect 22968 12656 22974 12668
rect 23020 12637 23048 12668
rect 23278 12656 23284 12668
rect 23336 12656 23342 12708
rect 23373 12699 23431 12705
rect 23373 12665 23385 12699
rect 23419 12696 23431 12699
rect 23646 12696 23652 12708
rect 23419 12668 23652 12696
rect 23419 12665 23431 12668
rect 23373 12659 23431 12665
rect 21717 12631 21775 12637
rect 21717 12628 21729 12631
rect 20720 12600 21729 12628
rect 21717 12597 21729 12600
rect 21763 12597 21775 12631
rect 21717 12591 21775 12597
rect 23005 12631 23063 12637
rect 23005 12597 23017 12631
rect 23051 12628 23063 12631
rect 23388 12628 23416 12659
rect 23646 12656 23652 12668
rect 23704 12656 23710 12708
rect 23051 12600 23416 12628
rect 23051 12597 23063 12600
rect 23005 12591 23063 12597
rect 24290 12588 24296 12640
rect 24348 12628 24354 12640
rect 24937 12631 24995 12637
rect 24937 12628 24949 12631
rect 24348 12600 24949 12628
rect 24348 12588 24354 12600
rect 24937 12597 24949 12600
rect 24983 12597 24995 12631
rect 24937 12591 24995 12597
rect 632 12538 26392 12560
rect 632 12486 9843 12538
rect 9895 12486 9907 12538
rect 9959 12486 9971 12538
rect 10023 12486 10035 12538
rect 10087 12486 19176 12538
rect 19228 12486 19240 12538
rect 19292 12486 19304 12538
rect 19356 12486 19368 12538
rect 19420 12486 26392 12538
rect 632 12464 26392 12486
rect 10582 12424 10588 12436
rect 10495 12396 10588 12424
rect 10582 12384 10588 12396
rect 10640 12424 10646 12436
rect 12238 12424 12244 12436
rect 10640 12396 12244 12424
rect 10640 12384 10646 12396
rect 12238 12384 12244 12396
rect 12296 12384 12302 12436
rect 13069 12427 13127 12433
rect 13069 12393 13081 12427
rect 13115 12424 13127 12427
rect 13342 12424 13348 12436
rect 13115 12396 13348 12424
rect 13115 12393 13127 12396
rect 13069 12387 13127 12393
rect 13342 12384 13348 12396
rect 13400 12384 13406 12436
rect 13802 12424 13808 12436
rect 13763 12396 13808 12424
rect 13802 12384 13808 12396
rect 13860 12384 13866 12436
rect 13986 12384 13992 12436
rect 14044 12424 14050 12436
rect 14173 12427 14231 12433
rect 14173 12424 14185 12427
rect 14044 12396 14185 12424
rect 14044 12384 14050 12396
rect 14173 12393 14185 12396
rect 14219 12393 14231 12427
rect 16102 12424 16108 12436
rect 16063 12396 16108 12424
rect 14173 12387 14231 12393
rect 16102 12384 16108 12396
rect 16160 12384 16166 12436
rect 16654 12384 16660 12436
rect 16712 12424 16718 12436
rect 17301 12427 17359 12433
rect 17301 12424 17313 12427
rect 16712 12396 17313 12424
rect 16712 12384 16718 12396
rect 17301 12393 17313 12396
rect 17347 12393 17359 12427
rect 17301 12387 17359 12393
rect 19506 12384 19512 12436
rect 19564 12424 19570 12436
rect 19693 12427 19751 12433
rect 19693 12424 19705 12427
rect 19564 12396 19705 12424
rect 19564 12384 19570 12396
rect 19693 12393 19705 12396
rect 19739 12393 19751 12427
rect 19693 12387 19751 12393
rect 19782 12384 19788 12436
rect 19840 12424 19846 12436
rect 20886 12424 20892 12436
rect 19840 12396 20892 12424
rect 19840 12384 19846 12396
rect 20886 12384 20892 12396
rect 20944 12424 20950 12436
rect 21073 12427 21131 12433
rect 21073 12424 21085 12427
rect 20944 12396 21085 12424
rect 20944 12384 20950 12396
rect 21073 12393 21085 12396
rect 21119 12393 21131 12427
rect 21073 12387 21131 12393
rect 22269 12427 22327 12433
rect 22269 12393 22281 12427
rect 22315 12424 22327 12427
rect 22910 12424 22916 12436
rect 22315 12396 22916 12424
rect 22315 12393 22327 12396
rect 22269 12387 22327 12393
rect 22910 12384 22916 12396
rect 22968 12384 22974 12436
rect 25026 12433 25032 12436
rect 24983 12427 25032 12433
rect 24983 12393 24995 12427
rect 25029 12393 25032 12427
rect 24983 12387 25032 12393
rect 25026 12384 25032 12387
rect 25084 12384 25090 12436
rect 12514 12356 12520 12368
rect 12475 12328 12520 12356
rect 12514 12316 12520 12328
rect 12572 12316 12578 12368
rect 16473 12359 16531 12365
rect 16473 12325 16485 12359
rect 16519 12356 16531 12359
rect 16746 12356 16752 12368
rect 16519 12328 16752 12356
rect 16519 12325 16531 12328
rect 16473 12319 16531 12325
rect 16746 12316 16752 12328
rect 16804 12316 16810 12368
rect 17022 12356 17028 12368
rect 16983 12328 17028 12356
rect 17022 12316 17028 12328
rect 17080 12316 17086 12368
rect 18954 12316 18960 12368
rect 19012 12356 19018 12368
rect 19417 12359 19475 12365
rect 19417 12356 19429 12359
rect 19012 12328 19429 12356
rect 19012 12316 19018 12328
rect 19417 12325 19429 12328
rect 19463 12356 19475 12359
rect 19598 12356 19604 12368
rect 19463 12328 19604 12356
rect 19463 12325 19475 12328
rect 19417 12319 19475 12325
rect 19598 12316 19604 12328
rect 19656 12316 19662 12368
rect 20610 12316 20616 12368
rect 20668 12356 20674 12368
rect 21670 12359 21728 12365
rect 21670 12356 21682 12359
rect 20668 12328 21682 12356
rect 20668 12316 20674 12328
rect 21670 12325 21682 12328
rect 21716 12325 21728 12359
rect 21670 12319 21728 12325
rect 23002 12316 23008 12368
rect 23060 12356 23066 12368
rect 23465 12359 23523 12365
rect 23465 12356 23477 12359
rect 23060 12328 23477 12356
rect 23060 12316 23066 12328
rect 23465 12325 23477 12328
rect 23511 12356 23523 12359
rect 23830 12356 23836 12368
rect 23511 12328 23836 12356
rect 23511 12325 23523 12328
rect 23465 12319 23523 12325
rect 23830 12316 23836 12328
rect 23888 12316 23894 12368
rect 24290 12316 24296 12368
rect 24348 12316 24354 12368
rect 8101 12291 8159 12297
rect 8101 12257 8113 12291
rect 8147 12288 8159 12291
rect 8650 12288 8656 12300
rect 8147 12260 8656 12288
rect 8147 12257 8159 12260
rect 8101 12251 8159 12257
rect 8650 12248 8656 12260
rect 8708 12248 8714 12300
rect 10033 12291 10091 12297
rect 10033 12257 10045 12291
rect 10079 12288 10091 12291
rect 10214 12288 10220 12300
rect 10079 12260 10220 12288
rect 10079 12257 10091 12260
rect 10033 12251 10091 12257
rect 10214 12248 10220 12260
rect 10272 12248 10278 12300
rect 10490 12248 10496 12300
rect 10548 12288 10554 12300
rect 11042 12288 11048 12300
rect 10548 12260 11048 12288
rect 10548 12248 10554 12260
rect 11042 12248 11048 12260
rect 11100 12288 11106 12300
rect 13161 12291 13219 12297
rect 13161 12288 13173 12291
rect 11100 12260 13173 12288
rect 11100 12248 11106 12260
rect 13161 12257 13173 12260
rect 13207 12257 13219 12291
rect 13161 12251 13219 12257
rect 10953 12223 11011 12229
rect 10953 12189 10965 12223
rect 10999 12220 11011 12223
rect 11410 12220 11416 12232
rect 10999 12192 11416 12220
rect 10999 12189 11011 12192
rect 10953 12183 11011 12189
rect 11410 12180 11416 12192
rect 11468 12180 11474 12232
rect 13176 12220 13204 12251
rect 18126 12248 18132 12300
rect 18184 12288 18190 12300
rect 18310 12288 18316 12300
rect 18184 12260 18316 12288
rect 18184 12248 18190 12260
rect 18310 12248 18316 12260
rect 18368 12248 18374 12300
rect 19049 12291 19107 12297
rect 19049 12257 19061 12291
rect 19095 12288 19107 12291
rect 19690 12288 19696 12300
rect 19095 12260 19696 12288
rect 19095 12257 19107 12260
rect 19049 12251 19107 12257
rect 19690 12248 19696 12260
rect 19748 12248 19754 12300
rect 21349 12291 21407 12297
rect 21349 12257 21361 12291
rect 21395 12288 21407 12291
rect 21898 12288 21904 12300
rect 21395 12260 21904 12288
rect 21395 12257 21407 12260
rect 21349 12251 21407 12257
rect 21898 12248 21904 12260
rect 21956 12288 21962 12300
rect 23186 12288 23192 12300
rect 21956 12260 23192 12288
rect 21956 12248 21962 12260
rect 23186 12248 23192 12260
rect 23244 12248 23250 12300
rect 13434 12220 13440 12232
rect 13176 12192 13440 12220
rect 13434 12180 13440 12192
rect 13492 12180 13498 12232
rect 13529 12223 13587 12229
rect 13529 12189 13541 12223
rect 13575 12220 13587 12223
rect 13618 12220 13624 12232
rect 13575 12192 13624 12220
rect 13575 12189 13587 12192
rect 13529 12183 13587 12189
rect 13618 12180 13624 12192
rect 13676 12180 13682 12232
rect 15277 12223 15335 12229
rect 15277 12189 15289 12223
rect 15323 12220 15335 12223
rect 15734 12220 15740 12232
rect 15323 12192 15740 12220
rect 15323 12189 15335 12192
rect 15277 12183 15335 12189
rect 15734 12180 15740 12192
rect 15792 12180 15798 12232
rect 16381 12223 16439 12229
rect 16381 12189 16393 12223
rect 16427 12220 16439 12223
rect 16654 12220 16660 12232
rect 16427 12192 16660 12220
rect 16427 12189 16439 12192
rect 16381 12183 16439 12189
rect 16654 12180 16660 12192
rect 16712 12180 16718 12232
rect 18681 12223 18739 12229
rect 18681 12220 18693 12223
rect 17776 12192 18693 12220
rect 14538 12152 14544 12164
rect 14499 12124 14544 12152
rect 14538 12112 14544 12124
rect 14596 12112 14602 12164
rect 8282 12084 8288 12096
rect 8243 12056 8288 12084
rect 8282 12044 8288 12056
rect 8340 12044 8346 12096
rect 9938 12084 9944 12096
rect 9899 12056 9944 12084
rect 9938 12044 9944 12056
rect 9996 12044 10002 12096
rect 11226 12093 11232 12096
rect 10217 12087 10275 12093
rect 10217 12053 10229 12087
rect 10263 12084 10275 12087
rect 11210 12087 11232 12093
rect 11210 12084 11222 12087
rect 10263 12056 11222 12084
rect 10263 12053 10275 12056
rect 10217 12047 10275 12053
rect 11210 12053 11222 12056
rect 11210 12047 11232 12053
rect 11226 12044 11232 12047
rect 11284 12044 11290 12096
rect 11318 12044 11324 12096
rect 11376 12084 11382 12096
rect 11502 12084 11508 12096
rect 11376 12056 11421 12084
rect 11463 12056 11508 12084
rect 11376 12044 11382 12056
rect 11502 12044 11508 12056
rect 11560 12044 11566 12096
rect 11962 12044 11968 12096
rect 12020 12084 12026 12096
rect 12149 12087 12207 12093
rect 12149 12084 12161 12087
rect 12020 12056 12161 12084
rect 12020 12044 12026 12056
rect 12149 12053 12161 12056
rect 12195 12084 12207 12087
rect 12330 12084 12336 12096
rect 12195 12056 12336 12084
rect 12195 12053 12207 12056
rect 12149 12047 12207 12053
rect 12330 12044 12336 12056
rect 12388 12044 12394 12096
rect 13342 12093 13348 12096
rect 13326 12087 13348 12093
rect 13326 12053 13338 12087
rect 13326 12047 13348 12053
rect 13342 12044 13348 12047
rect 13400 12044 13406 12096
rect 13437 12087 13495 12093
rect 13437 12053 13449 12087
rect 13483 12084 13495 12087
rect 14078 12084 14084 12096
rect 13483 12056 14084 12084
rect 13483 12053 13495 12056
rect 13437 12047 13495 12053
rect 14078 12044 14084 12056
rect 14136 12044 14142 12096
rect 15826 12084 15832 12096
rect 15787 12056 15832 12084
rect 15826 12044 15832 12056
rect 15884 12044 15890 12096
rect 17298 12044 17304 12096
rect 17356 12084 17362 12096
rect 17776 12093 17804 12192
rect 18681 12189 18693 12192
rect 18727 12220 18739 12223
rect 18862 12220 18868 12232
rect 18727 12192 18868 12220
rect 18727 12189 18739 12192
rect 18681 12183 18739 12189
rect 18862 12180 18868 12192
rect 18920 12220 18926 12232
rect 20242 12220 20248 12232
rect 18920 12192 20248 12220
rect 18920 12180 18926 12192
rect 20242 12180 20248 12192
rect 20300 12180 20306 12232
rect 23373 12223 23431 12229
rect 23373 12189 23385 12223
rect 23419 12220 23431 12223
rect 23462 12220 23468 12232
rect 23419 12192 23468 12220
rect 23419 12189 23431 12192
rect 23373 12183 23431 12189
rect 23462 12180 23468 12192
rect 23520 12180 23526 12232
rect 23646 12220 23652 12232
rect 23607 12192 23652 12220
rect 23646 12180 23652 12192
rect 23704 12180 23710 12232
rect 18034 12112 18040 12164
rect 18092 12152 18098 12164
rect 18451 12155 18509 12161
rect 18451 12152 18463 12155
rect 18092 12124 18463 12152
rect 18092 12112 18098 12124
rect 18451 12121 18463 12124
rect 18497 12152 18509 12155
rect 18770 12152 18776 12164
rect 18497 12124 18776 12152
rect 18497 12121 18509 12124
rect 18451 12115 18509 12121
rect 18770 12112 18776 12124
rect 18828 12112 18834 12164
rect 19598 12112 19604 12164
rect 19656 12152 19662 12164
rect 20702 12152 20708 12164
rect 19656 12124 20708 12152
rect 19656 12112 19662 12124
rect 20702 12112 20708 12124
rect 20760 12112 20766 12164
rect 23554 12112 23560 12164
rect 23612 12152 23618 12164
rect 24106 12152 24112 12164
rect 23612 12124 24112 12152
rect 23612 12112 23618 12124
rect 24106 12112 24112 12124
rect 24164 12112 24170 12164
rect 24308 12096 24336 12316
rect 24842 12248 24848 12300
rect 24900 12297 24906 12300
rect 24900 12291 24938 12297
rect 24926 12257 24938 12291
rect 24900 12251 24938 12257
rect 24900 12248 24906 12251
rect 17761 12087 17819 12093
rect 17761 12084 17773 12087
rect 17356 12056 17773 12084
rect 17356 12044 17362 12056
rect 17761 12053 17773 12056
rect 17807 12053 17819 12087
rect 18218 12084 18224 12096
rect 18179 12056 18224 12084
rect 17761 12047 17819 12053
rect 18218 12044 18224 12056
rect 18276 12044 18282 12096
rect 18586 12044 18592 12096
rect 18644 12084 18650 12096
rect 20245 12087 20303 12093
rect 18644 12056 18689 12084
rect 18644 12044 18650 12056
rect 20245 12053 20257 12087
rect 20291 12084 20303 12087
rect 20334 12084 20340 12096
rect 20291 12056 20340 12084
rect 20291 12053 20303 12056
rect 20245 12047 20303 12053
rect 20334 12044 20340 12056
rect 20392 12044 20398 12096
rect 22542 12084 22548 12096
rect 22503 12056 22548 12084
rect 22542 12044 22548 12056
rect 22600 12044 22606 12096
rect 24290 12044 24296 12096
rect 24348 12044 24354 12096
rect 632 11994 26392 12016
rect 632 11942 5176 11994
rect 5228 11942 5240 11994
rect 5292 11942 5304 11994
rect 5356 11942 5368 11994
rect 5420 11942 14510 11994
rect 14562 11942 14574 11994
rect 14626 11942 14638 11994
rect 14690 11942 14702 11994
rect 14754 11942 23843 11994
rect 23895 11942 23907 11994
rect 23959 11942 23971 11994
rect 24023 11942 24035 11994
rect 24087 11942 26392 11994
rect 632 11920 26392 11942
rect 7730 11880 7736 11892
rect 7691 11852 7736 11880
rect 7730 11840 7736 11852
rect 7788 11840 7794 11892
rect 8650 11880 8656 11892
rect 8611 11852 8656 11880
rect 8650 11840 8656 11852
rect 8708 11840 8714 11892
rect 9386 11880 9392 11892
rect 9347 11852 9392 11880
rect 9386 11840 9392 11852
rect 9444 11840 9450 11892
rect 10125 11883 10183 11889
rect 10125 11849 10137 11883
rect 10171 11880 10183 11883
rect 10214 11880 10220 11892
rect 10171 11852 10220 11880
rect 10171 11849 10183 11852
rect 10125 11843 10183 11849
rect 10214 11840 10220 11852
rect 10272 11840 10278 11892
rect 11134 11840 11140 11892
rect 11192 11880 11198 11892
rect 11229 11883 11287 11889
rect 11229 11880 11241 11883
rect 11192 11852 11241 11880
rect 11192 11840 11198 11852
rect 11229 11849 11241 11852
rect 11275 11880 11287 11883
rect 11318 11880 11324 11892
rect 11275 11852 11324 11880
rect 11275 11849 11287 11852
rect 11229 11843 11287 11849
rect 11318 11840 11324 11852
rect 11376 11840 11382 11892
rect 13253 11883 13311 11889
rect 13253 11849 13265 11883
rect 13299 11880 13311 11883
rect 13618 11880 13624 11892
rect 13299 11852 13624 11880
rect 13299 11849 13311 11852
rect 13253 11843 13311 11849
rect 13618 11840 13624 11852
rect 13676 11840 13682 11892
rect 14170 11840 14176 11892
rect 14228 11880 14234 11892
rect 14265 11883 14323 11889
rect 14265 11880 14277 11883
rect 14228 11852 14277 11880
rect 14228 11840 14234 11852
rect 14265 11849 14277 11852
rect 14311 11849 14323 11883
rect 15182 11880 15188 11892
rect 15143 11852 15188 11880
rect 14265 11843 14323 11849
rect 15182 11840 15188 11852
rect 15240 11840 15246 11892
rect 16473 11883 16531 11889
rect 16473 11849 16485 11883
rect 16519 11880 16531 11883
rect 16746 11880 16752 11892
rect 16519 11852 16752 11880
rect 16519 11849 16531 11852
rect 16473 11843 16531 11849
rect 16746 11840 16752 11852
rect 16804 11840 16810 11892
rect 17298 11880 17304 11892
rect 17259 11852 17304 11880
rect 17298 11840 17304 11852
rect 17356 11840 17362 11892
rect 18678 11840 18684 11892
rect 18736 11880 18742 11892
rect 18846 11883 18904 11889
rect 18846 11880 18858 11883
rect 18736 11852 18858 11880
rect 18736 11840 18742 11852
rect 18846 11849 18858 11852
rect 18892 11880 18904 11883
rect 19782 11880 19788 11892
rect 18892 11852 19788 11880
rect 18892 11849 18904 11852
rect 18846 11843 18904 11849
rect 19782 11840 19788 11852
rect 19840 11840 19846 11892
rect 20245 11883 20303 11889
rect 20245 11849 20257 11883
rect 20291 11880 20303 11883
rect 20794 11880 20800 11892
rect 20291 11852 20800 11880
rect 20291 11849 20303 11852
rect 20245 11843 20303 11849
rect 9110 11812 9116 11824
rect 9071 11784 9116 11812
rect 9110 11772 9116 11784
rect 9168 11772 9174 11824
rect 12238 11812 12244 11824
rect 12199 11784 12244 11812
rect 12238 11772 12244 11784
rect 12296 11772 12302 11824
rect 13713 11815 13771 11821
rect 13713 11781 13725 11815
rect 13759 11812 13771 11815
rect 13943 11815 14001 11821
rect 13943 11812 13955 11815
rect 13759 11784 13955 11812
rect 13759 11781 13771 11784
rect 13713 11775 13771 11781
rect 13943 11781 13955 11784
rect 13989 11781 14001 11815
rect 13943 11775 14001 11781
rect 7181 11679 7239 11685
rect 7181 11645 7193 11679
rect 7227 11676 7239 11679
rect 7730 11676 7736 11688
rect 7227 11648 7736 11676
rect 7227 11645 7239 11648
rect 7181 11639 7239 11645
rect 7730 11636 7736 11648
rect 7788 11636 7794 11688
rect 8193 11679 8251 11685
rect 8193 11645 8205 11679
rect 8239 11676 8251 11679
rect 9128 11676 9156 11772
rect 12330 11744 12336 11756
rect 12291 11716 12336 11744
rect 12330 11704 12336 11716
rect 12388 11704 12394 11756
rect 8239 11648 9156 11676
rect 9205 11679 9263 11685
rect 8239 11645 8251 11648
rect 8193 11639 8251 11645
rect 9205 11645 9217 11679
rect 9251 11645 9263 11679
rect 9205 11639 9263 11645
rect 8098 11568 8104 11620
rect 8156 11608 8162 11620
rect 9220 11608 9248 11639
rect 9938 11636 9944 11688
rect 9996 11676 10002 11688
rect 10214 11676 10220 11688
rect 9996 11648 10220 11676
rect 9996 11636 10002 11648
rect 10214 11636 10220 11648
rect 10272 11636 10278 11688
rect 10766 11676 10772 11688
rect 10679 11648 10772 11676
rect 10766 11636 10772 11648
rect 10824 11676 10830 11688
rect 11502 11676 11508 11688
rect 10824 11648 11508 11676
rect 10824 11636 10830 11648
rect 11502 11636 11508 11648
rect 11560 11636 11566 11688
rect 12054 11676 12060 11688
rect 12022 11648 12060 11676
rect 12054 11636 12060 11648
rect 12112 11685 12118 11688
rect 12112 11679 12170 11685
rect 12112 11645 12124 11679
rect 12158 11676 12170 11679
rect 12422 11676 12428 11688
rect 12158 11648 12428 11676
rect 12158 11645 12170 11648
rect 12112 11639 12170 11645
rect 12112 11636 12118 11639
rect 12422 11636 12428 11648
rect 12480 11636 12486 11688
rect 13958 11676 13986 11775
rect 14078 11772 14084 11824
rect 14136 11812 14142 11824
rect 14998 11812 15004 11824
rect 14136 11784 15004 11812
rect 14136 11772 14142 11784
rect 14998 11772 15004 11784
rect 15056 11772 15062 11824
rect 18494 11772 18500 11824
rect 18552 11812 18558 11824
rect 18957 11815 19015 11821
rect 18957 11812 18969 11815
rect 18552 11784 18969 11812
rect 18552 11772 18558 11784
rect 18957 11781 18969 11784
rect 19003 11812 19015 11815
rect 19598 11812 19604 11824
rect 19003 11784 19604 11812
rect 19003 11781 19015 11784
rect 18957 11775 19015 11781
rect 19598 11772 19604 11784
rect 19656 11772 19662 11824
rect 14173 11747 14231 11753
rect 14173 11713 14185 11747
rect 14219 11744 14231 11747
rect 14262 11744 14268 11756
rect 14219 11716 14268 11744
rect 14219 11713 14231 11716
rect 14173 11707 14231 11713
rect 14262 11704 14268 11716
rect 14320 11704 14326 11756
rect 18034 11744 18040 11756
rect 15108 11716 18040 11744
rect 15108 11676 15136 11716
rect 18034 11704 18040 11716
rect 18092 11744 18098 11756
rect 18129 11747 18187 11753
rect 18129 11744 18141 11747
rect 18092 11716 18141 11744
rect 18092 11704 18098 11716
rect 18129 11713 18141 11716
rect 18175 11713 18187 11747
rect 18129 11707 18187 11713
rect 18862 11704 18868 11756
rect 18920 11744 18926 11756
rect 19049 11747 19107 11753
rect 19049 11744 19061 11747
rect 18920 11716 19061 11744
rect 18920 11704 18926 11716
rect 19049 11713 19061 11716
rect 19095 11713 19107 11747
rect 19049 11707 19107 11713
rect 13958 11648 15136 11676
rect 15182 11636 15188 11688
rect 15240 11676 15246 11688
rect 15369 11679 15427 11685
rect 15369 11676 15381 11679
rect 15240 11648 15381 11676
rect 15240 11636 15246 11648
rect 15369 11645 15381 11648
rect 15415 11645 15427 11679
rect 15826 11676 15832 11688
rect 15739 11648 15832 11676
rect 15369 11639 15427 11645
rect 15826 11636 15832 11648
rect 15884 11636 15890 11688
rect 17666 11636 17672 11688
rect 17724 11685 17730 11688
rect 17724 11679 17762 11685
rect 17750 11645 17762 11679
rect 17724 11639 17762 11645
rect 17807 11679 17865 11685
rect 17807 11645 17819 11679
rect 17853 11676 17865 11679
rect 18770 11676 18776 11688
rect 17853 11648 18776 11676
rect 17853 11645 17865 11648
rect 17807 11639 17865 11645
rect 17724 11636 17730 11639
rect 18770 11636 18776 11648
rect 18828 11636 18834 11688
rect 20444 11685 20472 11852
rect 20794 11840 20800 11852
rect 20852 11840 20858 11892
rect 23002 11880 23008 11892
rect 22963 11852 23008 11880
rect 23002 11840 23008 11852
rect 23060 11840 23066 11892
rect 24753 11883 24811 11889
rect 24753 11849 24765 11883
rect 24799 11880 24811 11883
rect 24842 11880 24848 11892
rect 24799 11852 24848 11880
rect 24799 11849 24811 11852
rect 24753 11843 24811 11849
rect 24842 11840 24848 11852
rect 24900 11840 24906 11892
rect 24293 11815 24351 11821
rect 24293 11812 24305 11815
rect 23388 11784 24305 11812
rect 20610 11704 20616 11756
rect 20668 11744 20674 11756
rect 20797 11747 20855 11753
rect 20797 11744 20809 11747
rect 20668 11716 20809 11744
rect 20668 11704 20674 11716
rect 20797 11713 20809 11716
rect 20843 11744 20855 11747
rect 21165 11747 21223 11753
rect 21165 11744 21177 11747
rect 20843 11716 21177 11744
rect 20843 11713 20855 11716
rect 20797 11707 20855 11713
rect 21165 11713 21177 11716
rect 21211 11744 21223 11747
rect 21530 11744 21536 11756
rect 21211 11716 21536 11744
rect 21211 11713 21223 11716
rect 21165 11707 21223 11713
rect 21530 11704 21536 11716
rect 21588 11744 21594 11756
rect 21588 11716 21713 11744
rect 21588 11704 21594 11716
rect 20404 11679 20472 11685
rect 20404 11645 20416 11679
rect 20450 11648 20472 11679
rect 21346 11676 21352 11688
rect 21307 11648 21352 11676
rect 20450 11645 20462 11648
rect 20404 11639 20462 11645
rect 21346 11636 21352 11648
rect 21404 11636 21410 11688
rect 9662 11608 9668 11620
rect 8156 11580 9668 11608
rect 8156 11568 8162 11580
rect 9662 11568 9668 11580
rect 9720 11568 9726 11620
rect 11962 11568 11968 11620
rect 12020 11608 12026 11620
rect 12020 11580 12065 11608
rect 12020 11568 12026 11580
rect 13710 11568 13716 11620
rect 13768 11608 13774 11620
rect 13805 11611 13863 11617
rect 13805 11608 13817 11611
rect 13768 11580 13817 11608
rect 13768 11568 13774 11580
rect 13805 11577 13817 11580
rect 13851 11608 13863 11611
rect 13986 11608 13992 11620
rect 13851 11580 13992 11608
rect 13851 11577 13863 11580
rect 13805 11571 13863 11577
rect 13986 11568 13992 11580
rect 14044 11568 14050 11620
rect 14909 11611 14967 11617
rect 14909 11577 14921 11611
rect 14955 11608 14967 11611
rect 14998 11608 15004 11620
rect 14955 11580 15004 11608
rect 14955 11577 14967 11580
rect 14909 11571 14967 11577
rect 14998 11568 15004 11580
rect 15056 11568 15062 11620
rect 15274 11568 15280 11620
rect 15332 11608 15338 11620
rect 15844 11608 15872 11636
rect 15332 11580 15872 11608
rect 15332 11568 15338 11580
rect 18586 11568 18592 11620
rect 18644 11608 18650 11620
rect 18681 11611 18739 11617
rect 18681 11608 18693 11611
rect 18644 11580 18693 11608
rect 18644 11568 18650 11580
rect 18681 11577 18693 11580
rect 18727 11577 18739 11611
rect 18681 11571 18739 11577
rect 19417 11611 19475 11617
rect 19417 11577 19429 11611
rect 19463 11608 19475 11611
rect 20886 11608 20892 11620
rect 19463 11580 20892 11608
rect 19463 11577 19475 11580
rect 19417 11571 19475 11577
rect 20886 11568 20892 11580
rect 20944 11568 20950 11620
rect 21685 11617 21713 11716
rect 23094 11704 23100 11756
rect 23152 11744 23158 11756
rect 23388 11753 23416 11784
rect 24293 11781 24305 11784
rect 24339 11781 24351 11815
rect 24293 11775 24351 11781
rect 23373 11747 23431 11753
rect 23373 11744 23385 11747
rect 23152 11716 23385 11744
rect 23152 11704 23158 11716
rect 23373 11713 23385 11716
rect 23419 11713 23431 11747
rect 23646 11744 23652 11756
rect 23607 11716 23652 11744
rect 23373 11707 23431 11713
rect 23646 11704 23652 11716
rect 23704 11704 23710 11756
rect 24842 11676 24848 11688
rect 24803 11648 24848 11676
rect 24842 11636 24848 11648
rect 24900 11676 24906 11688
rect 25397 11679 25455 11685
rect 25397 11676 25409 11679
rect 24900 11648 25409 11676
rect 24900 11636 24906 11648
rect 25397 11645 25409 11648
rect 25443 11645 25455 11679
rect 25397 11639 25455 11645
rect 21670 11611 21728 11617
rect 21670 11577 21682 11611
rect 21716 11577 21728 11611
rect 21670 11571 21728 11577
rect 23465 11611 23523 11617
rect 23465 11577 23477 11611
rect 23511 11608 23523 11611
rect 23554 11608 23560 11620
rect 23511 11580 23560 11608
rect 23511 11577 23523 11580
rect 23465 11571 23523 11577
rect 7362 11540 7368 11552
rect 7323 11512 7368 11540
rect 7362 11500 7368 11512
rect 7420 11500 7426 11552
rect 8374 11540 8380 11552
rect 8335 11512 8380 11540
rect 8374 11500 8380 11512
rect 8432 11500 8438 11552
rect 10493 11543 10551 11549
rect 10493 11509 10505 11543
rect 10539 11540 10551 11543
rect 10582 11540 10588 11552
rect 10539 11512 10588 11540
rect 10539 11509 10551 11512
rect 10493 11503 10551 11509
rect 10582 11500 10588 11512
rect 10640 11500 10646 11552
rect 11686 11540 11692 11552
rect 11647 11512 11692 11540
rect 11686 11500 11692 11512
rect 11744 11500 11750 11552
rect 12606 11540 12612 11552
rect 12567 11512 12612 11540
rect 12606 11500 12612 11512
rect 12664 11500 12670 11552
rect 15458 11540 15464 11552
rect 15419 11512 15464 11540
rect 15458 11500 15464 11512
rect 15516 11500 15522 11552
rect 16746 11540 16752 11552
rect 16707 11512 16752 11540
rect 16746 11500 16752 11512
rect 16804 11500 16810 11552
rect 18402 11500 18408 11552
rect 18460 11540 18466 11552
rect 18497 11543 18555 11549
rect 18497 11540 18509 11543
rect 18460 11512 18509 11540
rect 18460 11500 18466 11512
rect 18497 11509 18509 11512
rect 18543 11509 18555 11543
rect 18497 11503 18555 11509
rect 20475 11543 20533 11549
rect 20475 11509 20487 11543
rect 20521 11540 20533 11543
rect 20702 11540 20708 11552
rect 20521 11512 20708 11540
rect 20521 11509 20533 11512
rect 20475 11503 20533 11509
rect 20702 11500 20708 11512
rect 20760 11500 20766 11552
rect 22269 11543 22327 11549
rect 22269 11509 22281 11543
rect 22315 11540 22327 11543
rect 22637 11543 22695 11549
rect 22637 11540 22649 11543
rect 22315 11512 22649 11540
rect 22315 11509 22327 11512
rect 22269 11503 22327 11509
rect 22637 11509 22649 11512
rect 22683 11540 22695 11543
rect 23480 11540 23508 11571
rect 23554 11568 23560 11580
rect 23612 11568 23618 11620
rect 23646 11568 23652 11620
rect 23704 11608 23710 11620
rect 24934 11608 24940 11620
rect 23704 11580 24940 11608
rect 23704 11568 23710 11580
rect 24934 11568 24940 11580
rect 24992 11568 24998 11620
rect 22683 11512 23508 11540
rect 22683 11509 22695 11512
rect 22637 11503 22695 11509
rect 23738 11500 23744 11552
rect 23796 11540 23802 11552
rect 24290 11540 24296 11552
rect 23796 11512 24296 11540
rect 23796 11500 23802 11512
rect 24290 11500 24296 11512
rect 24348 11500 24354 11552
rect 24382 11500 24388 11552
rect 24440 11540 24446 11552
rect 25029 11543 25087 11549
rect 25029 11540 25041 11543
rect 24440 11512 25041 11540
rect 24440 11500 24446 11512
rect 25029 11509 25041 11512
rect 25075 11509 25087 11543
rect 25029 11503 25087 11509
rect 632 11450 26392 11472
rect 632 11398 9843 11450
rect 9895 11398 9907 11450
rect 9959 11398 9971 11450
rect 10023 11398 10035 11450
rect 10087 11398 19176 11450
rect 19228 11398 19240 11450
rect 19292 11398 19304 11450
rect 19356 11398 19368 11450
rect 19420 11398 26392 11450
rect 632 11376 26392 11398
rect 9386 11296 9392 11348
rect 9444 11336 9450 11348
rect 10033 11339 10091 11345
rect 10033 11336 10045 11339
rect 9444 11308 10045 11336
rect 9444 11296 9450 11308
rect 10033 11305 10045 11308
rect 10079 11336 10091 11339
rect 10214 11336 10220 11348
rect 10079 11308 10220 11336
rect 10079 11305 10091 11308
rect 10033 11299 10091 11305
rect 10214 11296 10220 11308
rect 10272 11296 10278 11348
rect 10953 11339 11011 11345
rect 10953 11305 10965 11339
rect 10999 11336 11011 11339
rect 11042 11336 11048 11348
rect 10999 11308 11048 11336
rect 10999 11305 11011 11308
rect 10953 11299 11011 11305
rect 11042 11296 11048 11308
rect 11100 11296 11106 11348
rect 12149 11339 12207 11345
rect 12149 11305 12161 11339
rect 12195 11336 12207 11339
rect 12238 11336 12244 11348
rect 12195 11308 12244 11336
rect 12195 11305 12207 11308
rect 12149 11299 12207 11305
rect 12238 11296 12244 11308
rect 12296 11296 12302 11348
rect 12422 11336 12428 11348
rect 12383 11308 12428 11336
rect 12422 11296 12428 11308
rect 12480 11296 12486 11348
rect 13434 11296 13440 11348
rect 13492 11336 13498 11348
rect 13621 11339 13679 11345
rect 13621 11336 13633 11339
rect 13492 11308 13633 11336
rect 13492 11296 13498 11308
rect 13621 11305 13633 11308
rect 13667 11305 13679 11339
rect 13621 11299 13679 11305
rect 13894 11296 13900 11348
rect 13952 11336 13958 11348
rect 13989 11339 14047 11345
rect 13989 11336 14001 11339
rect 13952 11308 14001 11336
rect 13952 11296 13958 11308
rect 13989 11305 14001 11308
rect 14035 11305 14047 11339
rect 13989 11299 14047 11305
rect 14449 11339 14507 11345
rect 14449 11305 14461 11339
rect 14495 11336 14507 11339
rect 14998 11336 15004 11348
rect 14495 11308 15004 11336
rect 14495 11305 14507 11308
rect 14449 11299 14507 11305
rect 14998 11296 15004 11308
rect 15056 11296 15062 11348
rect 16470 11336 16476 11348
rect 16431 11308 16476 11336
rect 16470 11296 16476 11308
rect 16528 11296 16534 11348
rect 21346 11296 21352 11348
rect 21404 11336 21410 11348
rect 22269 11339 22327 11345
rect 22269 11336 22281 11339
rect 21404 11308 22281 11336
rect 21404 11296 21410 11308
rect 22269 11305 22281 11308
rect 22315 11336 22327 11339
rect 23462 11336 23468 11348
rect 22315 11308 22864 11336
rect 23423 11308 23468 11336
rect 22315 11305 22327 11308
rect 22269 11299 22327 11305
rect 9294 11228 9300 11280
rect 9352 11268 9358 11280
rect 11686 11268 11692 11280
rect 9352 11240 11692 11268
rect 9352 11228 9358 11240
rect 8098 11200 8104 11212
rect 8059 11172 8104 11200
rect 8098 11160 8104 11172
rect 8156 11160 8162 11212
rect 9662 11160 9668 11212
rect 9720 11200 9726 11212
rect 11060 11209 11088 11240
rect 11686 11228 11692 11240
rect 11744 11228 11750 11280
rect 12330 11228 12336 11280
rect 12388 11268 12394 11280
rect 12609 11271 12667 11277
rect 12609 11268 12621 11271
rect 12388 11240 12621 11268
rect 12388 11228 12394 11240
rect 12609 11237 12621 11240
rect 12655 11237 12667 11271
rect 12609 11231 12667 11237
rect 14354 11228 14360 11280
rect 14412 11268 14418 11280
rect 14817 11271 14875 11277
rect 14817 11268 14829 11271
rect 14412 11240 14829 11268
rect 14412 11228 14418 11240
rect 14817 11237 14829 11240
rect 14863 11237 14875 11271
rect 14817 11231 14875 11237
rect 16289 11271 16347 11277
rect 16289 11237 16301 11271
rect 16335 11268 16347 11271
rect 17666 11268 17672 11280
rect 16335 11240 17672 11268
rect 16335 11237 16347 11240
rect 16289 11231 16347 11237
rect 17666 11228 17672 11240
rect 17724 11228 17730 11280
rect 18494 11228 18500 11280
rect 18552 11268 18558 11280
rect 19693 11271 19751 11277
rect 19693 11268 19705 11271
rect 18552 11240 19705 11268
rect 18552 11228 18558 11240
rect 19693 11237 19705 11240
rect 19739 11237 19751 11271
rect 19693 11231 19751 11237
rect 20702 11228 20708 11280
rect 20760 11268 20766 11280
rect 21898 11268 21904 11280
rect 20760 11240 21760 11268
rect 21859 11240 21904 11268
rect 20760 11228 20766 11240
rect 9849 11203 9907 11209
rect 9849 11200 9861 11203
rect 9720 11172 9861 11200
rect 9720 11160 9726 11172
rect 9849 11169 9861 11172
rect 9895 11169 9907 11203
rect 9849 11163 9907 11169
rect 11045 11203 11103 11209
rect 11045 11169 11057 11203
rect 11091 11169 11103 11203
rect 11045 11163 11103 11169
rect 13066 11160 13072 11212
rect 13124 11200 13130 11212
rect 13253 11203 13311 11209
rect 13253 11200 13265 11203
rect 13124 11172 13265 11200
rect 13124 11160 13130 11172
rect 13253 11169 13265 11172
rect 13299 11200 13311 11203
rect 13618 11200 13624 11212
rect 13299 11172 13624 11200
rect 13299 11169 13311 11172
rect 13253 11163 13311 11169
rect 13618 11160 13624 11172
rect 13676 11160 13682 11212
rect 16378 11160 16384 11212
rect 16436 11200 16442 11212
rect 16654 11200 16660 11212
rect 16436 11172 16660 11200
rect 16436 11160 16442 11172
rect 16654 11160 16660 11172
rect 16712 11160 16718 11212
rect 16841 11203 16899 11209
rect 16841 11169 16853 11203
rect 16887 11169 16899 11203
rect 16841 11163 16899 11169
rect 10585 11135 10643 11141
rect 10585 11101 10597 11135
rect 10631 11132 10643 11135
rect 11410 11132 11416 11144
rect 10631 11104 10996 11132
rect 11371 11104 11416 11132
rect 10631 11101 10643 11104
rect 10585 11095 10643 11101
rect 8282 11064 8288 11076
rect 8243 11036 8288 11064
rect 8282 11024 8288 11036
rect 8340 11024 8346 11076
rect 9757 11067 9815 11073
rect 9757 11033 9769 11067
rect 9803 11064 9815 11067
rect 10766 11064 10772 11076
rect 9803 11036 10772 11064
rect 9803 11033 9815 11036
rect 9757 11027 9815 11033
rect 10766 11024 10772 11036
rect 10824 11024 10830 11076
rect 10968 11064 10996 11104
rect 11410 11092 11416 11104
rect 11468 11092 11474 11144
rect 11502 11092 11508 11144
rect 11560 11132 11566 11144
rect 15182 11132 15188 11144
rect 11560 11104 11605 11132
rect 15143 11104 15188 11132
rect 11560 11092 11566 11104
rect 15182 11092 15188 11104
rect 15240 11092 15246 11144
rect 16194 11092 16200 11144
rect 16252 11132 16258 11144
rect 16856 11132 16884 11163
rect 17482 11160 17488 11212
rect 17540 11200 17546 11212
rect 18126 11200 18132 11212
rect 17540 11172 18132 11200
rect 17540 11160 17546 11172
rect 18126 11160 18132 11172
rect 18184 11200 18190 11212
rect 18681 11203 18739 11209
rect 18681 11200 18693 11203
rect 18184 11172 18693 11200
rect 18184 11160 18190 11172
rect 18681 11169 18693 11172
rect 18727 11200 18739 11203
rect 18770 11200 18776 11212
rect 18727 11172 18776 11200
rect 18727 11169 18739 11172
rect 18681 11163 18739 11169
rect 18770 11160 18776 11172
rect 18828 11160 18834 11212
rect 20426 11200 20432 11212
rect 20387 11172 20432 11200
rect 20426 11160 20432 11172
rect 20484 11160 20490 11212
rect 20886 11200 20892 11212
rect 20847 11172 20892 11200
rect 20886 11160 20892 11172
rect 20944 11200 20950 11212
rect 21441 11203 21499 11209
rect 21441 11200 21453 11203
rect 20944 11172 21453 11200
rect 20944 11160 20950 11172
rect 21441 11169 21453 11172
rect 21487 11169 21499 11203
rect 21441 11163 21499 11169
rect 17393 11135 17451 11141
rect 17393 11132 17405 11135
rect 16252 11104 17405 11132
rect 16252 11092 16258 11104
rect 17393 11101 17405 11104
rect 17439 11132 17451 11135
rect 18034 11132 18040 11144
rect 17439 11104 18040 11132
rect 17439 11101 17451 11104
rect 17393 11095 17451 11101
rect 18034 11092 18040 11104
rect 18092 11092 18098 11144
rect 18954 11092 18960 11144
rect 19012 11132 19018 11144
rect 19049 11135 19107 11141
rect 19049 11132 19061 11135
rect 19012 11104 19061 11132
rect 19012 11092 19018 11104
rect 19049 11101 19061 11104
rect 19095 11101 19107 11135
rect 20978 11132 20984 11144
rect 20939 11104 20984 11132
rect 19049 11095 19107 11101
rect 20978 11092 20984 11104
rect 21036 11092 21042 11144
rect 21732 11132 21760 11240
rect 21898 11228 21904 11240
rect 21956 11228 21962 11280
rect 22637 11271 22695 11277
rect 22637 11237 22649 11271
rect 22683 11268 22695 11271
rect 22726 11268 22732 11280
rect 22683 11240 22732 11268
rect 22683 11237 22695 11240
rect 22637 11231 22695 11237
rect 22726 11228 22732 11240
rect 22784 11228 22790 11280
rect 22836 11268 22864 11308
rect 23462 11296 23468 11308
rect 23520 11296 23526 11348
rect 24109 11339 24167 11345
rect 24109 11305 24121 11339
rect 24155 11305 24167 11339
rect 24109 11299 24167 11305
rect 24124 11268 24152 11299
rect 22836 11240 24152 11268
rect 24293 11203 24351 11209
rect 24293 11169 24305 11203
rect 24339 11169 24351 11203
rect 24474 11200 24480 11212
rect 24435 11172 24480 11200
rect 24293 11163 24351 11169
rect 22545 11135 22603 11141
rect 22545 11132 22557 11135
rect 21732 11104 22557 11132
rect 22545 11101 22557 11104
rect 22591 11132 22603 11135
rect 22634 11132 22640 11144
rect 22591 11104 22640 11132
rect 22591 11101 22603 11104
rect 22545 11095 22603 11101
rect 22634 11092 22640 11104
rect 22692 11092 22698 11144
rect 22910 11092 22916 11144
rect 22968 11132 22974 11144
rect 23005 11135 23063 11141
rect 23005 11132 23017 11135
rect 22968 11104 23017 11132
rect 22968 11092 22974 11104
rect 23005 11101 23017 11104
rect 23051 11101 23063 11135
rect 23005 11095 23063 11101
rect 11226 11073 11232 11076
rect 11210 11067 11232 11073
rect 11210 11064 11222 11067
rect 10968 11036 11222 11064
rect 11210 11033 11222 11036
rect 11284 11064 11290 11076
rect 11778 11064 11784 11076
rect 11284 11036 11784 11064
rect 11210 11027 11232 11033
rect 11226 11024 11232 11027
rect 11284 11024 11290 11036
rect 11778 11024 11784 11036
rect 11836 11024 11842 11076
rect 13894 11024 13900 11076
rect 13952 11064 13958 11076
rect 15093 11067 15151 11073
rect 15093 11064 15105 11067
rect 13952 11036 15105 11064
rect 13952 11024 13958 11036
rect 15093 11033 15105 11036
rect 15139 11064 15151 11067
rect 16102 11064 16108 11076
rect 15139 11036 16108 11064
rect 15139 11033 15151 11036
rect 15093 11027 15151 11033
rect 16102 11024 16108 11036
rect 16160 11024 16166 11076
rect 17853 11067 17911 11073
rect 17853 11033 17865 11067
rect 17899 11064 17911 11067
rect 18218 11064 18224 11076
rect 17899 11036 18224 11064
rect 17899 11033 17911 11036
rect 17853 11027 17911 11033
rect 18218 11024 18224 11036
rect 18276 11064 18282 11076
rect 19138 11064 19144 11076
rect 18276 11036 19000 11064
rect 19099 11036 19144 11064
rect 18276 11024 18282 11036
rect 11318 10996 11324 11008
rect 11279 10968 11324 10996
rect 11318 10956 11324 10968
rect 11376 10956 11382 11008
rect 14906 10956 14912 11008
rect 14964 11005 14970 11008
rect 14964 10999 15013 11005
rect 14964 10965 14967 10999
rect 15001 10965 15013 10999
rect 15274 10996 15280 11008
rect 15235 10968 15280 10996
rect 14964 10959 15013 10965
rect 14964 10956 14970 10959
rect 15274 10956 15280 10968
rect 15332 10956 15338 11008
rect 18494 10996 18500 11008
rect 18455 10968 18500 10996
rect 18494 10956 18500 10968
rect 18552 10956 18558 11008
rect 18678 10956 18684 11008
rect 18736 10996 18742 11008
rect 18972 11005 19000 11036
rect 19138 11024 19144 11036
rect 19196 11024 19202 11076
rect 24308 11064 24336 11163
rect 24474 11160 24480 11172
rect 24532 11160 24538 11212
rect 24308 11036 24428 11064
rect 24400 11008 24428 11036
rect 18819 10999 18877 11005
rect 18819 10996 18831 10999
rect 18736 10968 18831 10996
rect 18736 10956 18742 10968
rect 18819 10965 18831 10968
rect 18865 10965 18877 10999
rect 18819 10959 18877 10965
rect 18957 10999 19015 11005
rect 18957 10965 18969 10999
rect 19003 10996 19015 10999
rect 19414 10996 19420 11008
rect 19003 10968 19420 10996
rect 19003 10965 19015 10968
rect 18957 10959 19015 10965
rect 19414 10956 19420 10968
rect 19472 10956 19478 11008
rect 24382 10956 24388 11008
rect 24440 10956 24446 11008
rect 632 10906 26392 10928
rect 632 10854 5176 10906
rect 5228 10854 5240 10906
rect 5292 10854 5304 10906
rect 5356 10854 5368 10906
rect 5420 10854 14510 10906
rect 14562 10854 14574 10906
rect 14626 10854 14638 10906
rect 14690 10854 14702 10906
rect 14754 10854 23843 10906
rect 23895 10854 23907 10906
rect 23959 10854 23971 10906
rect 24023 10854 24035 10906
rect 24087 10854 26392 10906
rect 632 10832 26392 10854
rect 8098 10792 8104 10804
rect 8059 10764 8104 10792
rect 8098 10752 8104 10764
rect 8156 10752 8162 10804
rect 9662 10752 9668 10804
rect 9720 10792 9726 10804
rect 9849 10795 9907 10801
rect 9849 10792 9861 10795
rect 9720 10764 9861 10792
rect 9720 10752 9726 10764
rect 9849 10761 9861 10764
rect 9895 10761 9907 10795
rect 11318 10792 11324 10804
rect 11279 10764 11324 10792
rect 9849 10755 9907 10761
rect 11318 10752 11324 10764
rect 11376 10752 11382 10804
rect 11686 10792 11692 10804
rect 11647 10764 11692 10792
rect 11686 10752 11692 10764
rect 11744 10752 11750 10804
rect 13066 10792 13072 10804
rect 13027 10764 13072 10792
rect 13066 10752 13072 10764
rect 13124 10752 13130 10804
rect 13434 10792 13440 10804
rect 13395 10764 13440 10792
rect 13434 10752 13440 10764
rect 13492 10752 13498 10804
rect 13802 10792 13808 10804
rect 13763 10764 13808 10792
rect 13802 10752 13808 10764
rect 13860 10752 13866 10804
rect 14170 10801 14176 10804
rect 14154 10795 14176 10801
rect 14154 10792 14166 10795
rect 14083 10764 14166 10792
rect 14154 10761 14166 10764
rect 14228 10792 14234 10804
rect 14906 10792 14912 10804
rect 14228 10764 14912 10792
rect 14154 10755 14176 10761
rect 14170 10752 14176 10755
rect 14228 10752 14234 10764
rect 14906 10752 14912 10764
rect 14964 10752 14970 10804
rect 16102 10752 16108 10804
rect 16160 10792 16166 10804
rect 16565 10795 16623 10801
rect 16565 10792 16577 10795
rect 16160 10764 16577 10792
rect 16160 10752 16166 10764
rect 16565 10761 16577 10764
rect 16611 10792 16623 10795
rect 17298 10792 17304 10804
rect 16611 10764 17304 10792
rect 16611 10761 16623 10764
rect 16565 10755 16623 10761
rect 17298 10752 17304 10764
rect 17356 10752 17362 10804
rect 18678 10752 18684 10804
rect 18736 10792 18742 10804
rect 19279 10795 19337 10801
rect 19279 10792 19291 10795
rect 18736 10764 19291 10792
rect 18736 10752 18742 10764
rect 19279 10761 19291 10764
rect 19325 10792 19337 10795
rect 19506 10792 19512 10804
rect 19325 10764 19512 10792
rect 19325 10761 19337 10764
rect 19279 10755 19337 10761
rect 19506 10752 19512 10764
rect 19564 10792 19570 10804
rect 20153 10795 20211 10801
rect 20153 10792 20165 10795
rect 19564 10764 20165 10792
rect 19564 10752 19570 10764
rect 20153 10761 20165 10764
rect 20199 10761 20211 10795
rect 20153 10755 20211 10761
rect 21898 10752 21904 10804
rect 21956 10792 21962 10804
rect 22269 10795 22327 10801
rect 22269 10792 22281 10795
rect 21956 10764 22281 10792
rect 21956 10752 21962 10764
rect 22269 10761 22281 10764
rect 22315 10792 22327 10795
rect 22726 10792 22732 10804
rect 22315 10764 22732 10792
rect 22315 10761 22327 10764
rect 22269 10755 22327 10761
rect 22726 10752 22732 10764
rect 22784 10752 22790 10804
rect 24474 10752 24480 10804
rect 24532 10792 24538 10804
rect 24753 10795 24811 10801
rect 24753 10792 24765 10795
rect 24532 10764 24765 10792
rect 24532 10752 24538 10764
rect 24753 10761 24765 10764
rect 24799 10761 24811 10795
rect 24753 10755 24811 10761
rect 8466 10724 8472 10736
rect 8427 10696 8472 10724
rect 8466 10684 8472 10696
rect 8524 10684 8530 10736
rect 9205 10727 9263 10733
rect 9205 10693 9217 10727
rect 9251 10724 9263 10727
rect 9251 10696 12928 10724
rect 9251 10693 9263 10696
rect 9205 10687 9263 10693
rect 8285 10591 8343 10597
rect 8285 10557 8297 10591
rect 8331 10588 8343 10591
rect 9220 10588 9248 10687
rect 12057 10659 12115 10665
rect 12057 10625 12069 10659
rect 12103 10656 12115 10659
rect 12514 10656 12520 10668
rect 12103 10628 12520 10656
rect 12103 10625 12115 10628
rect 12057 10619 12115 10625
rect 12514 10616 12520 10628
rect 12572 10616 12578 10668
rect 9297 10591 9355 10597
rect 9297 10588 9309 10591
rect 8331 10560 8880 10588
rect 8331 10557 8343 10560
rect 8285 10551 8343 10557
rect 8852 10529 8880 10560
rect 9220 10560 9309 10588
rect 9220 10532 9248 10560
rect 9297 10557 9309 10560
rect 9343 10557 9355 10591
rect 10306 10588 10312 10600
rect 10267 10560 10312 10588
rect 9297 10551 9355 10557
rect 10306 10548 10312 10560
rect 10364 10548 10370 10600
rect 10766 10588 10772 10600
rect 10727 10560 10772 10588
rect 10766 10548 10772 10560
rect 10824 10548 10830 10600
rect 8837 10523 8895 10529
rect 8837 10489 8849 10523
rect 8883 10520 8895 10523
rect 9202 10520 9208 10532
rect 8883 10492 9208 10520
rect 8883 10489 8895 10492
rect 8837 10483 8895 10489
rect 9202 10480 9208 10492
rect 9260 10520 9266 10532
rect 11042 10520 11048 10532
rect 9260 10492 9353 10520
rect 11003 10492 11048 10520
rect 9260 10480 9266 10492
rect 11042 10480 11048 10492
rect 11100 10480 11106 10532
rect 11226 10480 11232 10532
rect 11284 10520 11290 10532
rect 12146 10520 12152 10532
rect 11284 10492 12152 10520
rect 11284 10480 11290 10492
rect 12146 10480 12152 10492
rect 12204 10480 12210 10532
rect 12701 10523 12759 10529
rect 12701 10489 12713 10523
rect 12747 10520 12759 10523
rect 12790 10520 12796 10532
rect 12747 10492 12796 10520
rect 12747 10489 12759 10492
rect 12701 10483 12759 10489
rect 12790 10480 12796 10492
rect 12848 10480 12854 10532
rect 12900 10520 12928 10696
rect 13820 10656 13848 10752
rect 13894 10684 13900 10736
rect 13952 10724 13958 10736
rect 14265 10727 14323 10733
rect 14265 10724 14277 10727
rect 13952 10696 14277 10724
rect 13952 10684 13958 10696
rect 14265 10693 14277 10696
rect 14311 10693 14323 10727
rect 19414 10724 19420 10736
rect 19327 10696 19420 10724
rect 14265 10687 14323 10693
rect 19414 10684 19420 10696
rect 19472 10724 19478 10736
rect 19690 10724 19696 10736
rect 19472 10696 19696 10724
rect 19472 10684 19478 10696
rect 19690 10684 19696 10696
rect 19748 10684 19754 10736
rect 21530 10684 21536 10736
rect 21588 10724 21594 10736
rect 22913 10727 22971 10733
rect 22913 10724 22925 10727
rect 21588 10696 22925 10724
rect 21588 10684 21594 10696
rect 22913 10693 22925 10696
rect 22959 10693 22971 10727
rect 24382 10724 24388 10736
rect 24343 10696 24388 10724
rect 22913 10687 22971 10693
rect 14357 10659 14415 10665
rect 14357 10656 14369 10659
rect 13820 10628 14369 10656
rect 14357 10625 14369 10628
rect 14403 10656 14415 10659
rect 15001 10659 15059 10665
rect 15001 10656 15013 10659
rect 14403 10628 15013 10656
rect 14403 10625 14415 10628
rect 14357 10619 14415 10625
rect 15001 10625 15013 10628
rect 15047 10656 15059 10659
rect 15182 10656 15188 10668
rect 15047 10628 15188 10656
rect 15047 10625 15059 10628
rect 15001 10619 15059 10625
rect 15182 10616 15188 10628
rect 15240 10656 15246 10668
rect 18681 10659 18739 10665
rect 18681 10656 18693 10659
rect 15240 10628 18693 10656
rect 15240 10616 15246 10628
rect 18681 10625 18693 10628
rect 18727 10656 18739 10659
rect 18954 10656 18960 10668
rect 18727 10628 18960 10656
rect 18727 10625 18739 10628
rect 18681 10619 18739 10625
rect 18954 10616 18960 10628
rect 19012 10656 19018 10668
rect 19509 10659 19567 10665
rect 19509 10656 19521 10659
rect 19012 10628 19521 10656
rect 19012 10616 19018 10628
rect 19509 10625 19521 10628
rect 19555 10625 19567 10659
rect 20610 10656 20616 10668
rect 20571 10628 20616 10656
rect 19509 10619 19567 10625
rect 20610 10616 20616 10628
rect 20668 10656 20674 10668
rect 21254 10656 21260 10668
rect 20668 10628 20748 10656
rect 21215 10628 21260 10656
rect 20668 10616 20674 10628
rect 13434 10548 13440 10600
rect 13492 10588 13498 10600
rect 13989 10591 14047 10597
rect 13989 10588 14001 10591
rect 13492 10560 14001 10588
rect 13492 10548 13498 10560
rect 13989 10557 14001 10560
rect 14035 10557 14047 10591
rect 13989 10551 14047 10557
rect 15645 10591 15703 10597
rect 15645 10557 15657 10591
rect 15691 10557 15703 10591
rect 17574 10588 17580 10600
rect 17535 10560 17580 10588
rect 15645 10551 15703 10557
rect 15553 10523 15611 10529
rect 15553 10520 15565 10523
rect 12900 10492 15565 10520
rect 15553 10489 15565 10492
rect 15599 10489 15611 10523
rect 15553 10483 15611 10489
rect 9478 10452 9484 10464
rect 9439 10424 9484 10452
rect 9478 10412 9484 10424
rect 9536 10412 9542 10464
rect 14630 10452 14636 10464
rect 14591 10424 14636 10452
rect 14630 10412 14636 10424
rect 14688 10412 14694 10464
rect 15366 10452 15372 10464
rect 15327 10424 15372 10452
rect 15366 10412 15372 10424
rect 15424 10452 15430 10464
rect 15660 10452 15688 10551
rect 17574 10548 17580 10560
rect 17632 10548 17638 10600
rect 18034 10588 18040 10600
rect 17995 10560 18040 10588
rect 18034 10548 18040 10560
rect 18092 10548 18098 10600
rect 20720 10597 20748 10628
rect 21254 10616 21260 10628
rect 21312 10616 21318 10668
rect 22928 10656 22956 10687
rect 24382 10684 24388 10696
rect 24440 10684 24446 10736
rect 22928 10628 23324 10656
rect 20705 10591 20763 10597
rect 20705 10557 20717 10591
rect 20751 10557 20763 10591
rect 20705 10551 20763 10557
rect 20886 10548 20892 10600
rect 20944 10588 20950 10600
rect 21165 10591 21223 10597
rect 21165 10588 21177 10591
rect 20944 10560 21177 10588
rect 20944 10548 20950 10560
rect 21165 10557 21177 10560
rect 21211 10588 21223 10591
rect 21717 10591 21775 10597
rect 21717 10588 21729 10591
rect 21211 10560 21729 10588
rect 21211 10557 21223 10560
rect 21165 10551 21223 10557
rect 21717 10557 21729 10560
rect 21763 10557 21775 10591
rect 21717 10551 21775 10557
rect 23189 10591 23247 10597
rect 23189 10557 23201 10591
rect 23235 10557 23247 10591
rect 23189 10551 23247 10557
rect 17206 10480 17212 10532
rect 17264 10520 17270 10532
rect 17301 10523 17359 10529
rect 17301 10520 17313 10523
rect 17264 10492 17313 10520
rect 17264 10480 17270 10492
rect 17301 10489 17313 10492
rect 17347 10520 17359 10523
rect 17482 10520 17488 10532
rect 17347 10492 17488 10520
rect 17347 10489 17359 10492
rect 17301 10483 17359 10489
rect 17482 10480 17488 10492
rect 17540 10480 17546 10532
rect 18310 10520 18316 10532
rect 18271 10492 18316 10520
rect 18310 10480 18316 10492
rect 18368 10480 18374 10532
rect 18494 10480 18500 10532
rect 18552 10520 18558 10532
rect 19141 10523 19199 10529
rect 19141 10520 19153 10523
rect 18552 10492 19153 10520
rect 18552 10480 18558 10492
rect 19141 10489 19153 10492
rect 19187 10489 19199 10523
rect 19874 10520 19880 10532
rect 19835 10492 19880 10520
rect 19141 10483 19199 10489
rect 19874 10480 19880 10492
rect 19932 10480 19938 10532
rect 22542 10520 22548 10532
rect 22503 10492 22548 10520
rect 22542 10480 22548 10492
rect 22600 10520 22606 10532
rect 23204 10520 23232 10551
rect 22600 10492 23232 10520
rect 23296 10520 23324 10628
rect 24934 10588 24940 10600
rect 24895 10560 24940 10588
rect 24934 10548 24940 10560
rect 24992 10588 24998 10600
rect 25489 10591 25547 10597
rect 25489 10588 25501 10591
rect 24992 10560 25501 10588
rect 24992 10548 24998 10560
rect 25489 10557 25501 10560
rect 25535 10557 25547 10591
rect 25489 10551 25547 10557
rect 23510 10523 23568 10529
rect 23510 10520 23522 10523
rect 23296 10492 23522 10520
rect 22600 10480 22606 10492
rect 23510 10489 23522 10492
rect 23556 10489 23568 10523
rect 23510 10483 23568 10489
rect 15424 10424 15688 10452
rect 15424 10412 15430 10424
rect 16654 10412 16660 10464
rect 16712 10452 16718 10464
rect 16930 10452 16936 10464
rect 16712 10424 16936 10452
rect 16712 10412 16718 10424
rect 16930 10412 16936 10424
rect 16988 10412 16994 10464
rect 24106 10452 24112 10464
rect 24067 10424 24112 10452
rect 24106 10412 24112 10424
rect 24164 10412 24170 10464
rect 24474 10412 24480 10464
rect 24532 10452 24538 10464
rect 25121 10455 25179 10461
rect 25121 10452 25133 10455
rect 24532 10424 25133 10452
rect 24532 10412 24538 10424
rect 25121 10421 25133 10424
rect 25167 10421 25179 10455
rect 25121 10415 25179 10421
rect 632 10362 26392 10384
rect 632 10310 9843 10362
rect 9895 10310 9907 10362
rect 9959 10310 9971 10362
rect 10023 10310 10035 10362
rect 10087 10310 19176 10362
rect 19228 10310 19240 10362
rect 19292 10310 19304 10362
rect 19356 10310 19368 10362
rect 19420 10310 26392 10362
rect 632 10288 26392 10310
rect 9849 10251 9907 10257
rect 9849 10217 9861 10251
rect 9895 10248 9907 10251
rect 10766 10248 10772 10260
rect 9895 10220 10772 10248
rect 9895 10217 9907 10220
rect 9849 10211 9907 10217
rect 10766 10208 10772 10220
rect 10824 10208 10830 10260
rect 11226 10248 11232 10260
rect 11187 10220 11232 10248
rect 11226 10208 11232 10220
rect 11284 10208 11290 10260
rect 11410 10208 11416 10260
rect 11468 10248 11474 10260
rect 11505 10251 11563 10257
rect 11505 10248 11517 10251
rect 11468 10220 11517 10248
rect 11468 10208 11474 10220
rect 11505 10217 11517 10220
rect 11551 10217 11563 10251
rect 11505 10211 11563 10217
rect 12054 10208 12060 10260
rect 12112 10208 12118 10260
rect 12146 10208 12152 10260
rect 12204 10248 12210 10260
rect 13069 10251 13127 10257
rect 13069 10248 13081 10251
rect 12204 10220 13081 10248
rect 12204 10208 12210 10220
rect 13069 10217 13081 10220
rect 13115 10217 13127 10251
rect 13069 10211 13127 10217
rect 13253 10251 13311 10257
rect 13253 10217 13265 10251
rect 13299 10248 13311 10251
rect 14170 10248 14176 10260
rect 13299 10220 14176 10248
rect 13299 10217 13311 10220
rect 13253 10211 13311 10217
rect 14170 10208 14176 10220
rect 14228 10208 14234 10260
rect 14354 10208 14360 10260
rect 14412 10248 14418 10260
rect 14541 10251 14599 10257
rect 14541 10248 14553 10251
rect 14412 10220 14553 10248
rect 14412 10208 14418 10220
rect 14541 10217 14553 10220
rect 14587 10217 14599 10251
rect 16194 10248 16200 10260
rect 16155 10220 16200 10248
rect 14541 10211 14599 10217
rect 16194 10208 16200 10220
rect 16252 10208 16258 10260
rect 17574 10248 17580 10260
rect 17535 10220 17580 10248
rect 17574 10208 17580 10220
rect 17632 10208 17638 10260
rect 18954 10208 18960 10260
rect 19012 10248 19018 10260
rect 19141 10251 19199 10257
rect 19141 10248 19153 10251
rect 19012 10220 19153 10248
rect 19012 10208 19018 10220
rect 19141 10217 19153 10220
rect 19187 10217 19199 10251
rect 19506 10248 19512 10260
rect 19467 10220 19512 10248
rect 19141 10211 19199 10217
rect 19506 10208 19512 10220
rect 19564 10208 19570 10260
rect 19690 10208 19696 10260
rect 19748 10248 19754 10260
rect 19877 10251 19935 10257
rect 19877 10248 19889 10251
rect 19748 10220 19889 10248
rect 19748 10208 19754 10220
rect 19877 10217 19889 10220
rect 19923 10217 19935 10251
rect 19877 10211 19935 10217
rect 20150 10208 20156 10260
rect 20208 10248 20214 10260
rect 20426 10248 20432 10260
rect 20208 10220 20432 10248
rect 20208 10208 20214 10220
rect 20426 10208 20432 10220
rect 20484 10248 20490 10260
rect 20613 10251 20671 10257
rect 20613 10248 20625 10251
rect 20484 10220 20625 10248
rect 20484 10208 20490 10220
rect 20613 10217 20625 10220
rect 20659 10217 20671 10251
rect 21898 10248 21904 10260
rect 21859 10220 21904 10248
rect 20613 10211 20671 10217
rect 21898 10208 21904 10220
rect 21956 10208 21962 10260
rect 22545 10251 22603 10257
rect 22545 10217 22557 10251
rect 22591 10248 22603 10251
rect 22634 10248 22640 10260
rect 22591 10220 22640 10248
rect 22591 10217 22603 10220
rect 22545 10211 22603 10217
rect 22634 10208 22640 10220
rect 22692 10208 22698 10260
rect 10674 10189 10680 10192
rect 10671 10180 10680 10189
rect 10635 10152 10680 10180
rect 10671 10143 10680 10152
rect 10674 10140 10680 10143
rect 10732 10140 10738 10192
rect 12072 10180 12100 10208
rect 12241 10183 12299 10189
rect 12241 10180 12253 10183
rect 12072 10152 12253 10180
rect 12241 10149 12253 10152
rect 12287 10149 12299 10183
rect 12241 10143 12299 10149
rect 16286 10140 16292 10192
rect 16344 10180 16350 10192
rect 16746 10189 16752 10192
rect 16743 10180 16752 10189
rect 16344 10152 16752 10180
rect 16344 10140 16350 10152
rect 16743 10143 16752 10152
rect 16746 10140 16752 10143
rect 16804 10140 16810 10192
rect 18494 10180 18500 10192
rect 18144 10152 18500 10180
rect 9202 10072 9208 10124
rect 9260 10112 9266 10124
rect 9297 10115 9355 10121
rect 9297 10112 9309 10115
rect 9260 10084 9309 10112
rect 9260 10072 9266 10084
rect 9297 10081 9309 10084
rect 9343 10081 9355 10115
rect 9297 10075 9355 10081
rect 10309 10115 10367 10121
rect 10309 10081 10321 10115
rect 10355 10112 10367 10115
rect 10490 10112 10496 10124
rect 10355 10084 10496 10112
rect 10355 10081 10367 10084
rect 10309 10075 10367 10081
rect 10490 10072 10496 10084
rect 10548 10072 10554 10124
rect 13526 10072 13532 10124
rect 13584 10112 13590 10124
rect 13621 10115 13679 10121
rect 13621 10112 13633 10115
rect 13584 10084 13633 10112
rect 13584 10072 13590 10084
rect 13621 10081 13633 10084
rect 13667 10081 13679 10115
rect 13621 10075 13679 10081
rect 13986 10072 13992 10124
rect 14044 10112 14050 10124
rect 14817 10115 14875 10121
rect 14817 10112 14829 10115
rect 14044 10084 14829 10112
rect 14044 10072 14050 10084
rect 14817 10081 14829 10084
rect 14863 10081 14875 10115
rect 14817 10075 14875 10081
rect 9478 10004 9484 10056
rect 9536 10044 9542 10056
rect 10398 10044 10404 10056
rect 9536 10016 10404 10044
rect 9536 10004 9542 10016
rect 10398 10004 10404 10016
rect 10456 10004 10462 10056
rect 12149 10047 12207 10053
rect 12149 10013 12161 10047
rect 12195 10044 12207 10047
rect 12790 10044 12796 10056
rect 12195 10016 12796 10044
rect 12195 10013 12207 10016
rect 12149 10007 12207 10013
rect 12790 10004 12796 10016
rect 12848 10004 12854 10056
rect 12698 9976 12704 9988
rect 12659 9948 12704 9976
rect 12698 9936 12704 9948
rect 12756 9936 12762 9988
rect 13529 9979 13587 9985
rect 13529 9945 13541 9979
rect 13575 9976 13587 9979
rect 13894 9976 13900 9988
rect 13575 9948 13900 9976
rect 13575 9945 13587 9948
rect 13529 9939 13587 9945
rect 13894 9936 13900 9948
rect 13952 9936 13958 9988
rect 14832 9976 14860 10075
rect 14906 10072 14912 10124
rect 14964 10112 14970 10124
rect 15274 10112 15280 10124
rect 14964 10084 15280 10112
rect 14964 10072 14970 10084
rect 15274 10072 15280 10084
rect 15332 10072 15338 10124
rect 16381 10115 16439 10121
rect 16381 10081 16393 10115
rect 16427 10112 16439 10115
rect 16470 10112 16476 10124
rect 16427 10084 16476 10112
rect 16427 10081 16439 10084
rect 16381 10075 16439 10081
rect 16470 10072 16476 10084
rect 16528 10072 16534 10124
rect 18144 10121 18172 10152
rect 18494 10140 18500 10152
rect 18552 10140 18558 10192
rect 21343 10183 21401 10189
rect 21343 10149 21355 10183
rect 21389 10180 21401 10183
rect 21530 10180 21536 10192
rect 21389 10152 21536 10180
rect 21389 10149 21401 10152
rect 21343 10143 21401 10149
rect 21530 10140 21536 10152
rect 21588 10140 21594 10192
rect 24106 10140 24112 10192
rect 24164 10180 24170 10192
rect 24201 10183 24259 10189
rect 24201 10180 24213 10183
rect 24164 10152 24213 10180
rect 24164 10140 24170 10152
rect 24201 10149 24213 10152
rect 24247 10149 24259 10183
rect 24201 10143 24259 10149
rect 18129 10115 18187 10121
rect 18129 10112 18141 10115
rect 17960 10084 18141 10112
rect 15553 10047 15611 10053
rect 15553 10013 15565 10047
rect 15599 10044 15611 10047
rect 16010 10044 16016 10056
rect 15599 10016 16016 10044
rect 15599 10013 15611 10016
rect 15553 10007 15611 10013
rect 16010 10004 16016 10016
rect 16068 10004 16074 10056
rect 16930 9976 16936 9988
rect 14832 9948 16936 9976
rect 9481 9911 9539 9917
rect 9481 9877 9493 9911
rect 9527 9908 9539 9911
rect 10125 9911 10183 9917
rect 10125 9908 10137 9911
rect 9527 9880 10137 9908
rect 9527 9877 9539 9880
rect 9481 9871 9539 9877
rect 10125 9877 10137 9880
rect 10171 9908 10183 9911
rect 10306 9908 10312 9920
rect 10171 9880 10312 9908
rect 10171 9877 10183 9880
rect 10125 9871 10183 9877
rect 10306 9868 10312 9880
rect 10364 9868 10370 9920
rect 11778 9868 11784 9920
rect 11836 9908 11842 9920
rect 11965 9911 12023 9917
rect 11965 9908 11977 9911
rect 11836 9880 11977 9908
rect 11836 9868 11842 9880
rect 11965 9877 11977 9880
rect 12011 9908 12023 9911
rect 13253 9911 13311 9917
rect 13253 9908 13265 9911
rect 12011 9880 13265 9908
rect 12011 9877 12023 9880
rect 11965 9871 12023 9877
rect 13253 9877 13265 9880
rect 13299 9877 13311 9911
rect 13802 9908 13808 9920
rect 13763 9880 13808 9908
rect 13253 9871 13311 9877
rect 13802 9868 13808 9880
rect 13860 9868 13866 9920
rect 14832 9908 14860 9948
rect 16930 9936 16936 9948
rect 16988 9936 16994 9988
rect 14906 9908 14912 9920
rect 14832 9880 14912 9908
rect 14906 9868 14912 9880
rect 14964 9868 14970 9920
rect 15826 9908 15832 9920
rect 15787 9880 15832 9908
rect 15826 9868 15832 9880
rect 15884 9868 15890 9920
rect 17301 9911 17359 9917
rect 17301 9877 17313 9911
rect 17347 9908 17359 9911
rect 17390 9908 17396 9920
rect 17347 9880 17396 9908
rect 17347 9877 17359 9880
rect 17301 9871 17359 9877
rect 17390 9868 17396 9880
rect 17448 9868 17454 9920
rect 17850 9868 17856 9920
rect 17908 9908 17914 9920
rect 17960 9917 17988 10084
rect 18129 10081 18141 10084
rect 18175 10081 18187 10115
rect 18129 10075 18187 10081
rect 18276 10115 18334 10121
rect 18276 10081 18288 10115
rect 18322 10112 18334 10115
rect 18678 10112 18684 10124
rect 18322 10084 18684 10112
rect 18322 10081 18334 10084
rect 18276 10075 18334 10081
rect 18678 10072 18684 10084
rect 18736 10072 18742 10124
rect 20978 10112 20984 10124
rect 20939 10084 20984 10112
rect 20978 10072 20984 10084
rect 21036 10112 21042 10124
rect 21622 10112 21628 10124
rect 21036 10084 21628 10112
rect 21036 10072 21042 10084
rect 21622 10072 21628 10084
rect 21680 10072 21686 10124
rect 23072 10115 23130 10121
rect 23072 10081 23084 10115
rect 23118 10112 23130 10115
rect 23462 10112 23468 10124
rect 23118 10084 23468 10112
rect 23118 10081 23130 10084
rect 23072 10075 23130 10081
rect 23462 10072 23468 10084
rect 23520 10072 23526 10124
rect 18497 10047 18555 10053
rect 18497 10013 18509 10047
rect 18543 10044 18555 10047
rect 18954 10044 18960 10056
rect 18543 10016 18960 10044
rect 18543 10013 18555 10016
rect 18497 10007 18555 10013
rect 18954 10004 18960 10016
rect 19012 10004 19018 10056
rect 22082 10004 22088 10056
rect 22140 10044 22146 10056
rect 24109 10047 24167 10053
rect 24109 10044 24121 10047
rect 22140 10016 24121 10044
rect 22140 10004 22146 10016
rect 24109 10013 24121 10016
rect 24155 10044 24167 10047
rect 24566 10044 24572 10056
rect 24155 10016 24572 10044
rect 24155 10013 24167 10016
rect 24109 10007 24167 10013
rect 24566 10004 24572 10016
rect 24624 10004 24630 10056
rect 24750 10044 24756 10056
rect 24711 10016 24756 10044
rect 24750 10004 24756 10016
rect 24808 10004 24814 10056
rect 17945 9911 18003 9917
rect 17945 9908 17957 9911
rect 17908 9880 17957 9908
rect 17908 9868 17914 9880
rect 17945 9877 17957 9880
rect 17991 9877 18003 9911
rect 18402 9908 18408 9920
rect 18363 9880 18408 9908
rect 17945 9871 18003 9877
rect 18402 9868 18408 9880
rect 18460 9868 18466 9920
rect 18586 9908 18592 9920
rect 18547 9880 18592 9908
rect 18586 9868 18592 9880
rect 18644 9868 18650 9920
rect 23143 9911 23201 9917
rect 23143 9877 23155 9911
rect 23189 9908 23201 9911
rect 23554 9908 23560 9920
rect 23189 9880 23560 9908
rect 23189 9877 23201 9880
rect 23143 9871 23201 9877
rect 23554 9868 23560 9880
rect 23612 9868 23618 9920
rect 632 9818 26392 9840
rect 632 9766 5176 9818
rect 5228 9766 5240 9818
rect 5292 9766 5304 9818
rect 5356 9766 5368 9818
rect 5420 9766 14510 9818
rect 14562 9766 14574 9818
rect 14626 9766 14638 9818
rect 14690 9766 14702 9818
rect 14754 9766 23843 9818
rect 23895 9766 23907 9818
rect 23959 9766 23971 9818
rect 24023 9766 24035 9818
rect 24087 9766 26392 9818
rect 632 9744 26392 9766
rect 7270 9664 7276 9716
rect 7328 9704 7334 9716
rect 8190 9704 8196 9716
rect 7328 9676 8196 9704
rect 7328 9664 7334 9676
rect 8190 9664 8196 9676
rect 8248 9664 8254 9716
rect 9021 9707 9079 9713
rect 9021 9673 9033 9707
rect 9067 9704 9079 9707
rect 9202 9704 9208 9716
rect 9067 9676 9208 9704
rect 9067 9673 9079 9676
rect 9021 9667 9079 9673
rect 9202 9664 9208 9676
rect 9260 9664 9266 9716
rect 11226 9704 11232 9716
rect 10508 9676 11232 9704
rect 9478 9596 9484 9648
rect 9536 9596 9542 9648
rect 10214 9596 10220 9648
rect 10272 9636 10278 9648
rect 10508 9636 10536 9676
rect 11226 9664 11232 9676
rect 11284 9664 11290 9716
rect 13526 9704 13532 9716
rect 13268 9676 13532 9704
rect 10272 9608 10536 9636
rect 10272 9596 10278 9608
rect 10582 9596 10588 9648
rect 10640 9636 10646 9648
rect 11321 9639 11379 9645
rect 11321 9636 11333 9639
rect 10640 9608 11333 9636
rect 10640 9596 10646 9608
rect 11321 9605 11333 9608
rect 11367 9605 11379 9639
rect 11321 9599 11379 9605
rect 11781 9639 11839 9645
rect 11781 9605 11793 9639
rect 11827 9636 11839 9639
rect 12054 9636 12060 9648
rect 11827 9608 12060 9636
rect 11827 9605 11839 9608
rect 11781 9599 11839 9605
rect 12054 9596 12060 9608
rect 12112 9596 12118 9648
rect 12977 9639 13035 9645
rect 12977 9605 12989 9639
rect 13023 9636 13035 9639
rect 13268 9636 13296 9676
rect 13526 9664 13532 9676
rect 13584 9664 13590 9716
rect 14906 9704 14912 9716
rect 14867 9676 14912 9704
rect 14906 9664 14912 9676
rect 14964 9664 14970 9716
rect 14998 9664 15004 9716
rect 15056 9704 15062 9716
rect 15185 9707 15243 9713
rect 15185 9704 15197 9707
rect 15056 9676 15197 9704
rect 15056 9664 15062 9676
rect 15185 9673 15197 9676
rect 15231 9673 15243 9707
rect 17298 9704 17304 9716
rect 17259 9676 17304 9704
rect 15185 9667 15243 9673
rect 17298 9664 17304 9676
rect 17356 9704 17362 9716
rect 18402 9704 18408 9716
rect 17356 9676 18408 9704
rect 17356 9664 17362 9676
rect 18402 9664 18408 9676
rect 18460 9704 18466 9716
rect 18681 9707 18739 9713
rect 18460 9676 18632 9704
rect 18460 9664 18466 9676
rect 13023 9608 13296 9636
rect 13023 9605 13035 9608
rect 12977 9599 13035 9605
rect 15918 9596 15924 9648
rect 15976 9636 15982 9648
rect 16013 9639 16071 9645
rect 16013 9636 16025 9639
rect 15976 9608 16025 9636
rect 15976 9596 15982 9608
rect 16013 9605 16025 9608
rect 16059 9605 16071 9639
rect 18604 9636 18632 9676
rect 18681 9673 18693 9707
rect 18727 9704 18739 9707
rect 18954 9704 18960 9716
rect 18727 9676 18960 9704
rect 18727 9673 18739 9676
rect 18681 9667 18739 9673
rect 18954 9664 18960 9676
rect 19012 9664 19018 9716
rect 19306 9707 19364 9713
rect 19306 9673 19318 9707
rect 19352 9704 19364 9707
rect 19506 9704 19512 9716
rect 19352 9676 19512 9704
rect 19352 9673 19364 9676
rect 19306 9667 19364 9673
rect 19506 9664 19512 9676
rect 19564 9704 19570 9716
rect 20153 9707 20211 9713
rect 20153 9704 20165 9707
rect 19564 9676 20165 9704
rect 19564 9664 19570 9676
rect 20153 9673 20165 9676
rect 20199 9673 20211 9707
rect 20153 9667 20211 9673
rect 21622 9664 21628 9716
rect 21680 9664 21686 9716
rect 21806 9664 21812 9716
rect 21864 9704 21870 9716
rect 22174 9704 22180 9716
rect 21864 9676 22180 9704
rect 21864 9664 21870 9676
rect 22174 9664 22180 9676
rect 22232 9664 22238 9716
rect 18604 9608 18908 9636
rect 16013 9599 16071 9605
rect 9294 9528 9300 9580
rect 9352 9568 9358 9580
rect 9496 9568 9524 9596
rect 9352 9540 9524 9568
rect 10125 9571 10183 9577
rect 9352 9528 9358 9540
rect 10125 9537 10137 9571
rect 10171 9568 10183 9571
rect 10674 9568 10680 9580
rect 10171 9540 10680 9568
rect 10171 9537 10183 9540
rect 10125 9531 10183 9537
rect 10674 9528 10680 9540
rect 10732 9528 10738 9580
rect 11045 9571 11103 9577
rect 11045 9537 11057 9571
rect 11091 9568 11103 9571
rect 12790 9568 12796 9580
rect 11091 9540 12796 9568
rect 11091 9537 11103 9540
rect 11045 9531 11103 9537
rect 12790 9528 12796 9540
rect 12848 9528 12854 9580
rect 15461 9571 15519 9577
rect 15461 9537 15473 9571
rect 15507 9568 15519 9571
rect 16838 9568 16844 9580
rect 15507 9540 16844 9568
rect 15507 9537 15519 9540
rect 15461 9531 15519 9537
rect 16838 9528 16844 9540
rect 16896 9528 16902 9580
rect 17666 9568 17672 9580
rect 17627 9540 17672 9568
rect 17666 9528 17672 9540
rect 17724 9528 17730 9580
rect 9164 9503 9222 9509
rect 9164 9469 9176 9503
rect 9210 9500 9222 9503
rect 9478 9500 9484 9512
rect 9210 9472 9484 9500
rect 9210 9469 9222 9472
rect 9164 9463 9222 9469
rect 9478 9460 9484 9472
rect 9536 9500 9542 9512
rect 9573 9503 9631 9509
rect 9573 9500 9585 9503
rect 9536 9472 9585 9500
rect 9536 9460 9542 9472
rect 9573 9469 9585 9472
rect 9619 9469 9631 9503
rect 9573 9463 9631 9469
rect 13345 9503 13403 9509
rect 13345 9469 13357 9503
rect 13391 9500 13403 9503
rect 13710 9500 13716 9512
rect 13391 9472 13716 9500
rect 13391 9469 13403 9472
rect 13345 9463 13403 9469
rect 13710 9460 13716 9472
rect 13768 9460 13774 9512
rect 13897 9503 13955 9509
rect 13897 9469 13909 9503
rect 13943 9469 13955 9503
rect 13897 9463 13955 9469
rect 9251 9435 9309 9441
rect 9251 9401 9263 9435
rect 9297 9432 9309 9435
rect 10398 9432 10404 9444
rect 9297 9404 10404 9432
rect 9297 9401 9309 9404
rect 9251 9395 9309 9401
rect 10398 9392 10404 9404
rect 10456 9392 10462 9444
rect 10490 9392 10496 9444
rect 10548 9432 10554 9444
rect 12609 9435 12667 9441
rect 10548 9404 10593 9432
rect 10548 9392 10554 9404
rect 12609 9401 12621 9435
rect 12655 9432 12667 9435
rect 13802 9432 13808 9444
rect 12655 9404 13808 9432
rect 12655 9401 12667 9404
rect 12609 9395 12667 9401
rect 13802 9392 13808 9404
rect 13860 9432 13866 9444
rect 13912 9432 13940 9463
rect 13986 9460 13992 9512
rect 14044 9500 14050 9512
rect 14265 9503 14323 9509
rect 14265 9500 14277 9503
rect 14044 9472 14277 9500
rect 14044 9460 14050 9472
rect 14265 9469 14277 9472
rect 14311 9469 14323 9503
rect 18880 9500 18908 9608
rect 18972 9568 19000 9664
rect 20794 9636 20800 9648
rect 20707 9608 20800 9636
rect 20794 9596 20800 9608
rect 20852 9636 20858 9648
rect 21073 9639 21131 9645
rect 21073 9636 21085 9639
rect 20852 9608 21085 9636
rect 20852 9596 20858 9608
rect 21073 9605 21085 9608
rect 21119 9636 21131 9639
rect 21530 9636 21536 9648
rect 21119 9608 21536 9636
rect 21119 9605 21131 9608
rect 21073 9599 21131 9605
rect 21530 9596 21536 9608
rect 21588 9596 21594 9648
rect 21640 9636 21668 9664
rect 22453 9639 22511 9645
rect 22453 9636 22465 9639
rect 21640 9608 22465 9636
rect 22453 9605 22465 9608
rect 22499 9605 22511 9639
rect 22453 9599 22511 9605
rect 19509 9571 19567 9577
rect 19509 9568 19521 9571
rect 18972 9540 19521 9568
rect 19509 9537 19521 9540
rect 19555 9537 19567 9571
rect 21254 9568 21260 9580
rect 21215 9540 21260 9568
rect 19509 9531 19567 9537
rect 21254 9528 21260 9540
rect 21312 9568 21318 9580
rect 22821 9571 22879 9577
rect 22821 9568 22833 9571
rect 21312 9540 22833 9568
rect 21312 9528 21318 9540
rect 22821 9537 22833 9540
rect 22867 9537 22879 9571
rect 25489 9571 25547 9577
rect 25489 9568 25501 9571
rect 22821 9531 22879 9537
rect 24032 9540 25501 9568
rect 18954 9500 18960 9512
rect 18867 9472 18960 9500
rect 14265 9463 14323 9469
rect 18954 9460 18960 9472
rect 19012 9500 19018 9512
rect 19371 9503 19429 9509
rect 19371 9500 19383 9503
rect 19012 9472 19383 9500
rect 19012 9460 19018 9472
rect 19371 9469 19383 9472
rect 19417 9469 19429 9503
rect 19371 9463 19429 9469
rect 22177 9503 22235 9509
rect 22177 9469 22189 9503
rect 22223 9500 22235 9503
rect 22634 9500 22640 9512
rect 22223 9472 22640 9500
rect 22223 9469 22235 9472
rect 22177 9463 22235 9469
rect 22634 9460 22640 9472
rect 22692 9500 22698 9512
rect 23370 9500 23376 9512
rect 22692 9472 23376 9500
rect 22692 9460 22698 9472
rect 23370 9460 23376 9472
rect 23428 9460 23434 9512
rect 13860 9404 13940 9432
rect 15553 9435 15611 9441
rect 13860 9392 13866 9404
rect 15553 9401 15565 9435
rect 15599 9432 15611 9435
rect 15826 9432 15832 9444
rect 15599 9404 15832 9432
rect 15599 9401 15611 9404
rect 15553 9395 15611 9401
rect 15826 9392 15832 9404
rect 15884 9392 15890 9444
rect 17025 9435 17083 9441
rect 17025 9401 17037 9435
rect 17071 9432 17083 9435
rect 17390 9432 17396 9444
rect 17071 9404 17396 9432
rect 17071 9401 17083 9404
rect 17025 9395 17083 9401
rect 17390 9392 17396 9404
rect 17448 9432 17454 9444
rect 17761 9435 17819 9441
rect 17448 9404 17620 9432
rect 17448 9392 17454 9404
rect 11962 9324 11968 9376
rect 12020 9364 12026 9376
rect 14541 9367 14599 9373
rect 12020 9336 12065 9364
rect 12020 9324 12026 9336
rect 14541 9333 14553 9367
rect 14587 9364 14599 9367
rect 14722 9364 14728 9376
rect 14587 9336 14728 9364
rect 14587 9333 14599 9336
rect 14541 9327 14599 9333
rect 14722 9324 14728 9336
rect 14780 9324 14786 9376
rect 16473 9367 16531 9373
rect 16473 9333 16485 9367
rect 16519 9364 16531 9367
rect 16746 9364 16752 9376
rect 16519 9336 16752 9364
rect 16519 9333 16531 9336
rect 16473 9327 16531 9333
rect 16746 9324 16752 9336
rect 16804 9324 16810 9376
rect 17592 9364 17620 9404
rect 17761 9401 17773 9435
rect 17807 9401 17819 9435
rect 17761 9395 17819 9401
rect 17776 9364 17804 9395
rect 17850 9392 17856 9444
rect 17908 9432 17914 9444
rect 18313 9435 18371 9441
rect 18313 9432 18325 9435
rect 17908 9404 18325 9432
rect 17908 9392 17914 9404
rect 18313 9401 18325 9404
rect 18359 9401 18371 9435
rect 18313 9395 18371 9401
rect 18862 9392 18868 9444
rect 18920 9432 18926 9444
rect 19141 9435 19199 9441
rect 19141 9432 19153 9435
rect 18920 9404 19153 9432
rect 18920 9392 18926 9404
rect 19141 9401 19153 9404
rect 19187 9401 19199 9435
rect 19141 9395 19199 9401
rect 21530 9392 21536 9444
rect 21588 9441 21594 9444
rect 21588 9435 21636 9441
rect 21588 9401 21590 9435
rect 21624 9401 21636 9435
rect 21588 9395 21636 9401
rect 21588 9392 21594 9395
rect 23922 9392 23928 9444
rect 23980 9432 23986 9444
rect 24032 9432 24060 9540
rect 25489 9537 25501 9540
rect 25535 9537 25547 9571
rect 25489 9531 25547 9537
rect 24842 9460 24848 9512
rect 24900 9500 24906 9512
rect 24900 9472 24945 9500
rect 24900 9460 24906 9472
rect 24201 9435 24259 9441
rect 24201 9432 24213 9435
rect 23980 9404 24213 9432
rect 23980 9392 23986 9404
rect 24201 9401 24213 9404
rect 24247 9401 24259 9435
rect 24201 9395 24259 9401
rect 24290 9392 24296 9444
rect 24348 9432 24354 9444
rect 24348 9404 24393 9432
rect 24348 9392 24354 9404
rect 24566 9392 24572 9444
rect 24624 9432 24630 9444
rect 25121 9435 25179 9441
rect 25121 9432 25133 9435
rect 24624 9404 25133 9432
rect 24624 9392 24630 9404
rect 25121 9401 25133 9404
rect 25167 9401 25179 9435
rect 25121 9395 25179 9401
rect 18402 9364 18408 9376
rect 17592 9336 18408 9364
rect 18402 9324 18408 9336
rect 18460 9324 18466 9376
rect 19782 9364 19788 9376
rect 19743 9336 19788 9364
rect 19782 9324 19788 9336
rect 19840 9324 19846 9376
rect 23462 9364 23468 9376
rect 23423 9336 23468 9364
rect 23462 9324 23468 9336
rect 23520 9324 23526 9376
rect 24017 9367 24075 9373
rect 24017 9333 24029 9367
rect 24063 9364 24075 9367
rect 24308 9364 24336 9392
rect 24063 9336 24336 9364
rect 24063 9333 24075 9336
rect 24017 9327 24075 9333
rect 632 9274 26392 9296
rect 632 9222 9843 9274
rect 9895 9222 9907 9274
rect 9959 9222 9971 9274
rect 10023 9222 10035 9274
rect 10087 9222 19176 9274
rect 19228 9222 19240 9274
rect 19292 9222 19304 9274
rect 19356 9222 19368 9274
rect 19420 9222 26392 9274
rect 632 9200 26392 9222
rect 10398 9120 10404 9172
rect 10456 9160 10462 9172
rect 10953 9163 11011 9169
rect 10953 9160 10965 9163
rect 10456 9132 10965 9160
rect 10456 9120 10462 9132
rect 10953 9129 10965 9132
rect 10999 9129 11011 9163
rect 12054 9160 12060 9172
rect 12015 9132 12060 9160
rect 10953 9123 11011 9129
rect 12054 9120 12060 9132
rect 12112 9120 12118 9172
rect 12425 9163 12483 9169
rect 12425 9129 12437 9163
rect 12471 9160 12483 9163
rect 12514 9160 12520 9172
rect 12471 9132 12520 9160
rect 12471 9129 12483 9132
rect 12425 9123 12483 9129
rect 12514 9120 12520 9132
rect 12572 9120 12578 9172
rect 12790 9160 12796 9172
rect 12751 9132 12796 9160
rect 12790 9120 12796 9132
rect 12848 9120 12854 9172
rect 14630 9160 14636 9172
rect 14591 9132 14636 9160
rect 14630 9120 14636 9132
rect 14688 9120 14694 9172
rect 16470 9160 16476 9172
rect 16431 9132 16476 9160
rect 16470 9120 16476 9132
rect 16528 9120 16534 9172
rect 18589 9163 18647 9169
rect 18589 9129 18601 9163
rect 18635 9160 18647 9163
rect 18678 9160 18684 9172
rect 18635 9132 18684 9160
rect 18635 9129 18647 9132
rect 18589 9123 18647 9129
rect 18678 9120 18684 9132
rect 18736 9120 18742 9172
rect 18954 9120 18960 9172
rect 19012 9160 19018 9172
rect 19141 9163 19199 9169
rect 19141 9160 19153 9163
rect 19012 9132 19153 9160
rect 19012 9120 19018 9132
rect 19141 9129 19153 9132
rect 19187 9129 19199 9163
rect 19141 9123 19199 9129
rect 19463 9163 19521 9169
rect 19463 9129 19475 9163
rect 19509 9160 19521 9163
rect 19598 9160 19604 9172
rect 19509 9132 19604 9160
rect 19509 9129 19521 9132
rect 19463 9123 19521 9129
rect 19598 9120 19604 9132
rect 19656 9120 19662 9172
rect 20978 9120 20984 9172
rect 21036 9160 21042 9172
rect 21346 9160 21352 9172
rect 21036 9132 21352 9160
rect 21036 9120 21042 9132
rect 21346 9120 21352 9132
rect 21404 9120 21410 9172
rect 24109 9163 24167 9169
rect 24109 9129 24121 9163
rect 24155 9160 24167 9163
rect 24198 9160 24204 9172
rect 24155 9132 24204 9160
rect 24155 9129 24167 9132
rect 24109 9123 24167 9129
rect 24198 9120 24204 9132
rect 24256 9160 24262 9172
rect 24256 9132 24520 9160
rect 24256 9120 24262 9132
rect 10674 9052 10680 9104
rect 10732 9092 10738 9104
rect 11226 9092 11232 9104
rect 10732 9064 11232 9092
rect 10732 9052 10738 9064
rect 11226 9052 11232 9064
rect 11284 9092 11290 9104
rect 11458 9095 11516 9101
rect 11458 9092 11470 9095
rect 11284 9064 11470 9092
rect 11284 9052 11290 9064
rect 11458 9061 11470 9064
rect 11504 9061 11516 9095
rect 13066 9092 13072 9104
rect 13027 9064 13072 9092
rect 11458 9055 11516 9061
rect 13066 9052 13072 9064
rect 13124 9052 13130 9104
rect 14998 9092 15004 9104
rect 14832 9064 15004 9092
rect 10214 9024 10220 9036
rect 10175 8996 10220 9024
rect 10214 8984 10220 8996
rect 10272 8984 10278 9036
rect 10309 9027 10367 9033
rect 10309 8993 10321 9027
rect 10355 9024 10367 9027
rect 10490 9024 10496 9036
rect 10355 8996 10496 9024
rect 10355 8993 10367 8996
rect 10309 8987 10367 8993
rect 10490 8984 10496 8996
rect 10548 9024 10554 9036
rect 10585 9027 10643 9033
rect 10585 9024 10597 9027
rect 10548 8996 10597 9024
rect 10548 8984 10554 8996
rect 10585 8993 10597 8996
rect 10631 8993 10643 9027
rect 10585 8987 10643 8993
rect 11042 8984 11048 9036
rect 11100 9024 11106 9036
rect 11137 9027 11195 9033
rect 11137 9024 11149 9027
rect 11100 8996 11149 9024
rect 11100 8984 11106 8996
rect 11137 8993 11149 8996
rect 11183 8993 11195 9027
rect 11137 8987 11195 8993
rect 13710 8984 13716 9036
rect 13768 9024 13774 9036
rect 14832 9033 14860 9064
rect 14998 9052 15004 9064
rect 15056 9092 15062 9104
rect 15550 9092 15556 9104
rect 15056 9064 15556 9092
rect 15056 9052 15062 9064
rect 15550 9052 15556 9064
rect 15608 9052 15614 9104
rect 16838 9092 16844 9104
rect 16799 9064 16844 9092
rect 16838 9052 16844 9064
rect 16896 9052 16902 9104
rect 17574 9052 17580 9104
rect 17632 9092 17638 9104
rect 17669 9095 17727 9101
rect 17669 9092 17681 9095
rect 17632 9064 17681 9092
rect 17632 9052 17638 9064
rect 17669 9061 17681 9064
rect 17715 9061 17727 9095
rect 17669 9055 17727 9061
rect 18862 9052 18868 9104
rect 18920 9092 18926 9104
rect 19785 9095 19843 9101
rect 19785 9092 19797 9095
rect 18920 9064 19797 9092
rect 18920 9052 18926 9064
rect 19785 9061 19797 9064
rect 19831 9061 19843 9095
rect 21438 9092 21444 9104
rect 21399 9064 21444 9092
rect 19785 9055 19843 9061
rect 21438 9052 21444 9064
rect 21496 9052 21502 9104
rect 21993 9095 22051 9101
rect 21993 9061 22005 9095
rect 22039 9092 22051 9095
rect 22729 9095 22787 9101
rect 22729 9092 22741 9095
rect 22039 9064 22741 9092
rect 22039 9061 22051 9064
rect 21993 9055 22051 9061
rect 22729 9061 22741 9064
rect 22775 9092 22787 9095
rect 22910 9092 22916 9104
rect 22775 9064 22916 9092
rect 22775 9061 22787 9064
rect 22729 9055 22787 9061
rect 22910 9052 22916 9064
rect 22968 9052 22974 9104
rect 23005 9095 23063 9101
rect 23005 9061 23017 9095
rect 23051 9092 23063 9095
rect 23370 9092 23376 9104
rect 23051 9064 23376 9092
rect 23051 9061 23063 9064
rect 23005 9055 23063 9061
rect 23370 9052 23376 9064
rect 23428 9052 23434 9104
rect 24290 9052 24296 9104
rect 24348 9092 24354 9104
rect 24385 9095 24443 9101
rect 24385 9092 24397 9095
rect 24348 9064 24397 9092
rect 24348 9052 24354 9064
rect 24385 9061 24397 9064
rect 24431 9061 24443 9095
rect 24385 9055 24443 9061
rect 14817 9027 14875 9033
rect 14817 9024 14829 9027
rect 13768 8996 14829 9024
rect 13768 8984 13774 8996
rect 14817 8993 14829 8996
rect 14863 8993 14875 9027
rect 14817 8987 14875 8993
rect 14906 8984 14912 9036
rect 14964 9024 14970 9036
rect 15645 9027 15703 9033
rect 15645 9024 15657 9027
rect 14964 8996 15657 9024
rect 14964 8984 14970 8996
rect 15645 8993 15657 8996
rect 15691 8993 15703 9027
rect 15645 8987 15703 8993
rect 19392 9027 19450 9033
rect 19392 8993 19404 9027
rect 19438 9024 19450 9027
rect 19690 9024 19696 9036
rect 19438 8996 19696 9024
rect 19438 8993 19450 8996
rect 19392 8987 19450 8993
rect 19690 8984 19696 8996
rect 19748 8984 19754 9036
rect 24492 9033 24520 9132
rect 24477 9027 24535 9033
rect 24477 8993 24489 9027
rect 24523 8993 24535 9027
rect 24477 8987 24535 8993
rect 11962 8916 11968 8968
rect 12020 8956 12026 8968
rect 12974 8956 12980 8968
rect 12020 8928 12980 8956
rect 12020 8916 12026 8928
rect 12974 8916 12980 8928
rect 13032 8916 13038 8968
rect 13342 8956 13348 8968
rect 13303 8928 13348 8956
rect 13342 8916 13348 8928
rect 13400 8916 13406 8968
rect 13802 8916 13808 8968
rect 13860 8956 13866 8968
rect 15553 8959 15611 8965
rect 15553 8956 15565 8959
rect 13860 8928 15565 8956
rect 13860 8916 13866 8928
rect 15553 8925 15565 8928
rect 15599 8925 15611 8959
rect 15553 8919 15611 8925
rect 16930 8916 16936 8968
rect 16988 8956 16994 8968
rect 17577 8959 17635 8965
rect 17577 8956 17589 8959
rect 16988 8928 17589 8956
rect 16988 8916 16994 8928
rect 17577 8925 17589 8928
rect 17623 8925 17635 8959
rect 17850 8956 17856 8968
rect 17811 8928 17856 8956
rect 17577 8919 17635 8925
rect 17850 8916 17856 8928
rect 17908 8916 17914 8968
rect 21349 8959 21407 8965
rect 21349 8925 21361 8959
rect 21395 8956 21407 8959
rect 21530 8956 21536 8968
rect 21395 8928 21536 8956
rect 21395 8925 21407 8928
rect 21349 8919 21407 8925
rect 21530 8916 21536 8928
rect 21588 8916 21594 8968
rect 23186 8956 23192 8968
rect 23147 8928 23192 8956
rect 23186 8916 23192 8928
rect 23244 8916 23250 8968
rect 15642 8888 15648 8900
rect 15603 8860 15648 8888
rect 15642 8848 15648 8860
rect 15700 8848 15706 8900
rect 17393 8891 17451 8897
rect 17393 8857 17405 8891
rect 17439 8888 17451 8891
rect 17666 8888 17672 8900
rect 17439 8860 17672 8888
rect 17439 8857 17451 8860
rect 17393 8851 17451 8857
rect 17666 8848 17672 8860
rect 17724 8848 17730 8900
rect 13894 8820 13900 8832
rect 13855 8792 13900 8820
rect 13894 8780 13900 8792
rect 13952 8780 13958 8832
rect 20886 8820 20892 8832
rect 20847 8792 20892 8820
rect 20886 8780 20892 8792
rect 20944 8780 20950 8832
rect 23462 8780 23468 8832
rect 23520 8820 23526 8832
rect 25118 8820 25124 8832
rect 23520 8792 25124 8820
rect 23520 8780 23526 8792
rect 25118 8780 25124 8792
rect 25176 8780 25182 8832
rect 632 8730 26392 8752
rect 632 8678 5176 8730
rect 5228 8678 5240 8730
rect 5292 8678 5304 8730
rect 5356 8678 5368 8730
rect 5420 8678 14510 8730
rect 14562 8678 14574 8730
rect 14626 8678 14638 8730
rect 14690 8678 14702 8730
rect 14754 8678 23843 8730
rect 23895 8678 23907 8730
rect 23959 8678 23971 8730
rect 24023 8678 24035 8730
rect 24087 8678 26392 8730
rect 632 8656 26392 8678
rect 9481 8619 9539 8625
rect 9481 8585 9493 8619
rect 9527 8616 9539 8619
rect 10214 8616 10220 8628
rect 9527 8588 10220 8616
rect 9527 8585 9539 8588
rect 9481 8579 9539 8585
rect 10214 8576 10220 8588
rect 10272 8576 10278 8628
rect 11226 8616 11232 8628
rect 11187 8588 11232 8616
rect 11226 8576 11232 8588
rect 11284 8576 11290 8628
rect 13434 8616 13440 8628
rect 13395 8588 13440 8616
rect 13434 8576 13440 8588
rect 13492 8576 13498 8628
rect 14998 8616 15004 8628
rect 14959 8588 15004 8616
rect 14998 8576 15004 8588
rect 15056 8576 15062 8628
rect 15734 8576 15740 8628
rect 15792 8616 15798 8628
rect 16930 8616 16936 8628
rect 15792 8588 16936 8616
rect 15792 8576 15798 8588
rect 16930 8576 16936 8588
rect 16988 8576 16994 8628
rect 19233 8619 19291 8625
rect 19233 8585 19245 8619
rect 19279 8616 19291 8619
rect 19966 8616 19972 8628
rect 19279 8588 19972 8616
rect 19279 8585 19291 8588
rect 19233 8579 19291 8585
rect 9386 8508 9392 8560
rect 9444 8548 9450 8560
rect 9757 8551 9815 8557
rect 9757 8548 9769 8551
rect 9444 8520 9769 8548
rect 9444 8508 9450 8520
rect 9757 8517 9769 8520
rect 9803 8517 9815 8551
rect 9757 8511 9815 8517
rect 11781 8551 11839 8557
rect 11781 8517 11793 8551
rect 11827 8548 11839 8551
rect 12054 8548 12060 8560
rect 11827 8520 12060 8548
rect 11827 8517 11839 8520
rect 11781 8511 11839 8517
rect 9772 8412 9800 8511
rect 12054 8508 12060 8520
rect 12112 8508 12118 8560
rect 14262 8548 14268 8560
rect 14223 8520 14268 8548
rect 14262 8508 14268 8520
rect 14320 8508 14326 8560
rect 10490 8480 10496 8492
rect 10451 8452 10496 8480
rect 10490 8440 10496 8452
rect 10548 8440 10554 8492
rect 9941 8415 9999 8421
rect 9941 8412 9953 8415
rect 9772 8384 9953 8412
rect 9941 8381 9953 8384
rect 9987 8381 9999 8415
rect 10398 8412 10404 8424
rect 10359 8384 10404 8412
rect 9941 8375 9999 8381
rect 10398 8372 10404 8384
rect 10456 8372 10462 8424
rect 12072 8421 12100 8508
rect 12701 8483 12759 8489
rect 12701 8449 12713 8483
rect 12747 8480 12759 8483
rect 12977 8483 13035 8489
rect 12977 8480 12989 8483
rect 12747 8452 12989 8480
rect 12747 8449 12759 8452
rect 12701 8443 12759 8449
rect 12977 8449 12989 8452
rect 13023 8480 13035 8483
rect 13066 8480 13072 8492
rect 13023 8452 13072 8480
rect 13023 8449 13035 8452
rect 12977 8443 13035 8449
rect 13066 8440 13072 8452
rect 13124 8440 13130 8492
rect 15461 8483 15519 8489
rect 15461 8449 15473 8483
rect 15507 8480 15519 8483
rect 15642 8480 15648 8492
rect 15507 8452 15648 8480
rect 15507 8449 15519 8452
rect 15461 8443 15519 8449
rect 15642 8440 15648 8452
rect 15700 8480 15706 8492
rect 16102 8480 16108 8492
rect 15700 8452 16108 8480
rect 15700 8440 15706 8452
rect 16102 8440 16108 8452
rect 16160 8440 16166 8492
rect 17393 8483 17451 8489
rect 17393 8449 17405 8483
rect 17439 8480 17451 8483
rect 17574 8480 17580 8492
rect 17439 8452 17580 8480
rect 17439 8449 17451 8452
rect 17393 8443 17451 8449
rect 17574 8440 17580 8452
rect 17632 8440 17638 8492
rect 12057 8415 12115 8421
rect 12057 8381 12069 8415
rect 12103 8381 12115 8415
rect 12057 8375 12115 8381
rect 13434 8372 13440 8424
rect 13492 8412 13498 8424
rect 13529 8415 13587 8421
rect 13529 8412 13541 8415
rect 13492 8384 13541 8412
rect 13492 8372 13498 8384
rect 13529 8381 13541 8384
rect 13575 8381 13587 8415
rect 13529 8375 13587 8381
rect 13802 8372 13808 8424
rect 13860 8412 13866 8424
rect 13989 8415 14047 8421
rect 13989 8412 14001 8415
rect 13860 8384 14001 8412
rect 13860 8372 13866 8384
rect 13989 8381 14001 8384
rect 14035 8381 14047 8415
rect 13989 8375 14047 8381
rect 14357 8415 14415 8421
rect 14357 8381 14369 8415
rect 14403 8381 14415 8415
rect 16378 8412 16384 8424
rect 16339 8384 16384 8412
rect 14357 8375 14415 8381
rect 8926 8344 8932 8356
rect 8887 8316 8932 8344
rect 8926 8304 8932 8316
rect 8984 8304 8990 8356
rect 13894 8304 13900 8356
rect 13952 8344 13958 8356
rect 14372 8344 14400 8375
rect 16378 8372 16384 8384
rect 16436 8372 16442 8424
rect 18221 8415 18279 8421
rect 18221 8381 18233 8415
rect 18267 8412 18279 8415
rect 18402 8412 18408 8424
rect 18267 8384 18408 8412
rect 18267 8381 18279 8384
rect 18221 8375 18279 8381
rect 18402 8372 18408 8384
rect 18460 8372 18466 8424
rect 18954 8372 18960 8424
rect 19012 8412 19018 8424
rect 19340 8421 19368 8588
rect 19966 8576 19972 8588
rect 20024 8616 20030 8628
rect 20150 8616 20156 8628
rect 20024 8588 20156 8616
rect 20024 8576 20030 8588
rect 20150 8576 20156 8588
rect 20208 8576 20214 8628
rect 20610 8576 20616 8628
rect 20668 8616 20674 8628
rect 20705 8619 20763 8625
rect 20705 8616 20717 8619
rect 20668 8588 20717 8616
rect 20668 8576 20674 8588
rect 20705 8585 20717 8588
rect 20751 8585 20763 8619
rect 20705 8579 20763 8585
rect 19325 8415 19383 8421
rect 19325 8412 19337 8415
rect 19012 8384 19337 8412
rect 19012 8372 19018 8384
rect 19325 8381 19337 8384
rect 19371 8381 19383 8415
rect 19782 8412 19788 8424
rect 19743 8384 19788 8412
rect 19325 8375 19383 8381
rect 19782 8372 19788 8384
rect 19840 8372 19846 8424
rect 20242 8372 20248 8424
rect 20300 8412 20306 8424
rect 20720 8412 20748 8579
rect 21438 8576 21444 8628
rect 21496 8616 21502 8628
rect 21898 8616 21904 8628
rect 21496 8588 21904 8616
rect 21496 8576 21502 8588
rect 21898 8576 21904 8588
rect 21956 8576 21962 8628
rect 22634 8616 22640 8628
rect 22595 8588 22640 8616
rect 22634 8576 22640 8588
rect 22692 8576 22698 8628
rect 23002 8616 23008 8628
rect 22963 8588 23008 8616
rect 23002 8576 23008 8588
rect 23060 8616 23066 8628
rect 23370 8616 23376 8628
rect 23060 8588 23376 8616
rect 23060 8576 23066 8588
rect 23370 8576 23376 8588
rect 23428 8576 23434 8628
rect 24198 8576 24204 8628
rect 24256 8616 24262 8628
rect 24385 8619 24443 8625
rect 24385 8616 24397 8619
rect 24256 8588 24397 8616
rect 24256 8576 24262 8588
rect 24385 8585 24397 8588
rect 24431 8585 24443 8619
rect 24934 8616 24940 8628
rect 24895 8588 24940 8616
rect 24385 8579 24443 8585
rect 24934 8576 24940 8588
rect 24992 8576 24998 8628
rect 23186 8508 23192 8560
rect 23244 8548 23250 8560
rect 23244 8520 23600 8548
rect 23244 8508 23250 8520
rect 23572 8489 23600 8520
rect 23557 8483 23615 8489
rect 23557 8449 23569 8483
rect 23603 8449 23615 8483
rect 23557 8443 23615 8449
rect 24198 8440 24204 8492
rect 24256 8480 24262 8492
rect 24474 8480 24480 8492
rect 24256 8452 24480 8480
rect 24256 8440 24262 8452
rect 24474 8440 24480 8452
rect 24532 8440 24538 8492
rect 20889 8415 20947 8421
rect 20889 8412 20901 8415
rect 20300 8384 20901 8412
rect 20300 8372 20306 8384
rect 20889 8381 20901 8384
rect 20935 8381 20947 8415
rect 20889 8375 20947 8381
rect 20978 8372 20984 8424
rect 21036 8412 21042 8424
rect 21349 8415 21407 8421
rect 21349 8412 21361 8415
rect 21036 8384 21361 8412
rect 21036 8372 21042 8384
rect 21349 8381 21361 8384
rect 21395 8381 21407 8415
rect 24750 8412 24756 8424
rect 24711 8384 24756 8412
rect 21349 8375 21407 8381
rect 24750 8372 24756 8384
rect 24808 8412 24814 8424
rect 25305 8415 25363 8421
rect 25305 8412 25317 8415
rect 24808 8384 25317 8412
rect 24808 8372 24814 8384
rect 25305 8381 25317 8384
rect 25351 8381 25363 8415
rect 25305 8375 25363 8381
rect 15366 8344 15372 8356
rect 13952 8316 14400 8344
rect 15279 8316 15372 8344
rect 13952 8304 13958 8316
rect 15366 8304 15372 8316
rect 15424 8344 15430 8356
rect 15823 8347 15881 8353
rect 15823 8344 15835 8347
rect 15424 8316 15835 8344
rect 15424 8304 15430 8316
rect 15823 8313 15835 8316
rect 15869 8344 15881 8347
rect 16746 8344 16752 8356
rect 15869 8316 16752 8344
rect 15869 8313 15881 8316
rect 15823 8307 15881 8313
rect 16746 8304 16752 8316
rect 16804 8304 16810 8356
rect 18865 8347 18923 8353
rect 18865 8313 18877 8347
rect 18911 8344 18923 8347
rect 19800 8344 19828 8372
rect 20058 8344 20064 8356
rect 18911 8316 19828 8344
rect 20019 8316 20064 8344
rect 18911 8313 18923 8316
rect 18865 8307 18923 8313
rect 20058 8304 20064 8316
rect 20116 8304 20122 8356
rect 23278 8344 23284 8356
rect 23239 8316 23284 8344
rect 23278 8304 23284 8316
rect 23336 8304 23342 8356
rect 23370 8304 23376 8356
rect 23428 8344 23434 8356
rect 23428 8316 23473 8344
rect 23428 8304 23434 8316
rect 21162 8276 21168 8288
rect 21123 8248 21168 8276
rect 21162 8236 21168 8248
rect 21220 8236 21226 8288
rect 632 8186 26392 8208
rect 632 8134 9843 8186
rect 9895 8134 9907 8186
rect 9959 8134 9971 8186
rect 10023 8134 10035 8186
rect 10087 8134 19176 8186
rect 19228 8134 19240 8186
rect 19292 8134 19304 8186
rect 19356 8134 19368 8186
rect 19420 8134 26392 8186
rect 632 8112 26392 8134
rect 10033 8075 10091 8081
rect 10033 8041 10045 8075
rect 10079 8072 10091 8075
rect 10398 8072 10404 8084
rect 10079 8044 10404 8072
rect 10079 8041 10091 8044
rect 10033 8035 10091 8041
rect 10398 8032 10404 8044
rect 10456 8032 10462 8084
rect 10582 8072 10588 8084
rect 10543 8044 10588 8072
rect 10582 8032 10588 8044
rect 10640 8032 10646 8084
rect 11042 8032 11048 8084
rect 11100 8072 11106 8084
rect 11321 8075 11379 8081
rect 11321 8072 11333 8075
rect 11100 8044 11333 8072
rect 11100 8032 11106 8044
rect 11321 8041 11333 8044
rect 11367 8041 11379 8075
rect 11321 8035 11379 8041
rect 12057 8075 12115 8081
rect 12057 8041 12069 8075
rect 12103 8072 12115 8075
rect 12606 8072 12612 8084
rect 12103 8044 12612 8072
rect 12103 8041 12115 8044
rect 12057 8035 12115 8041
rect 12606 8032 12612 8044
rect 12664 8032 12670 8084
rect 12974 8072 12980 8084
rect 12935 8044 12980 8072
rect 12974 8032 12980 8044
rect 13032 8032 13038 8084
rect 13802 8032 13808 8084
rect 13860 8072 13866 8084
rect 14173 8075 14231 8081
rect 14173 8072 14185 8075
rect 13860 8044 14185 8072
rect 13860 8032 13866 8044
rect 14173 8041 14185 8044
rect 14219 8072 14231 8075
rect 14354 8072 14360 8084
rect 14219 8044 14360 8072
rect 14219 8041 14231 8044
rect 14173 8035 14231 8041
rect 14354 8032 14360 8044
rect 14412 8032 14418 8084
rect 14633 8075 14691 8081
rect 14633 8041 14645 8075
rect 14679 8072 14691 8075
rect 14906 8072 14912 8084
rect 14679 8044 14912 8072
rect 14679 8041 14691 8044
rect 14633 8035 14691 8041
rect 14906 8032 14912 8044
rect 14964 8032 14970 8084
rect 15737 8075 15795 8081
rect 15737 8041 15749 8075
rect 15783 8072 15795 8075
rect 15826 8072 15832 8084
rect 15783 8044 15832 8072
rect 15783 8041 15795 8044
rect 15737 8035 15795 8041
rect 15826 8032 15832 8044
rect 15884 8032 15890 8084
rect 16102 8032 16108 8084
rect 16160 8072 16166 8084
rect 16381 8075 16439 8081
rect 16381 8072 16393 8075
rect 16160 8044 16393 8072
rect 16160 8032 16166 8044
rect 16381 8041 16393 8044
rect 16427 8041 16439 8075
rect 17758 8072 17764 8084
rect 17719 8044 17764 8072
rect 16381 8035 16439 8041
rect 17758 8032 17764 8044
rect 17816 8032 17822 8084
rect 18402 8072 18408 8084
rect 18363 8044 18408 8072
rect 18402 8032 18408 8044
rect 18460 8032 18466 8084
rect 19690 8032 19696 8084
rect 19748 8072 19754 8084
rect 19785 8075 19843 8081
rect 19785 8072 19797 8075
rect 19748 8044 19797 8072
rect 19748 8032 19754 8044
rect 19785 8041 19797 8044
rect 19831 8041 19843 8075
rect 19785 8035 19843 8041
rect 21622 8032 21628 8084
rect 21680 8072 21686 8084
rect 23278 8072 23284 8084
rect 21680 8044 21725 8072
rect 23239 8044 23284 8072
rect 21680 8032 21686 8044
rect 23278 8032 23284 8044
rect 23336 8032 23342 8084
rect 15179 8007 15237 8013
rect 15179 7973 15191 8007
rect 15225 8004 15237 8007
rect 15366 8004 15372 8016
rect 15225 7976 15372 8004
rect 15225 7973 15237 7976
rect 15179 7967 15237 7973
rect 15366 7964 15372 7976
rect 15424 7964 15430 8016
rect 16930 7964 16936 8016
rect 16988 8004 16994 8016
rect 20794 8013 20800 8016
rect 17162 8007 17220 8013
rect 17162 8004 17174 8007
rect 16988 7976 17174 8004
rect 16988 7964 16994 7976
rect 17162 7973 17174 7976
rect 17208 7973 17220 8007
rect 20791 8004 20800 8013
rect 20755 7976 20800 8004
rect 17162 7967 17220 7973
rect 20791 7967 20800 7976
rect 20794 7964 20800 7967
rect 20852 7964 20858 8016
rect 22361 8007 22419 8013
rect 22361 7973 22373 8007
rect 22407 8004 22419 8007
rect 22450 8004 22456 8016
rect 22407 7976 22456 8004
rect 22407 7973 22419 7976
rect 22361 7967 22419 7973
rect 22450 7964 22456 7976
rect 22508 7964 22514 8016
rect 8190 7936 8196 7948
rect 8151 7908 8196 7936
rect 8190 7896 8196 7908
rect 8248 7896 8254 7948
rect 9386 7896 9392 7948
rect 9444 7936 9450 7948
rect 10309 7939 10367 7945
rect 10309 7936 10321 7939
rect 9444 7908 10321 7936
rect 9444 7896 9450 7908
rect 10309 7905 10321 7908
rect 10355 7936 10367 7939
rect 10766 7936 10772 7948
rect 10355 7908 10772 7936
rect 10355 7905 10367 7908
rect 10309 7899 10367 7905
rect 10766 7896 10772 7908
rect 10824 7896 10830 7948
rect 10861 7939 10919 7945
rect 10861 7905 10873 7939
rect 10907 7936 10919 7939
rect 11502 7936 11508 7948
rect 10907 7908 11508 7936
rect 10907 7905 10919 7908
rect 10861 7899 10919 7905
rect 11502 7896 11508 7908
rect 11560 7896 11566 7948
rect 12216 7939 12274 7945
rect 12216 7905 12228 7939
rect 12262 7936 12274 7939
rect 12514 7936 12520 7948
rect 12262 7908 12520 7936
rect 12262 7905 12274 7908
rect 12216 7899 12274 7905
rect 12514 7896 12520 7908
rect 12572 7896 12578 7948
rect 13250 7936 13256 7948
rect 13211 7908 13256 7936
rect 13250 7896 13256 7908
rect 13308 7936 13314 7948
rect 14630 7936 14636 7948
rect 13308 7908 14636 7936
rect 13308 7896 13314 7908
rect 14630 7896 14636 7908
rect 14688 7896 14694 7948
rect 14814 7936 14820 7948
rect 14775 7908 14820 7936
rect 14814 7896 14820 7908
rect 14872 7896 14878 7948
rect 16194 7896 16200 7948
rect 16252 7936 16258 7948
rect 16841 7939 16899 7945
rect 16841 7936 16853 7939
rect 16252 7908 16853 7936
rect 16252 7896 16258 7908
rect 16841 7905 16853 7908
rect 16887 7936 16899 7939
rect 17022 7936 17028 7948
rect 16887 7908 17028 7936
rect 16887 7905 16899 7908
rect 16841 7899 16899 7905
rect 17022 7896 17028 7908
rect 17080 7896 17086 7948
rect 18954 7936 18960 7948
rect 18915 7908 18960 7936
rect 18954 7896 18960 7908
rect 19012 7896 19018 7948
rect 19046 7896 19052 7948
rect 19104 7936 19110 7948
rect 19233 7939 19291 7945
rect 19233 7936 19245 7939
rect 19104 7908 19245 7936
rect 19104 7896 19110 7908
rect 19233 7905 19245 7908
rect 19279 7905 19291 7939
rect 19233 7899 19291 7905
rect 23186 7896 23192 7948
rect 23244 7936 23250 7948
rect 23833 7939 23891 7945
rect 23833 7936 23845 7939
rect 23244 7908 23845 7936
rect 23244 7896 23250 7908
rect 23833 7905 23845 7908
rect 23879 7905 23891 7939
rect 23833 7899 23891 7905
rect 8282 7868 8288 7880
rect 8243 7840 8288 7868
rect 8282 7828 8288 7840
rect 8340 7828 8346 7880
rect 9297 7871 9355 7877
rect 9297 7837 9309 7871
rect 9343 7868 9355 7871
rect 10398 7868 10404 7880
rect 9343 7840 10404 7868
rect 9343 7837 9355 7840
rect 9297 7831 9355 7837
rect 10398 7828 10404 7840
rect 10456 7828 10462 7880
rect 13894 7868 13900 7880
rect 13855 7840 13900 7868
rect 13894 7828 13900 7840
rect 13952 7828 13958 7880
rect 14354 7828 14360 7880
rect 14412 7868 14418 7880
rect 16013 7871 16071 7877
rect 16013 7868 16025 7871
rect 14412 7840 16025 7868
rect 14412 7828 14418 7840
rect 16013 7837 16025 7840
rect 16059 7837 16071 7871
rect 16013 7831 16071 7837
rect 19509 7871 19567 7877
rect 19509 7837 19521 7871
rect 19555 7868 19567 7871
rect 20429 7871 20487 7877
rect 20429 7868 20441 7871
rect 19555 7840 20441 7868
rect 19555 7837 19567 7840
rect 19509 7831 19567 7837
rect 20429 7837 20441 7840
rect 20475 7868 20487 7871
rect 20886 7868 20892 7880
rect 20475 7840 20892 7868
rect 20475 7837 20487 7840
rect 20429 7831 20487 7837
rect 20886 7828 20892 7840
rect 20944 7828 20950 7880
rect 22269 7871 22327 7877
rect 22269 7837 22281 7871
rect 22315 7868 22327 7871
rect 22358 7868 22364 7880
rect 22315 7840 22364 7868
rect 22315 7837 22327 7840
rect 22269 7831 22327 7837
rect 22358 7828 22364 7840
rect 22416 7828 22422 7880
rect 22542 7868 22548 7880
rect 22503 7840 22548 7868
rect 22542 7828 22548 7840
rect 22600 7868 22606 7880
rect 23557 7871 23615 7877
rect 23557 7868 23569 7871
rect 22600 7840 23569 7868
rect 22600 7828 22606 7840
rect 23557 7837 23569 7840
rect 23603 7837 23615 7871
rect 23738 7868 23744 7880
rect 23699 7840 23744 7868
rect 23557 7831 23615 7837
rect 23738 7828 23744 7840
rect 23796 7828 23802 7880
rect 12330 7809 12336 7812
rect 12287 7803 12336 7809
rect 12287 7769 12299 7803
rect 12333 7769 12336 7803
rect 12287 7763 12336 7769
rect 12330 7760 12336 7763
rect 12388 7760 12394 7812
rect 18126 7732 18132 7744
rect 18087 7704 18132 7732
rect 18126 7692 18132 7704
rect 18184 7692 18190 7744
rect 21346 7732 21352 7744
rect 21307 7704 21352 7732
rect 21346 7692 21352 7704
rect 21404 7692 21410 7744
rect 632 7642 26392 7664
rect 632 7590 5176 7642
rect 5228 7590 5240 7642
rect 5292 7590 5304 7642
rect 5356 7590 5368 7642
rect 5420 7590 14510 7642
rect 14562 7590 14574 7642
rect 14626 7590 14638 7642
rect 14690 7590 14702 7642
rect 14754 7590 23843 7642
rect 23895 7590 23907 7642
rect 23959 7590 23971 7642
rect 24023 7590 24035 7642
rect 24087 7590 26392 7642
rect 632 7568 26392 7590
rect 7641 7531 7699 7537
rect 7641 7497 7653 7531
rect 7687 7528 7699 7531
rect 8190 7528 8196 7540
rect 7687 7500 8196 7528
rect 7687 7497 7699 7500
rect 7641 7491 7699 7497
rect 8190 7488 8196 7500
rect 8248 7488 8254 7540
rect 10217 7531 10275 7537
rect 10217 7497 10229 7531
rect 10263 7528 10275 7531
rect 10306 7528 10312 7540
rect 10263 7500 10312 7528
rect 10263 7497 10275 7500
rect 10217 7491 10275 7497
rect 10306 7488 10312 7500
rect 10364 7488 10370 7540
rect 11413 7531 11471 7537
rect 11413 7497 11425 7531
rect 11459 7528 11471 7531
rect 11502 7528 11508 7540
rect 11459 7500 11508 7528
rect 11459 7497 11471 7500
rect 11413 7491 11471 7497
rect 7730 7392 7736 7404
rect 7691 7364 7736 7392
rect 7730 7352 7736 7364
rect 7788 7352 7794 7404
rect 8653 7395 8711 7401
rect 8653 7361 8665 7395
rect 8699 7392 8711 7395
rect 9386 7392 9392 7404
rect 8699 7364 9392 7392
rect 8699 7361 8711 7364
rect 8653 7355 8711 7361
rect 9036 7333 9064 7364
rect 9386 7352 9392 7364
rect 9444 7352 9450 7404
rect 9849 7395 9907 7401
rect 9849 7361 9861 7395
rect 9895 7392 9907 7395
rect 9895 7364 10904 7392
rect 9895 7361 9907 7364
rect 9849 7355 9907 7361
rect 9021 7327 9079 7333
rect 9021 7293 9033 7327
rect 9067 7293 9079 7327
rect 9294 7324 9300 7336
rect 9255 7296 9300 7324
rect 9021 7287 9079 7293
rect 9294 7284 9300 7296
rect 9352 7284 9358 7336
rect 10306 7324 10312 7336
rect 10267 7296 10312 7324
rect 10306 7284 10312 7296
rect 10364 7284 10370 7336
rect 10876 7333 10904 7364
rect 10861 7327 10919 7333
rect 10861 7293 10873 7327
rect 10907 7324 10919 7327
rect 11428 7324 11456 7491
rect 11502 7488 11508 7500
rect 11560 7488 11566 7540
rect 13069 7531 13127 7537
rect 13069 7497 13081 7531
rect 13115 7528 13127 7531
rect 13250 7528 13256 7540
rect 13115 7500 13256 7528
rect 13115 7497 13127 7500
rect 13069 7491 13127 7497
rect 13250 7488 13256 7500
rect 13308 7488 13314 7540
rect 13434 7488 13440 7540
rect 13492 7528 13498 7540
rect 13621 7531 13679 7537
rect 13621 7528 13633 7531
rect 13492 7500 13633 7528
rect 13492 7488 13498 7500
rect 13621 7497 13633 7500
rect 13667 7528 13679 7531
rect 13713 7531 13771 7537
rect 13713 7528 13725 7531
rect 13667 7500 13725 7528
rect 13667 7497 13679 7500
rect 13621 7491 13679 7497
rect 13713 7497 13725 7500
rect 13759 7497 13771 7531
rect 15366 7528 15372 7540
rect 15327 7500 15372 7528
rect 13713 7491 13771 7497
rect 15366 7488 15372 7500
rect 15424 7488 15430 7540
rect 15737 7531 15795 7537
rect 15737 7497 15749 7531
rect 15783 7528 15795 7531
rect 15826 7528 15832 7540
rect 15783 7500 15832 7528
rect 15783 7497 15795 7500
rect 15737 7491 15795 7497
rect 15826 7488 15832 7500
rect 15884 7488 15890 7540
rect 17022 7488 17028 7540
rect 17080 7528 17086 7540
rect 17209 7531 17267 7537
rect 17209 7528 17221 7531
rect 17080 7500 17221 7528
rect 17080 7488 17086 7500
rect 17209 7497 17221 7500
rect 17255 7497 17267 7531
rect 17209 7491 17267 7497
rect 18954 7488 18960 7540
rect 19012 7528 19018 7540
rect 19049 7531 19107 7537
rect 19049 7528 19061 7531
rect 19012 7500 19061 7528
rect 19012 7488 19018 7500
rect 19049 7497 19061 7500
rect 19095 7497 19107 7531
rect 19049 7491 19107 7497
rect 19509 7531 19567 7537
rect 19509 7497 19521 7531
rect 19555 7528 19567 7531
rect 20150 7528 20156 7540
rect 19555 7500 20156 7528
rect 19555 7497 19567 7500
rect 19509 7491 19567 7497
rect 14630 7460 14636 7472
rect 14591 7432 14636 7460
rect 14630 7420 14636 7432
rect 14688 7420 14694 7472
rect 13437 7395 13495 7401
rect 13437 7392 13449 7395
rect 12256 7364 13449 7392
rect 12256 7333 12284 7364
rect 13437 7361 13449 7364
rect 13483 7392 13495 7395
rect 17850 7392 17856 7404
rect 13483 7364 14768 7392
rect 17811 7364 17856 7392
rect 13483 7361 13495 7364
rect 13437 7355 13495 7361
rect 12241 7327 12299 7333
rect 12241 7324 12253 7327
rect 10907 7296 11456 7324
rect 11704 7296 12253 7324
rect 10907 7293 10919 7296
rect 10861 7287 10919 7293
rect 9481 7259 9539 7265
rect 9481 7225 9493 7259
rect 9527 7256 9539 7259
rect 10214 7256 10220 7268
rect 9527 7228 10220 7256
rect 9527 7225 9539 7228
rect 9481 7219 9539 7225
rect 10214 7216 10220 7228
rect 10272 7216 10278 7268
rect 10324 7188 10352 7284
rect 11042 7256 11048 7268
rect 11003 7228 11048 7256
rect 11042 7216 11048 7228
rect 11100 7216 11106 7268
rect 11704 7200 11732 7296
rect 12241 7293 12253 7296
rect 12287 7293 12299 7327
rect 12241 7287 12299 7293
rect 12517 7327 12575 7333
rect 12517 7293 12529 7327
rect 12563 7324 12575 7327
rect 12606 7324 12612 7336
rect 12563 7296 12612 7324
rect 12563 7293 12575 7296
rect 12517 7287 12575 7293
rect 12606 7284 12612 7296
rect 12664 7284 12670 7336
rect 13621 7327 13679 7333
rect 13621 7293 13633 7327
rect 13667 7324 13679 7327
rect 13897 7327 13955 7333
rect 13897 7324 13909 7327
rect 13667 7296 13909 7324
rect 13667 7293 13679 7296
rect 13621 7287 13679 7293
rect 13897 7293 13909 7296
rect 13943 7293 13955 7327
rect 14354 7324 14360 7336
rect 14315 7296 14360 7324
rect 13897 7287 13955 7293
rect 14354 7284 14360 7296
rect 14412 7284 14418 7336
rect 14740 7333 14768 7364
rect 17850 7352 17856 7364
rect 17908 7352 17914 7404
rect 18402 7392 18408 7404
rect 18363 7364 18408 7392
rect 18402 7352 18408 7364
rect 18460 7352 18466 7404
rect 19616 7336 19644 7500
rect 20150 7488 20156 7500
rect 20208 7488 20214 7540
rect 20705 7531 20763 7537
rect 20705 7497 20717 7531
rect 20751 7528 20763 7531
rect 20794 7528 20800 7540
rect 20751 7500 20800 7528
rect 20751 7497 20763 7500
rect 20705 7491 20763 7497
rect 20794 7488 20800 7500
rect 20852 7528 20858 7540
rect 20981 7531 21039 7537
rect 20981 7528 20993 7531
rect 20852 7500 20993 7528
rect 20852 7488 20858 7500
rect 20981 7497 20993 7500
rect 21027 7497 21039 7531
rect 20981 7491 21039 7497
rect 20150 7392 20156 7404
rect 20111 7364 20156 7392
rect 20150 7352 20156 7364
rect 20208 7352 20214 7404
rect 14725 7327 14783 7333
rect 14725 7293 14737 7327
rect 14771 7324 14783 7327
rect 14906 7324 14912 7336
rect 14771 7296 14912 7324
rect 14771 7293 14783 7296
rect 14725 7287 14783 7293
rect 14906 7284 14912 7296
rect 14964 7284 14970 7336
rect 15826 7284 15832 7336
rect 15884 7324 15890 7336
rect 15921 7327 15979 7333
rect 15921 7324 15933 7327
rect 15884 7296 15933 7324
rect 15884 7284 15890 7296
rect 15921 7293 15933 7296
rect 15967 7293 15979 7327
rect 19598 7324 19604 7336
rect 19511 7296 19604 7324
rect 15921 7287 15979 7293
rect 19598 7284 19604 7296
rect 19656 7284 19662 7336
rect 19782 7284 19788 7336
rect 19840 7324 19846 7336
rect 20061 7327 20119 7333
rect 20061 7324 20073 7327
rect 19840 7296 20073 7324
rect 19840 7284 19846 7296
rect 20061 7293 20073 7296
rect 20107 7293 20119 7327
rect 20061 7287 20119 7293
rect 20996 7268 21024 7491
rect 21346 7488 21352 7540
rect 21404 7528 21410 7540
rect 22450 7528 22456 7540
rect 21404 7500 22456 7528
rect 21404 7488 21410 7500
rect 22450 7488 22456 7500
rect 22508 7488 22514 7540
rect 21162 7392 21168 7404
rect 21123 7364 21168 7392
rect 21162 7352 21168 7364
rect 21220 7352 21226 7404
rect 22542 7352 22548 7404
rect 22600 7392 22606 7404
rect 23281 7395 23339 7401
rect 23281 7392 23293 7395
rect 22600 7364 23293 7392
rect 22600 7352 22606 7364
rect 23281 7361 23293 7364
rect 23327 7361 23339 7395
rect 23554 7392 23560 7404
rect 23515 7364 23560 7392
rect 23281 7355 23339 7361
rect 23554 7352 23560 7364
rect 23612 7352 23618 7404
rect 22085 7327 22143 7333
rect 22085 7293 22097 7327
rect 22131 7324 22143 7327
rect 24750 7324 24756 7336
rect 22131 7296 23048 7324
rect 24711 7296 24756 7324
rect 22131 7293 22143 7296
rect 22085 7287 22143 7293
rect 16930 7256 16936 7268
rect 16891 7228 16936 7256
rect 16930 7216 16936 7228
rect 16988 7216 16994 7268
rect 18126 7256 18132 7268
rect 18087 7228 18132 7256
rect 18126 7216 18132 7228
rect 18184 7216 18190 7268
rect 18221 7259 18279 7265
rect 18221 7225 18233 7259
rect 18267 7225 18279 7259
rect 20978 7256 20984 7268
rect 20891 7228 20984 7256
rect 18221 7219 18279 7225
rect 11686 7188 11692 7200
rect 10324 7160 11692 7188
rect 11686 7148 11692 7160
rect 11744 7148 11750 7200
rect 11962 7148 11968 7200
rect 12020 7188 12026 7200
rect 12057 7191 12115 7197
rect 12057 7188 12069 7191
rect 12020 7160 12069 7188
rect 12020 7148 12026 7160
rect 12057 7157 12069 7160
rect 12103 7157 12115 7191
rect 16102 7188 16108 7200
rect 16063 7160 16108 7188
rect 12057 7151 12115 7157
rect 16102 7148 16108 7160
rect 16160 7148 16166 7200
rect 17850 7148 17856 7200
rect 17908 7188 17914 7200
rect 18236 7188 18264 7219
rect 20978 7216 20984 7228
rect 21036 7256 21042 7268
rect 23020 7265 23048 7296
rect 24750 7284 24756 7296
rect 24808 7324 24814 7336
rect 25305 7327 25363 7333
rect 25305 7324 25317 7327
rect 24808 7296 25317 7324
rect 24808 7284 24814 7296
rect 25305 7293 25317 7296
rect 25351 7293 25363 7327
rect 25305 7287 25363 7293
rect 21486 7259 21544 7265
rect 21486 7256 21498 7259
rect 21036 7228 21498 7256
rect 21036 7216 21042 7228
rect 21486 7225 21498 7228
rect 21532 7225 21544 7259
rect 21486 7219 21544 7225
rect 23005 7259 23063 7265
rect 23005 7225 23017 7259
rect 23051 7256 23063 7259
rect 23373 7259 23431 7265
rect 23373 7256 23385 7259
rect 23051 7228 23385 7256
rect 23051 7225 23063 7228
rect 23005 7219 23063 7225
rect 23373 7225 23385 7228
rect 23419 7256 23431 7259
rect 24658 7256 24664 7268
rect 23419 7228 24664 7256
rect 23419 7225 23431 7228
rect 23373 7219 23431 7225
rect 24658 7216 24664 7228
rect 24716 7216 24722 7268
rect 17908 7160 18264 7188
rect 17908 7148 17914 7160
rect 23186 7148 23192 7200
rect 23244 7188 23250 7200
rect 23738 7188 23744 7200
rect 23244 7160 23744 7188
rect 23244 7148 23250 7160
rect 23738 7148 23744 7160
rect 23796 7188 23802 7200
rect 24201 7191 24259 7197
rect 24201 7188 24213 7191
rect 23796 7160 24213 7188
rect 23796 7148 23802 7160
rect 24201 7157 24213 7160
rect 24247 7157 24259 7191
rect 24934 7188 24940 7200
rect 24895 7160 24940 7188
rect 24201 7151 24259 7157
rect 24934 7148 24940 7160
rect 24992 7148 24998 7200
rect 632 7098 26392 7120
rect 632 7046 9843 7098
rect 9895 7046 9907 7098
rect 9959 7046 9971 7098
rect 10023 7046 10035 7098
rect 10087 7046 19176 7098
rect 19228 7046 19240 7098
rect 19292 7046 19304 7098
rect 19356 7046 19368 7098
rect 19420 7046 26392 7098
rect 632 7024 26392 7046
rect 12514 6944 12520 6996
rect 12572 6984 12578 6996
rect 12609 6987 12667 6993
rect 12609 6984 12621 6987
rect 12572 6956 12621 6984
rect 12572 6944 12578 6956
rect 12609 6953 12621 6956
rect 12655 6953 12667 6987
rect 12609 6947 12667 6953
rect 14265 6987 14323 6993
rect 14265 6953 14277 6987
rect 14311 6984 14323 6987
rect 14354 6984 14360 6996
rect 14311 6956 14360 6984
rect 14311 6953 14323 6956
rect 14265 6947 14323 6953
rect 14354 6944 14360 6956
rect 14412 6944 14418 6996
rect 14814 6944 14820 6996
rect 14872 6984 14878 6996
rect 15277 6987 15335 6993
rect 15277 6984 15289 6987
rect 14872 6956 15289 6984
rect 14872 6944 14878 6956
rect 15277 6953 15289 6956
rect 15323 6953 15335 6987
rect 19046 6984 19052 6996
rect 19007 6956 19052 6984
rect 15277 6947 15335 6953
rect 19046 6944 19052 6956
rect 19104 6944 19110 6996
rect 19693 6987 19751 6993
rect 19693 6953 19705 6987
rect 19739 6984 19751 6987
rect 19782 6984 19788 6996
rect 19739 6956 19788 6984
rect 19739 6953 19751 6956
rect 19693 6947 19751 6953
rect 19782 6944 19788 6956
rect 19840 6944 19846 6996
rect 20886 6984 20892 6996
rect 20847 6956 20892 6984
rect 20886 6944 20892 6956
rect 20944 6944 20950 6996
rect 21162 6944 21168 6996
rect 21220 6984 21226 6996
rect 21257 6987 21315 6993
rect 21257 6984 21269 6987
rect 21220 6956 21269 6984
rect 21220 6944 21226 6956
rect 21257 6953 21269 6956
rect 21303 6953 21315 6987
rect 21257 6947 21315 6953
rect 22358 6944 22364 6996
rect 22416 6984 22422 6996
rect 22453 6987 22511 6993
rect 22453 6984 22465 6987
rect 22416 6956 22465 6984
rect 22416 6944 22422 6956
rect 22453 6953 22465 6956
rect 22499 6953 22511 6987
rect 22453 6947 22511 6953
rect 9294 6916 9300 6928
rect 9128 6888 9300 6916
rect 8098 6848 8104 6860
rect 8059 6820 8104 6848
rect 8098 6808 8104 6820
rect 8156 6808 8162 6860
rect 8837 6851 8895 6857
rect 8837 6817 8849 6851
rect 8883 6848 8895 6851
rect 9128 6848 9156 6888
rect 9294 6876 9300 6888
rect 9352 6876 9358 6928
rect 10211 6919 10269 6925
rect 10211 6885 10223 6919
rect 10257 6916 10269 6919
rect 13342 6916 13348 6928
rect 10257 6888 10628 6916
rect 13303 6888 13348 6916
rect 10257 6885 10269 6888
rect 10211 6879 10269 6885
rect 8883 6820 9156 6848
rect 9849 6851 9907 6857
rect 8883 6817 8895 6820
rect 8837 6811 8895 6817
rect 9849 6817 9861 6851
rect 9895 6848 9907 6851
rect 10490 6848 10496 6860
rect 9895 6820 10496 6848
rect 9895 6817 9907 6820
rect 9849 6811 9907 6817
rect 10490 6808 10496 6820
rect 10548 6808 10554 6860
rect 10600 6848 10628 6888
rect 13342 6876 13348 6888
rect 13400 6876 13406 6928
rect 17758 6876 17764 6928
rect 17816 6916 17822 6928
rect 18129 6919 18187 6925
rect 18129 6916 18141 6919
rect 17816 6888 18141 6916
rect 17816 6876 17822 6888
rect 18129 6885 18141 6888
rect 18175 6885 18187 6919
rect 18129 6879 18187 6885
rect 21622 6876 21628 6928
rect 21680 6916 21686 6928
rect 22177 6919 22235 6925
rect 21680 6888 21725 6916
rect 21680 6876 21686 6888
rect 22177 6885 22189 6919
rect 22223 6916 22235 6919
rect 22542 6916 22548 6928
rect 22223 6888 22548 6916
rect 22223 6885 22235 6888
rect 22177 6879 22235 6885
rect 22542 6876 22548 6888
rect 22600 6876 22606 6928
rect 23373 6919 23431 6925
rect 23373 6885 23385 6919
rect 23419 6916 23431 6919
rect 23646 6916 23652 6928
rect 23419 6888 23652 6916
rect 23419 6885 23431 6888
rect 23373 6879 23431 6885
rect 23646 6876 23652 6888
rect 23704 6876 23710 6928
rect 10674 6848 10680 6860
rect 10600 6820 10680 6848
rect 10674 6808 10680 6820
rect 10732 6808 10738 6860
rect 10766 6808 10772 6860
rect 10824 6848 10830 6860
rect 11045 6851 11103 6857
rect 11045 6848 11057 6851
rect 10824 6820 11057 6848
rect 10824 6808 10830 6820
rect 11045 6817 11057 6820
rect 11091 6817 11103 6851
rect 11686 6848 11692 6860
rect 11647 6820 11692 6848
rect 11045 6811 11103 6817
rect 11686 6808 11692 6820
rect 11744 6808 11750 6860
rect 12146 6848 12152 6860
rect 12107 6820 12152 6848
rect 12146 6808 12152 6820
rect 12204 6808 12210 6860
rect 14884 6851 14942 6857
rect 14884 6817 14896 6851
rect 14930 6848 14942 6851
rect 15734 6848 15740 6860
rect 14930 6820 15740 6848
rect 14930 6817 14942 6820
rect 14884 6811 14942 6817
rect 15734 6808 15740 6820
rect 15792 6808 15798 6860
rect 16378 6848 16384 6860
rect 16339 6820 16384 6848
rect 16378 6808 16384 6820
rect 16436 6808 16442 6860
rect 20426 6808 20432 6860
rect 20484 6857 20490 6860
rect 20610 6857 20616 6860
rect 20484 6851 20522 6857
rect 20510 6817 20522 6851
rect 20484 6811 20522 6817
rect 20567 6851 20616 6857
rect 20567 6817 20579 6851
rect 20613 6817 20616 6851
rect 20567 6811 20616 6817
rect 20484 6808 20490 6811
rect 20610 6808 20616 6811
rect 20668 6808 20674 6860
rect 24566 6808 24572 6860
rect 24624 6848 24630 6860
rect 24753 6851 24811 6857
rect 24753 6848 24765 6851
rect 24624 6820 24765 6848
rect 24624 6808 24630 6820
rect 24753 6817 24765 6820
rect 24799 6817 24811 6851
rect 24753 6811 24811 6817
rect 12330 6780 12336 6792
rect 12291 6752 12336 6780
rect 12330 6740 12336 6752
rect 12388 6740 12394 6792
rect 13250 6780 13256 6792
rect 13211 6752 13256 6780
rect 13250 6740 13256 6752
rect 13308 6740 13314 6792
rect 13897 6783 13955 6789
rect 13897 6749 13909 6783
rect 13943 6780 13955 6783
rect 16010 6780 16016 6792
rect 13943 6752 16016 6780
rect 13943 6749 13955 6752
rect 13897 6743 13955 6749
rect 16010 6740 16016 6752
rect 16068 6740 16074 6792
rect 16565 6783 16623 6789
rect 16565 6749 16577 6783
rect 16611 6780 16623 6783
rect 16746 6780 16752 6792
rect 16611 6752 16752 6780
rect 16611 6749 16623 6752
rect 16565 6743 16623 6749
rect 16746 6740 16752 6752
rect 16804 6740 16810 6792
rect 18034 6780 18040 6792
rect 17995 6752 18040 6780
rect 18034 6740 18040 6752
rect 18092 6740 18098 6792
rect 18402 6780 18408 6792
rect 18363 6752 18408 6780
rect 18402 6740 18408 6752
rect 18460 6740 18466 6792
rect 21346 6740 21352 6792
rect 21404 6780 21410 6792
rect 21533 6783 21591 6789
rect 21533 6780 21545 6783
rect 21404 6752 21545 6780
rect 21404 6740 21410 6752
rect 21533 6749 21545 6752
rect 21579 6749 21591 6783
rect 21533 6743 21591 6749
rect 23094 6740 23100 6792
rect 23152 6780 23158 6792
rect 23281 6783 23339 6789
rect 23281 6780 23293 6783
rect 23152 6752 23293 6780
rect 23152 6740 23158 6752
rect 23281 6749 23293 6752
rect 23327 6749 23339 6783
rect 23554 6780 23560 6792
rect 23515 6752 23560 6780
rect 23281 6743 23339 6749
rect 23554 6740 23560 6752
rect 23612 6740 23618 6792
rect 10766 6644 10772 6656
rect 10727 6616 10772 6644
rect 10766 6604 10772 6616
rect 10824 6604 10830 6656
rect 14955 6647 15013 6653
rect 14955 6613 14967 6647
rect 15001 6644 15013 6647
rect 15090 6644 15096 6656
rect 15001 6616 15096 6644
rect 15001 6613 15013 6616
rect 14955 6607 15013 6613
rect 15090 6604 15096 6616
rect 15148 6604 15154 6656
rect 15734 6644 15740 6656
rect 15695 6616 15740 6644
rect 15734 6604 15740 6616
rect 15792 6604 15798 6656
rect 24937 6647 24995 6653
rect 24937 6613 24949 6647
rect 24983 6644 24995 6647
rect 25854 6644 25860 6656
rect 24983 6616 25860 6644
rect 24983 6613 24995 6616
rect 24937 6607 24995 6613
rect 25854 6604 25860 6616
rect 25912 6604 25918 6656
rect 632 6554 26392 6576
rect 632 6502 5176 6554
rect 5228 6502 5240 6554
rect 5292 6502 5304 6554
rect 5356 6502 5368 6554
rect 5420 6502 14510 6554
rect 14562 6502 14574 6554
rect 14626 6502 14638 6554
rect 14690 6502 14702 6554
rect 14754 6502 23843 6554
rect 23895 6502 23907 6554
rect 23959 6502 23971 6554
rect 24023 6502 24035 6554
rect 24087 6502 26392 6554
rect 632 6480 26392 6502
rect 6534 6449 6540 6452
rect 6491 6443 6540 6449
rect 6491 6409 6503 6443
rect 6537 6409 6540 6443
rect 6491 6403 6540 6409
rect 6534 6400 6540 6403
rect 6592 6400 6598 6452
rect 9665 6443 9723 6449
rect 9665 6409 9677 6443
rect 9711 6440 9723 6443
rect 10033 6443 10091 6449
rect 10033 6440 10045 6443
rect 9711 6412 10045 6440
rect 9711 6409 9723 6412
rect 9665 6403 9723 6409
rect 10033 6409 10045 6412
rect 10079 6440 10091 6443
rect 10398 6440 10404 6452
rect 10079 6412 10404 6440
rect 10079 6409 10091 6412
rect 10033 6403 10091 6409
rect 10398 6400 10404 6412
rect 10456 6440 10462 6452
rect 10674 6440 10680 6452
rect 10456 6412 10680 6440
rect 10456 6400 10462 6412
rect 10674 6400 10680 6412
rect 10732 6440 10738 6452
rect 11410 6440 11416 6452
rect 10732 6412 11416 6440
rect 10732 6400 10738 6412
rect 11410 6400 11416 6412
rect 11468 6440 11474 6452
rect 11689 6443 11747 6449
rect 11689 6440 11701 6443
rect 11468 6412 11701 6440
rect 11468 6400 11474 6412
rect 11689 6409 11701 6412
rect 11735 6409 11747 6443
rect 11689 6403 11747 6409
rect 8098 6304 8104 6316
rect 8059 6276 8104 6304
rect 8098 6264 8104 6276
rect 8156 6264 8162 6316
rect 6166 6196 6172 6248
rect 6224 6236 6230 6248
rect 6399 6239 6457 6245
rect 6399 6236 6411 6239
rect 6224 6208 6411 6236
rect 6224 6196 6230 6208
rect 6399 6205 6411 6208
rect 6445 6236 6457 6239
rect 6813 6239 6871 6245
rect 6813 6236 6825 6239
rect 6445 6208 6825 6236
rect 6445 6205 6457 6208
rect 6399 6199 6457 6205
rect 6813 6205 6825 6208
rect 6859 6205 6871 6239
rect 6813 6199 6871 6205
rect 7600 6239 7658 6245
rect 7600 6205 7612 6239
rect 7646 6236 7658 6239
rect 8116 6236 8144 6264
rect 7646 6208 8144 6236
rect 8469 6239 8527 6245
rect 7646 6205 7658 6208
rect 7600 6199 7658 6205
rect 8469 6205 8481 6239
rect 8515 6236 8527 6239
rect 9202 6236 9208 6248
rect 8515 6208 9208 6236
rect 8515 6205 8527 6208
rect 8469 6199 8527 6205
rect 9202 6196 9208 6208
rect 9260 6196 9266 6248
rect 10125 6239 10183 6245
rect 10125 6205 10137 6239
rect 10171 6236 10183 6239
rect 10858 6236 10864 6248
rect 10171 6208 10864 6236
rect 10171 6205 10183 6208
rect 10125 6199 10183 6205
rect 10858 6196 10864 6208
rect 10916 6196 10922 6248
rect 7730 6177 7736 6180
rect 7687 6171 7736 6177
rect 7687 6137 7699 6171
rect 7733 6137 7736 6171
rect 7687 6131 7736 6137
rect 7730 6128 7736 6131
rect 7788 6128 7794 6180
rect 10398 6128 10404 6180
rect 10456 6177 10462 6180
rect 10456 6171 10504 6177
rect 10456 6137 10458 6171
rect 10492 6137 10504 6171
rect 11704 6168 11732 6403
rect 13250 6400 13256 6452
rect 13308 6440 13314 6452
rect 13529 6443 13587 6449
rect 13529 6440 13541 6443
rect 13308 6412 13541 6440
rect 13308 6400 13314 6412
rect 13529 6409 13541 6412
rect 13575 6409 13587 6443
rect 13529 6403 13587 6409
rect 17758 6400 17764 6452
rect 17816 6440 17822 6452
rect 18589 6443 18647 6449
rect 18589 6440 18601 6443
rect 17816 6412 18601 6440
rect 17816 6400 17822 6412
rect 18589 6409 18601 6412
rect 18635 6409 18647 6443
rect 19598 6440 19604 6452
rect 19559 6412 19604 6440
rect 18589 6403 18647 6409
rect 19598 6400 19604 6412
rect 19656 6400 19662 6452
rect 20978 6400 20984 6452
rect 21036 6440 21042 6452
rect 21073 6443 21131 6449
rect 21073 6440 21085 6443
rect 21036 6412 21085 6440
rect 21036 6400 21042 6412
rect 21073 6409 21085 6412
rect 21119 6440 21131 6443
rect 21165 6443 21223 6449
rect 21165 6440 21177 6443
rect 21119 6412 21177 6440
rect 21119 6409 21131 6412
rect 21073 6403 21131 6409
rect 21165 6409 21177 6412
rect 21211 6409 21223 6443
rect 21165 6403 21223 6409
rect 23005 6443 23063 6449
rect 23005 6409 23017 6443
rect 23051 6440 23063 6443
rect 23646 6440 23652 6452
rect 23051 6412 23652 6440
rect 23051 6409 23063 6412
rect 23005 6403 23063 6409
rect 23646 6400 23652 6412
rect 23704 6400 23710 6452
rect 24566 6440 24572 6452
rect 24527 6412 24572 6440
rect 24566 6400 24572 6412
rect 24624 6400 24630 6452
rect 15093 6375 15151 6381
rect 15093 6341 15105 6375
rect 15139 6372 15151 6375
rect 15274 6372 15280 6384
rect 15139 6344 15280 6372
rect 15139 6341 15151 6344
rect 15093 6335 15151 6341
rect 15274 6332 15280 6344
rect 15332 6372 15338 6384
rect 15332 6344 17436 6372
rect 15332 6332 15338 6344
rect 11965 6307 12023 6313
rect 11965 6273 11977 6307
rect 12011 6304 12023 6307
rect 12054 6304 12060 6316
rect 12011 6276 12060 6304
rect 12011 6273 12023 6276
rect 11965 6267 12023 6273
rect 12054 6264 12060 6276
rect 12112 6264 12118 6316
rect 13253 6307 13311 6313
rect 13253 6273 13265 6307
rect 13299 6304 13311 6307
rect 13342 6304 13348 6316
rect 13299 6276 13348 6304
rect 13299 6273 13311 6276
rect 13253 6267 13311 6273
rect 13342 6264 13348 6276
rect 13400 6264 13406 6316
rect 14173 6307 14231 6313
rect 14173 6273 14185 6307
rect 14219 6304 14231 6307
rect 14262 6304 14268 6316
rect 14219 6276 14268 6304
rect 14219 6273 14231 6276
rect 14173 6267 14231 6273
rect 14262 6264 14268 6276
rect 14320 6264 14326 6316
rect 16010 6304 16016 6316
rect 15971 6276 16016 6304
rect 16010 6264 16016 6276
rect 16068 6264 16074 6316
rect 16286 6304 16292 6316
rect 16247 6276 16292 6304
rect 16286 6264 16292 6276
rect 16344 6264 16350 6316
rect 12327 6171 12385 6177
rect 12327 6168 12339 6171
rect 11704 6140 12339 6168
rect 10456 6131 10504 6137
rect 12327 6137 12339 6140
rect 12373 6168 12385 6171
rect 13066 6168 13072 6180
rect 12373 6140 13072 6168
rect 12373 6137 12385 6140
rect 12327 6131 12385 6137
rect 10456 6128 10462 6131
rect 13066 6128 13072 6140
rect 13124 6168 13130 6180
rect 14081 6171 14139 6177
rect 14081 6168 14093 6171
rect 13124 6140 14093 6168
rect 13124 6128 13130 6140
rect 14081 6137 14093 6140
rect 14127 6168 14139 6171
rect 14535 6171 14593 6177
rect 14535 6168 14547 6171
rect 14127 6140 14547 6168
rect 14127 6137 14139 6140
rect 14081 6131 14139 6137
rect 14535 6137 14547 6140
rect 14581 6168 14593 6171
rect 15182 6168 15188 6180
rect 14581 6140 15188 6168
rect 14581 6137 14593 6140
rect 14535 6131 14593 6137
rect 15182 6128 15188 6140
rect 15240 6128 15246 6180
rect 16105 6171 16163 6177
rect 16105 6137 16117 6171
rect 16151 6168 16163 6171
rect 16378 6168 16384 6180
rect 16151 6140 16384 6168
rect 16151 6137 16163 6140
rect 16105 6131 16163 6137
rect 8834 6100 8840 6112
rect 8795 6072 8840 6100
rect 8834 6060 8840 6072
rect 8892 6060 8898 6112
rect 10674 6060 10680 6112
rect 10732 6100 10738 6112
rect 11045 6103 11103 6109
rect 11045 6100 11057 6103
rect 10732 6072 11057 6100
rect 10732 6060 10738 6072
rect 11045 6069 11057 6072
rect 11091 6069 11103 6103
rect 11045 6063 11103 6069
rect 11413 6103 11471 6109
rect 11413 6069 11425 6103
rect 11459 6100 11471 6103
rect 11686 6100 11692 6112
rect 11459 6072 11692 6100
rect 11459 6069 11471 6072
rect 11413 6063 11471 6069
rect 11686 6060 11692 6072
rect 11744 6060 11750 6112
rect 12885 6103 12943 6109
rect 12885 6069 12897 6103
rect 12931 6100 12943 6103
rect 13250 6100 13256 6112
rect 12931 6072 13256 6100
rect 12931 6069 12943 6072
rect 12885 6063 12943 6069
rect 13250 6060 13256 6072
rect 13308 6060 13314 6112
rect 15461 6103 15519 6109
rect 15461 6069 15473 6103
rect 15507 6100 15519 6103
rect 15829 6103 15887 6109
rect 15829 6100 15841 6103
rect 15507 6072 15841 6100
rect 15507 6069 15519 6072
rect 15461 6063 15519 6069
rect 15829 6069 15841 6072
rect 15875 6100 15887 6103
rect 16120 6100 16148 6131
rect 16378 6128 16384 6140
rect 16436 6128 16442 6180
rect 17408 6109 17436 6344
rect 17666 6304 17672 6316
rect 17627 6276 17672 6304
rect 17666 6264 17672 6276
rect 17724 6264 17730 6316
rect 18126 6304 18132 6316
rect 18087 6276 18132 6304
rect 18126 6264 18132 6276
rect 18184 6264 18190 6316
rect 22637 6307 22695 6313
rect 22637 6304 22649 6307
rect 20260 6276 22649 6304
rect 19598 6196 19604 6248
rect 19656 6236 19662 6248
rect 19785 6239 19843 6245
rect 19785 6236 19797 6239
rect 19656 6208 19797 6236
rect 19656 6196 19662 6208
rect 19785 6205 19797 6208
rect 19831 6205 19843 6239
rect 19785 6199 19843 6205
rect 19874 6196 19880 6248
rect 19932 6236 19938 6248
rect 20260 6245 20288 6276
rect 22637 6273 22649 6276
rect 22683 6304 22695 6307
rect 22683 6276 23692 6304
rect 22683 6273 22695 6276
rect 22637 6267 22695 6273
rect 20245 6239 20303 6245
rect 20245 6236 20257 6239
rect 19932 6208 20257 6236
rect 19932 6196 19938 6208
rect 20245 6205 20257 6208
rect 20291 6205 20303 6239
rect 20245 6199 20303 6205
rect 20889 6239 20947 6245
rect 20889 6205 20901 6239
rect 20935 6236 20947 6239
rect 21349 6239 21407 6245
rect 21349 6236 21361 6239
rect 20935 6208 21361 6236
rect 20935 6205 20947 6208
rect 20889 6199 20947 6205
rect 21349 6205 21361 6208
rect 21395 6236 21407 6239
rect 23186 6236 23192 6248
rect 21395 6208 23048 6236
rect 23147 6208 23192 6236
rect 21395 6205 21407 6208
rect 21349 6199 21407 6205
rect 17761 6171 17819 6177
rect 17761 6137 17773 6171
rect 17807 6137 17819 6171
rect 17761 6131 17819 6137
rect 20521 6171 20579 6177
rect 20521 6137 20533 6171
rect 20567 6168 20579 6171
rect 20978 6168 20984 6180
rect 20567 6140 20984 6168
rect 20567 6137 20579 6140
rect 20521 6131 20579 6137
rect 15875 6072 16148 6100
rect 17393 6103 17451 6109
rect 15875 6069 15887 6072
rect 15829 6063 15887 6069
rect 17393 6069 17405 6103
rect 17439 6100 17451 6103
rect 17776 6100 17804 6131
rect 20978 6128 20984 6140
rect 21036 6128 21042 6180
rect 21711 6171 21769 6177
rect 21711 6137 21723 6171
rect 21757 6137 21769 6171
rect 23020 6168 23048 6208
rect 23186 6196 23192 6208
rect 23244 6196 23250 6248
rect 23664 6245 23692 6276
rect 23649 6239 23707 6245
rect 23649 6205 23661 6239
rect 23695 6205 23707 6239
rect 24750 6236 24756 6248
rect 24711 6208 24756 6236
rect 23649 6199 23707 6205
rect 24750 6196 24756 6208
rect 24808 6236 24814 6248
rect 25305 6239 25363 6245
rect 25305 6236 25317 6239
rect 24808 6208 25317 6236
rect 24808 6196 24814 6208
rect 25305 6205 25317 6208
rect 25351 6205 25363 6239
rect 25305 6199 25363 6205
rect 23020 6140 23324 6168
rect 21711 6131 21769 6137
rect 17439 6072 17804 6100
rect 17439 6069 17451 6072
rect 17393 6063 17451 6069
rect 20794 6060 20800 6112
rect 20852 6100 20858 6112
rect 21073 6103 21131 6109
rect 21073 6100 21085 6103
rect 20852 6072 21085 6100
rect 20852 6060 20858 6072
rect 21073 6069 21085 6072
rect 21119 6100 21131 6103
rect 21732 6100 21760 6131
rect 21898 6100 21904 6112
rect 21119 6072 21904 6100
rect 21119 6069 21131 6072
rect 21073 6063 21131 6069
rect 21898 6060 21904 6072
rect 21956 6060 21962 6112
rect 22266 6100 22272 6112
rect 22227 6072 22272 6100
rect 22266 6060 22272 6072
rect 22324 6060 22330 6112
rect 23296 6109 23324 6140
rect 23281 6103 23339 6109
rect 23281 6069 23293 6103
rect 23327 6069 23339 6103
rect 23281 6063 23339 6069
rect 23738 6060 23744 6112
rect 23796 6100 23802 6112
rect 24937 6103 24995 6109
rect 24937 6100 24949 6103
rect 23796 6072 24949 6100
rect 23796 6060 23802 6072
rect 24937 6069 24949 6072
rect 24983 6069 24995 6103
rect 24937 6063 24995 6069
rect 632 6010 26392 6032
rect 632 5958 9843 6010
rect 9895 5958 9907 6010
rect 9959 5958 9971 6010
rect 10023 5958 10035 6010
rect 10087 5958 19176 6010
rect 19228 5958 19240 6010
rect 19292 5958 19304 6010
rect 19356 5958 19368 6010
rect 19420 5958 26392 6010
rect 632 5936 26392 5958
rect 10490 5896 10496 5908
rect 10451 5868 10496 5896
rect 10490 5856 10496 5868
rect 10548 5856 10554 5908
rect 10858 5896 10864 5908
rect 10819 5868 10864 5896
rect 10858 5856 10864 5868
rect 10916 5896 10922 5908
rect 11870 5896 11876 5908
rect 10916 5868 11876 5896
rect 10916 5856 10922 5868
rect 11870 5856 11876 5868
rect 11928 5856 11934 5908
rect 12054 5856 12060 5908
rect 12112 5896 12118 5908
rect 12609 5899 12667 5905
rect 12609 5896 12621 5899
rect 12112 5868 12621 5896
rect 12112 5856 12118 5868
rect 12609 5865 12621 5868
rect 12655 5865 12667 5899
rect 14262 5896 14268 5908
rect 14223 5868 14268 5896
rect 12609 5859 12667 5865
rect 14262 5856 14268 5868
rect 14320 5856 14326 5908
rect 16010 5896 16016 5908
rect 15971 5868 16016 5896
rect 16010 5856 16016 5868
rect 16068 5856 16074 5908
rect 17666 5896 17672 5908
rect 17627 5868 17672 5896
rect 17666 5856 17672 5868
rect 17724 5856 17730 5908
rect 18034 5896 18040 5908
rect 17995 5868 18040 5896
rect 18034 5856 18040 5868
rect 18092 5856 18098 5908
rect 18770 5856 18776 5908
rect 18828 5896 18834 5908
rect 19233 5899 19291 5905
rect 19233 5896 19245 5899
rect 18828 5868 19245 5896
rect 18828 5856 18834 5868
rect 19233 5865 19245 5868
rect 19279 5896 19291 5899
rect 20521 5899 20579 5905
rect 20521 5896 20533 5899
rect 19279 5868 20533 5896
rect 19279 5865 19291 5868
rect 19233 5859 19291 5865
rect 20521 5865 20533 5868
rect 20567 5865 20579 5899
rect 20521 5859 20579 5865
rect 21533 5899 21591 5905
rect 21533 5865 21545 5899
rect 21579 5896 21591 5899
rect 21622 5896 21628 5908
rect 21579 5868 21628 5896
rect 21579 5865 21591 5868
rect 21533 5859 21591 5865
rect 21622 5856 21628 5868
rect 21680 5856 21686 5908
rect 22450 5856 22456 5908
rect 22508 5896 22514 5908
rect 22508 5868 23968 5896
rect 22508 5856 22514 5868
rect 9202 5788 9208 5840
rect 9260 5828 9266 5840
rect 9665 5831 9723 5837
rect 9665 5828 9677 5831
rect 9260 5800 9677 5828
rect 9260 5788 9266 5800
rect 9665 5797 9677 5800
rect 9711 5828 9723 5831
rect 10030 5828 10036 5840
rect 9711 5800 10036 5828
rect 9711 5797 9723 5800
rect 9665 5791 9723 5797
rect 10030 5788 10036 5800
rect 10088 5828 10094 5840
rect 10766 5828 10772 5840
rect 10088 5800 10772 5828
rect 10088 5788 10094 5800
rect 10766 5788 10772 5800
rect 10824 5788 10830 5840
rect 11410 5837 11416 5840
rect 11407 5828 11416 5837
rect 11371 5800 11416 5828
rect 11407 5791 11416 5800
rect 11410 5788 11416 5791
rect 11468 5788 11474 5840
rect 12146 5788 12152 5840
rect 12204 5828 12210 5840
rect 12241 5831 12299 5837
rect 12241 5828 12253 5831
rect 12204 5800 12253 5828
rect 12204 5788 12210 5800
rect 12241 5797 12253 5800
rect 12287 5797 12299 5831
rect 12241 5791 12299 5797
rect 13069 5831 13127 5837
rect 13069 5797 13081 5831
rect 13115 5828 13127 5831
rect 13250 5828 13256 5840
rect 13115 5800 13256 5828
rect 13115 5797 13127 5800
rect 13069 5791 13127 5797
rect 13250 5788 13256 5800
rect 13308 5788 13314 5840
rect 15182 5837 15188 5840
rect 15179 5828 15188 5837
rect 15143 5800 15188 5828
rect 15179 5791 15188 5800
rect 15182 5788 15188 5791
rect 15240 5788 15246 5840
rect 16746 5828 16752 5840
rect 16707 5800 16752 5828
rect 16746 5788 16752 5800
rect 16804 5788 16810 5840
rect 19598 5828 19604 5840
rect 18420 5800 19604 5828
rect 6442 5720 6448 5772
rect 6500 5760 6506 5772
rect 6572 5763 6630 5769
rect 6572 5760 6584 5763
rect 6500 5732 6584 5760
rect 6500 5720 6506 5732
rect 6572 5729 6584 5732
rect 6618 5729 6630 5763
rect 6572 5723 6630 5729
rect 7638 5720 7644 5772
rect 7696 5760 7702 5772
rect 8190 5760 8196 5772
rect 7696 5732 8196 5760
rect 7696 5720 7702 5732
rect 8190 5720 8196 5732
rect 8248 5720 8254 5772
rect 11042 5760 11048 5772
rect 11003 5732 11048 5760
rect 11042 5720 11048 5732
rect 11100 5720 11106 5772
rect 14354 5720 14360 5772
rect 14412 5760 14418 5772
rect 14814 5760 14820 5772
rect 14412 5732 14820 5760
rect 14412 5720 14418 5732
rect 14814 5720 14820 5732
rect 14872 5720 14878 5772
rect 17850 5720 17856 5772
rect 17908 5760 17914 5772
rect 18420 5769 18448 5800
rect 19598 5788 19604 5800
rect 19656 5788 19662 5840
rect 19874 5828 19880 5840
rect 19835 5800 19880 5828
rect 19874 5788 19880 5800
rect 19932 5788 19938 5840
rect 20245 5831 20303 5837
rect 20245 5797 20257 5831
rect 20291 5828 20303 5831
rect 20334 5828 20340 5840
rect 20291 5800 20340 5828
rect 20291 5797 20303 5800
rect 20245 5791 20303 5797
rect 20334 5788 20340 5800
rect 20392 5788 20398 5840
rect 20610 5788 20616 5840
rect 20668 5828 20674 5840
rect 21346 5828 21352 5840
rect 20668 5800 21352 5828
rect 20668 5788 20674 5800
rect 21346 5788 21352 5800
rect 21404 5828 21410 5840
rect 21809 5831 21867 5837
rect 21809 5828 21821 5831
rect 21404 5800 21821 5828
rect 21404 5788 21410 5800
rect 21809 5797 21821 5800
rect 21855 5797 21867 5831
rect 21809 5791 21867 5797
rect 21898 5788 21904 5840
rect 21956 5828 21962 5840
rect 22314 5831 22372 5837
rect 22314 5828 22326 5831
rect 21956 5800 22326 5828
rect 21956 5788 21962 5800
rect 22314 5797 22326 5800
rect 22360 5797 22372 5831
rect 23186 5828 23192 5840
rect 23147 5800 23192 5828
rect 22314 5791 22372 5797
rect 23186 5788 23192 5800
rect 23244 5788 23250 5840
rect 23940 5837 23968 5868
rect 23925 5831 23983 5837
rect 23925 5797 23937 5831
rect 23971 5828 23983 5831
rect 24474 5828 24480 5840
rect 23971 5800 24480 5828
rect 23971 5797 23983 5800
rect 23925 5791 23983 5797
rect 24474 5788 24480 5800
rect 24532 5788 24538 5840
rect 18405 5763 18463 5769
rect 18405 5760 18417 5763
rect 17908 5732 18417 5760
rect 17908 5720 17914 5732
rect 18405 5729 18417 5732
rect 18451 5729 18463 5763
rect 18586 5760 18592 5772
rect 18547 5732 18592 5760
rect 18405 5723 18463 5729
rect 18586 5720 18592 5732
rect 18644 5720 18650 5772
rect 19966 5720 19972 5772
rect 20024 5760 20030 5772
rect 20429 5763 20487 5769
rect 20429 5760 20441 5763
rect 20024 5732 20441 5760
rect 20024 5720 20030 5732
rect 20429 5729 20441 5732
rect 20475 5760 20487 5763
rect 20702 5760 20708 5772
rect 20475 5732 20708 5760
rect 20475 5729 20487 5732
rect 20429 5723 20487 5729
rect 20702 5720 20708 5732
rect 20760 5720 20766 5772
rect 20889 5763 20947 5769
rect 20889 5729 20901 5763
rect 20935 5729 20947 5763
rect 20889 5723 20947 5729
rect 8285 5695 8343 5701
rect 8285 5661 8297 5695
rect 8331 5692 8343 5695
rect 8926 5692 8932 5704
rect 8331 5664 8932 5692
rect 8331 5661 8343 5664
rect 8285 5655 8343 5661
rect 8926 5652 8932 5664
rect 8984 5652 8990 5704
rect 9294 5652 9300 5704
rect 9352 5692 9358 5704
rect 9573 5695 9631 5701
rect 9573 5692 9585 5695
rect 9352 5664 9585 5692
rect 9352 5652 9358 5664
rect 9573 5661 9585 5664
rect 9619 5661 9631 5695
rect 9573 5655 9631 5661
rect 9754 5652 9760 5704
rect 9812 5692 9818 5704
rect 9849 5695 9907 5701
rect 9849 5692 9861 5695
rect 9812 5664 9861 5692
rect 9812 5652 9818 5664
rect 9849 5661 9861 5664
rect 9895 5661 9907 5695
rect 9849 5655 9907 5661
rect 12977 5695 13035 5701
rect 12977 5661 12989 5695
rect 13023 5692 13035 5695
rect 13158 5692 13164 5704
rect 13023 5664 13164 5692
rect 13023 5661 13035 5664
rect 12977 5655 13035 5661
rect 13158 5652 13164 5664
rect 13216 5652 13222 5704
rect 13342 5692 13348 5704
rect 13303 5664 13348 5692
rect 13342 5652 13348 5664
rect 13400 5652 13406 5704
rect 16654 5692 16660 5704
rect 16615 5664 16660 5692
rect 16654 5652 16660 5664
rect 16712 5652 16718 5704
rect 16933 5695 16991 5701
rect 16933 5661 16945 5695
rect 16979 5661 16991 5695
rect 18678 5692 18684 5704
rect 18639 5664 18684 5692
rect 16933 5655 16991 5661
rect 6675 5627 6733 5633
rect 6675 5593 6687 5627
rect 6721 5624 6733 5627
rect 7730 5624 7736 5636
rect 6721 5596 7736 5624
rect 6721 5593 6733 5596
rect 6675 5587 6733 5593
rect 7730 5584 7736 5596
rect 7788 5584 7794 5636
rect 16286 5584 16292 5636
rect 16344 5624 16350 5636
rect 16948 5624 16976 5655
rect 18678 5652 18684 5664
rect 18736 5652 18742 5704
rect 20242 5652 20248 5704
rect 20300 5692 20306 5704
rect 20904 5692 20932 5723
rect 20978 5720 20984 5772
rect 21036 5760 21042 5772
rect 21036 5732 22036 5760
rect 21036 5720 21042 5732
rect 22008 5701 22036 5732
rect 23094 5720 23100 5772
rect 23152 5760 23158 5772
rect 23557 5763 23615 5769
rect 23557 5760 23569 5763
rect 23152 5732 23569 5760
rect 23152 5720 23158 5732
rect 23557 5729 23569 5732
rect 23603 5729 23615 5763
rect 23557 5723 23615 5729
rect 20300 5664 20932 5692
rect 21993 5695 22051 5701
rect 20300 5652 20306 5664
rect 21993 5661 22005 5695
rect 22039 5692 22051 5695
rect 22082 5692 22088 5704
rect 22039 5664 22088 5692
rect 22039 5661 22051 5664
rect 21993 5655 22051 5661
rect 22082 5652 22088 5664
rect 22140 5652 22146 5704
rect 23002 5652 23008 5704
rect 23060 5692 23066 5704
rect 23833 5695 23891 5701
rect 23833 5692 23845 5695
rect 23060 5664 23845 5692
rect 23060 5652 23066 5664
rect 23833 5661 23845 5664
rect 23879 5692 23891 5695
rect 24290 5692 24296 5704
rect 23879 5664 24296 5692
rect 23879 5661 23891 5664
rect 23833 5655 23891 5661
rect 24290 5652 24296 5664
rect 24348 5652 24354 5704
rect 24382 5624 24388 5636
rect 16344 5596 16976 5624
rect 24343 5596 24388 5624
rect 16344 5584 16350 5596
rect 24382 5584 24388 5596
rect 24440 5584 24446 5636
rect 11965 5559 12023 5565
rect 11965 5525 11977 5559
rect 12011 5556 12023 5559
rect 12238 5556 12244 5568
rect 12011 5528 12244 5556
rect 12011 5525 12023 5528
rect 11965 5519 12023 5525
rect 12238 5516 12244 5528
rect 12296 5516 12302 5568
rect 15550 5516 15556 5568
rect 15608 5556 15614 5568
rect 15737 5559 15795 5565
rect 15737 5556 15749 5559
rect 15608 5528 15749 5556
rect 15608 5516 15614 5528
rect 15737 5525 15749 5528
rect 15783 5525 15795 5559
rect 22910 5556 22916 5568
rect 22871 5528 22916 5556
rect 15737 5519 15795 5525
rect 22910 5516 22916 5528
rect 22968 5516 22974 5568
rect 632 5466 26392 5488
rect 632 5414 5176 5466
rect 5228 5414 5240 5466
rect 5292 5414 5304 5466
rect 5356 5414 5368 5466
rect 5420 5414 14510 5466
rect 14562 5414 14574 5466
rect 14626 5414 14638 5466
rect 14690 5414 14702 5466
rect 14754 5414 23843 5466
rect 23895 5414 23907 5466
rect 23959 5414 23971 5466
rect 24023 5414 24035 5466
rect 24087 5414 26392 5466
rect 632 5392 26392 5414
rect 6169 5355 6227 5361
rect 6169 5321 6181 5355
rect 6215 5352 6227 5355
rect 6442 5352 6448 5364
rect 6215 5324 6448 5352
rect 6215 5321 6227 5324
rect 6169 5315 6227 5321
rect 6442 5312 6448 5324
rect 6500 5312 6506 5364
rect 7365 5355 7423 5361
rect 7365 5321 7377 5355
rect 7411 5352 7423 5355
rect 7638 5352 7644 5364
rect 7411 5324 7644 5352
rect 7411 5321 7423 5324
rect 7365 5315 7423 5321
rect 7638 5312 7644 5324
rect 7696 5312 7702 5364
rect 8834 5352 8840 5364
rect 8795 5324 8840 5352
rect 8834 5312 8840 5324
rect 8892 5312 8898 5364
rect 10030 5352 10036 5364
rect 9991 5324 10036 5352
rect 10030 5312 10036 5324
rect 10088 5312 10094 5364
rect 11042 5312 11048 5364
rect 11100 5352 11106 5364
rect 11689 5355 11747 5361
rect 11689 5352 11701 5355
rect 11100 5324 11701 5352
rect 11100 5312 11106 5324
rect 11689 5321 11701 5324
rect 11735 5321 11747 5355
rect 11689 5315 11747 5321
rect 14173 5355 14231 5361
rect 14173 5321 14185 5355
rect 14219 5352 14231 5355
rect 14354 5352 14360 5364
rect 14219 5324 14360 5352
rect 14219 5321 14231 5324
rect 14173 5315 14231 5321
rect 14354 5312 14360 5324
rect 14412 5312 14418 5364
rect 16746 5312 16752 5364
rect 16804 5352 16810 5364
rect 16933 5355 16991 5361
rect 16933 5352 16945 5355
rect 16804 5324 16945 5352
rect 16804 5312 16810 5324
rect 16933 5321 16945 5324
rect 16979 5321 16991 5355
rect 17850 5352 17856 5364
rect 17811 5324 17856 5352
rect 16933 5315 16991 5321
rect 17850 5312 17856 5324
rect 17908 5312 17914 5364
rect 18586 5312 18592 5364
rect 18644 5352 18650 5364
rect 20061 5355 20119 5361
rect 20061 5352 20073 5355
rect 18644 5324 20073 5352
rect 18644 5312 18650 5324
rect 20061 5321 20073 5324
rect 20107 5352 20119 5355
rect 20242 5352 20248 5364
rect 20107 5324 20248 5352
rect 20107 5321 20119 5324
rect 20061 5315 20119 5321
rect 20242 5312 20248 5324
rect 20300 5312 20306 5364
rect 20521 5355 20579 5361
rect 20521 5321 20533 5355
rect 20567 5352 20579 5355
rect 20794 5352 20800 5364
rect 20567 5324 20800 5352
rect 20567 5321 20579 5324
rect 20521 5315 20579 5321
rect 20794 5312 20800 5324
rect 20852 5312 20858 5364
rect 24290 5312 24296 5364
rect 24348 5312 24354 5364
rect 24474 5352 24480 5364
rect 24435 5324 24480 5352
rect 24474 5312 24480 5324
rect 24532 5312 24538 5364
rect 9294 5244 9300 5296
rect 9352 5284 9358 5296
rect 10401 5287 10459 5293
rect 10401 5284 10413 5287
rect 9352 5256 10413 5284
rect 9352 5244 9358 5256
rect 10401 5253 10413 5256
rect 10447 5253 10459 5287
rect 10401 5247 10459 5253
rect 16565 5287 16623 5293
rect 16565 5253 16577 5287
rect 16611 5284 16623 5287
rect 17022 5284 17028 5296
rect 16611 5256 17028 5284
rect 16611 5253 16623 5256
rect 16565 5247 16623 5253
rect 17022 5244 17028 5256
rect 17080 5244 17086 5296
rect 19785 5287 19843 5293
rect 19785 5253 19797 5287
rect 19831 5284 19843 5287
rect 19966 5284 19972 5296
rect 19831 5256 19972 5284
rect 19831 5253 19843 5256
rect 19785 5247 19843 5253
rect 19966 5244 19972 5256
rect 20024 5244 20030 5296
rect 24308 5284 24336 5312
rect 24845 5287 24903 5293
rect 24845 5284 24857 5287
rect 24308 5256 24857 5284
rect 24845 5253 24857 5256
rect 24891 5253 24903 5287
rect 24845 5247 24903 5253
rect 6445 5219 6503 5225
rect 6445 5185 6457 5219
rect 6491 5216 6503 5219
rect 6534 5216 6540 5228
rect 6491 5188 6540 5216
rect 6491 5185 6503 5188
rect 6445 5179 6503 5185
rect 6534 5176 6540 5188
rect 6592 5176 6598 5228
rect 9754 5216 9760 5228
rect 9715 5188 9760 5216
rect 9754 5176 9760 5188
rect 9812 5216 9818 5228
rect 10306 5216 10312 5228
rect 9812 5188 10312 5216
rect 9812 5176 9818 5188
rect 10306 5176 10312 5188
rect 10364 5176 10370 5228
rect 12330 5176 12336 5228
rect 12388 5216 12394 5228
rect 12517 5219 12575 5225
rect 12517 5216 12529 5219
rect 12388 5188 12529 5216
rect 12388 5176 12394 5188
rect 12517 5185 12529 5188
rect 12563 5185 12575 5219
rect 12517 5179 12575 5185
rect 15182 5176 15188 5228
rect 15240 5216 15246 5228
rect 15737 5219 15795 5225
rect 15737 5216 15749 5219
rect 15240 5188 15749 5216
rect 15240 5176 15246 5188
rect 15737 5185 15749 5188
rect 15783 5216 15795 5219
rect 15783 5188 16608 5216
rect 15783 5185 15795 5188
rect 15737 5179 15795 5185
rect 6997 5151 7055 5157
rect 6997 5117 7009 5151
rect 7043 5148 7055 5151
rect 8098 5148 8104 5160
rect 7043 5120 8104 5148
rect 7043 5117 7055 5120
rect 6997 5111 7055 5117
rect 8098 5108 8104 5120
rect 8156 5108 8162 5160
rect 10912 5151 10970 5157
rect 10912 5117 10924 5151
rect 10958 5148 10970 5151
rect 11778 5148 11784 5160
rect 10958 5120 11784 5148
rect 10958 5117 10970 5120
rect 10912 5111 10970 5117
rect 11778 5108 11784 5120
rect 11836 5108 11842 5160
rect 14541 5151 14599 5157
rect 14541 5117 14553 5151
rect 14587 5148 14599 5151
rect 15274 5148 15280 5160
rect 14587 5120 15280 5148
rect 14587 5117 14599 5120
rect 14541 5111 14599 5117
rect 15274 5108 15280 5120
rect 15332 5108 15338 5160
rect 16381 5151 16439 5157
rect 16381 5148 16393 5151
rect 16212 5120 16393 5148
rect 8190 5080 8196 5092
rect 8151 5052 8196 5080
rect 8190 5040 8196 5052
rect 8248 5040 8254 5092
rect 9113 5083 9171 5089
rect 9113 5080 9125 5083
rect 8484 5052 9125 5080
rect 8484 5024 8512 5052
rect 9113 5049 9125 5052
rect 9159 5049 9171 5083
rect 9113 5043 9171 5049
rect 9205 5083 9263 5089
rect 9205 5049 9217 5083
rect 9251 5049 9263 5083
rect 9205 5043 9263 5049
rect 10999 5083 11057 5089
rect 10999 5049 11011 5083
rect 11045 5080 11057 5083
rect 11962 5080 11968 5092
rect 11045 5052 11968 5080
rect 11045 5049 11057 5052
rect 10999 5043 11057 5049
rect 8466 5012 8472 5024
rect 8427 4984 8472 5012
rect 8466 4972 8472 4984
rect 8524 4972 8530 5024
rect 8834 4972 8840 5024
rect 8892 5012 8898 5024
rect 9220 5012 9248 5043
rect 11962 5040 11968 5052
rect 12020 5040 12026 5092
rect 12425 5083 12483 5089
rect 12425 5049 12437 5083
rect 12471 5080 12483 5083
rect 12879 5083 12937 5089
rect 12879 5080 12891 5083
rect 12471 5052 12891 5080
rect 12471 5049 12483 5052
rect 12425 5043 12483 5049
rect 12879 5049 12891 5052
rect 12925 5080 12937 5083
rect 13066 5080 13072 5092
rect 12925 5052 13072 5080
rect 12925 5049 12937 5052
rect 12879 5043 12937 5049
rect 8892 4984 9248 5012
rect 8892 4972 8898 4984
rect 11318 4972 11324 5024
rect 11376 5012 11382 5024
rect 11413 5015 11471 5021
rect 11413 5012 11425 5015
rect 11376 4984 11425 5012
rect 11376 4972 11382 4984
rect 11413 4981 11425 4984
rect 11459 5012 11471 5015
rect 12440 5012 12468 5043
rect 13066 5040 13072 5052
rect 13124 5040 13130 5092
rect 13250 5040 13256 5092
rect 13308 5080 13314 5092
rect 14630 5080 14636 5092
rect 13308 5052 13756 5080
rect 14591 5052 14636 5080
rect 13308 5040 13314 5052
rect 13728 5024 13756 5052
rect 14630 5040 14636 5052
rect 14688 5040 14694 5092
rect 11459 4984 12468 5012
rect 13437 5015 13495 5021
rect 11459 4981 11471 4984
rect 11413 4975 11471 4981
rect 13437 4981 13449 5015
rect 13483 5012 13495 5015
rect 13526 5012 13532 5024
rect 13483 4984 13532 5012
rect 13483 4981 13495 4984
rect 13437 4975 13495 4981
rect 13526 4972 13532 4984
rect 13584 4972 13590 5024
rect 13710 5012 13716 5024
rect 13671 4984 13716 5012
rect 13710 4972 13716 4984
rect 13768 4972 13774 5024
rect 16102 4972 16108 5024
rect 16160 5012 16166 5024
rect 16212 5021 16240 5120
rect 16381 5117 16393 5120
rect 16427 5117 16439 5151
rect 16580 5148 16608 5188
rect 16654 5176 16660 5228
rect 16712 5216 16718 5228
rect 17301 5219 17359 5225
rect 17301 5216 17313 5219
rect 16712 5188 17313 5216
rect 16712 5176 16718 5188
rect 17301 5185 17313 5188
rect 17347 5185 17359 5219
rect 17301 5179 17359 5185
rect 18313 5219 18371 5225
rect 18313 5185 18325 5219
rect 18359 5216 18371 5219
rect 18770 5216 18776 5228
rect 18359 5188 18776 5216
rect 18359 5185 18371 5188
rect 18313 5179 18371 5185
rect 18770 5176 18776 5188
rect 18828 5176 18834 5228
rect 20242 5176 20248 5228
rect 20300 5216 20306 5228
rect 20613 5219 20671 5225
rect 20613 5216 20625 5219
rect 20300 5188 20625 5216
rect 20300 5176 20306 5188
rect 20613 5185 20625 5188
rect 20659 5216 20671 5219
rect 22361 5219 22419 5225
rect 22361 5216 22373 5219
rect 20659 5188 22373 5216
rect 20659 5185 20671 5188
rect 20613 5179 20671 5185
rect 22361 5185 22373 5188
rect 22407 5185 22419 5219
rect 22361 5179 22419 5185
rect 23370 5176 23376 5228
rect 23428 5216 23434 5228
rect 23557 5219 23615 5225
rect 23557 5216 23569 5219
rect 23428 5188 23569 5216
rect 23428 5176 23434 5188
rect 23557 5185 23569 5188
rect 23603 5216 23615 5219
rect 24290 5216 24296 5228
rect 23603 5188 24296 5216
rect 23603 5185 23615 5188
rect 23557 5179 23615 5185
rect 24290 5176 24296 5188
rect 24348 5176 24354 5228
rect 19233 5151 19291 5157
rect 16580 5120 16976 5148
rect 16381 5111 16439 5117
rect 16948 5092 16976 5120
rect 19233 5117 19245 5151
rect 19279 5148 19291 5151
rect 19966 5148 19972 5160
rect 19279 5120 19972 5148
rect 19279 5117 19291 5120
rect 19233 5111 19291 5117
rect 19966 5108 19972 5120
rect 20024 5108 20030 5160
rect 25026 5148 25032 5160
rect 24987 5120 25032 5148
rect 25026 5108 25032 5120
rect 25084 5148 25090 5160
rect 25581 5151 25639 5157
rect 25581 5148 25593 5151
rect 25084 5120 25593 5148
rect 25084 5108 25090 5120
rect 25581 5117 25593 5120
rect 25627 5117 25639 5151
rect 25581 5111 25639 5117
rect 16930 5040 16936 5092
rect 16988 5080 16994 5092
rect 18221 5083 18279 5089
rect 18221 5080 18233 5083
rect 16988 5052 18233 5080
rect 16988 5040 16994 5052
rect 18221 5049 18233 5052
rect 18267 5080 18279 5083
rect 18675 5083 18733 5089
rect 18675 5080 18687 5083
rect 18267 5052 18687 5080
rect 18267 5049 18279 5052
rect 18221 5043 18279 5049
rect 18675 5049 18687 5052
rect 18721 5080 18733 5083
rect 18770 5080 18776 5092
rect 18721 5052 18776 5080
rect 18721 5049 18733 5052
rect 18675 5043 18733 5049
rect 18770 5040 18776 5052
rect 18828 5040 18834 5092
rect 20794 5040 20800 5092
rect 20852 5080 20858 5092
rect 20934 5083 20992 5089
rect 20934 5080 20946 5083
rect 20852 5052 20946 5080
rect 20852 5040 20858 5052
rect 20934 5049 20946 5052
rect 20980 5080 20992 5083
rect 21993 5083 22051 5089
rect 21993 5080 22005 5083
rect 20980 5052 22005 5080
rect 20980 5049 20992 5052
rect 20934 5043 20992 5049
rect 21993 5049 22005 5052
rect 22039 5049 22051 5083
rect 23649 5083 23707 5089
rect 23649 5080 23661 5083
rect 21993 5043 22051 5049
rect 23020 5052 23661 5080
rect 23020 5024 23048 5052
rect 23649 5049 23661 5052
rect 23695 5049 23707 5083
rect 23649 5043 23707 5049
rect 24201 5083 24259 5089
rect 24201 5049 24213 5083
rect 24247 5080 24259 5083
rect 24290 5080 24296 5092
rect 24247 5052 24296 5080
rect 24247 5049 24259 5052
rect 24201 5043 24259 5049
rect 24290 5040 24296 5052
rect 24348 5040 24354 5092
rect 16197 5015 16255 5021
rect 16197 5012 16209 5015
rect 16160 4984 16209 5012
rect 16160 4972 16166 4984
rect 16197 4981 16209 4984
rect 16243 4981 16255 5015
rect 21530 5012 21536 5024
rect 21491 4984 21536 5012
rect 16197 4975 16255 4981
rect 21530 4972 21536 4984
rect 21588 4972 21594 5024
rect 23002 5012 23008 5024
rect 22963 4984 23008 5012
rect 23002 4972 23008 4984
rect 23060 4972 23066 5024
rect 25210 5012 25216 5024
rect 25171 4984 25216 5012
rect 25210 4972 25216 4984
rect 25268 4972 25274 5024
rect 632 4922 26392 4944
rect 632 4870 9843 4922
rect 9895 4870 9907 4922
rect 9959 4870 9971 4922
rect 10023 4870 10035 4922
rect 10087 4870 19176 4922
rect 19228 4870 19240 4922
rect 19292 4870 19304 4922
rect 19356 4870 19368 4922
rect 19420 4870 26392 4922
rect 632 4848 26392 4870
rect 5663 4811 5721 4817
rect 5663 4777 5675 4811
rect 5709 4808 5721 4811
rect 5798 4808 5804 4820
rect 5709 4780 5804 4808
rect 5709 4777 5721 4780
rect 5663 4771 5721 4777
rect 5798 4768 5804 4780
rect 5856 4768 5862 4820
rect 10306 4808 10312 4820
rect 10267 4780 10312 4808
rect 10306 4768 10312 4780
rect 10364 4768 10370 4820
rect 11778 4808 11784 4820
rect 11739 4780 11784 4808
rect 11778 4768 11784 4780
rect 11836 4768 11842 4820
rect 12330 4768 12336 4820
rect 12388 4808 12394 4820
rect 12517 4811 12575 4817
rect 12517 4808 12529 4811
rect 12388 4780 12529 4808
rect 12388 4768 12394 4780
rect 12517 4777 12529 4780
rect 12563 4777 12575 4811
rect 12517 4771 12575 4777
rect 12977 4811 13035 4817
rect 12977 4777 12989 4811
rect 13023 4808 13035 4811
rect 13158 4808 13164 4820
rect 13023 4780 13164 4808
rect 13023 4777 13035 4780
rect 12977 4771 13035 4777
rect 13158 4768 13164 4780
rect 13216 4768 13222 4820
rect 18221 4811 18279 4817
rect 18221 4777 18233 4811
rect 18267 4808 18279 4811
rect 18586 4808 18592 4820
rect 18267 4780 18592 4808
rect 18267 4777 18279 4780
rect 18221 4771 18279 4777
rect 18586 4768 18592 4780
rect 18644 4768 18650 4820
rect 21346 4808 21352 4820
rect 21307 4780 21352 4808
rect 21346 4768 21352 4780
rect 21404 4768 21410 4820
rect 22082 4808 22088 4820
rect 22043 4780 22088 4808
rect 22082 4768 22088 4780
rect 22140 4768 22146 4820
rect 23370 4808 23376 4820
rect 23331 4780 23376 4808
rect 23370 4768 23376 4780
rect 23428 4768 23434 4820
rect 10855 4743 10913 4749
rect 10855 4709 10867 4743
rect 10901 4740 10913 4743
rect 11318 4740 11324 4752
rect 10901 4712 11324 4740
rect 10901 4709 10913 4712
rect 10855 4703 10913 4709
rect 11318 4700 11324 4712
rect 11376 4700 11382 4752
rect 13345 4743 13403 4749
rect 13345 4709 13357 4743
rect 13391 4740 13403 4743
rect 13434 4740 13440 4752
rect 13391 4712 13440 4740
rect 13391 4709 13403 4712
rect 13345 4703 13403 4709
rect 13434 4700 13440 4712
rect 13492 4740 13498 4752
rect 14630 4740 14636 4752
rect 13492 4712 14636 4740
rect 13492 4700 13498 4712
rect 14630 4700 14636 4712
rect 14688 4700 14694 4752
rect 16559 4743 16617 4749
rect 16559 4709 16571 4743
rect 16605 4740 16617 4743
rect 16930 4740 16936 4752
rect 16605 4712 16936 4740
rect 16605 4709 16617 4712
rect 16559 4703 16617 4709
rect 16930 4700 16936 4712
rect 16988 4700 16994 4752
rect 18770 4700 18776 4752
rect 18828 4740 18834 4752
rect 20794 4749 20800 4752
rect 18951 4743 19009 4749
rect 18951 4740 18963 4743
rect 18828 4712 18963 4740
rect 18828 4700 18834 4712
rect 18951 4709 18963 4712
rect 18997 4740 19009 4743
rect 20791 4740 20800 4749
rect 18997 4712 20800 4740
rect 18997 4709 19009 4712
rect 18951 4703 19009 4709
rect 20791 4703 20800 4712
rect 20794 4700 20800 4703
rect 20852 4700 20858 4752
rect 23646 4740 23652 4752
rect 23607 4712 23652 4740
rect 23646 4700 23652 4712
rect 23704 4700 23710 4752
rect 4580 4675 4638 4681
rect 4580 4641 4592 4675
rect 4626 4672 4638 4675
rect 4786 4672 4792 4684
rect 4626 4644 4792 4672
rect 4626 4641 4638 4644
rect 4580 4635 4638 4641
rect 4786 4632 4792 4644
rect 4844 4632 4850 4684
rect 5592 4675 5650 4681
rect 5592 4641 5604 4675
rect 5638 4672 5650 4675
rect 5706 4672 5712 4684
rect 5638 4644 5712 4672
rect 5638 4641 5650 4644
rect 5592 4635 5650 4641
rect 5706 4632 5712 4644
rect 5764 4632 5770 4684
rect 8190 4672 8196 4684
rect 8151 4644 8196 4672
rect 8190 4632 8196 4644
rect 8248 4632 8254 4684
rect 9478 4672 9484 4684
rect 9439 4644 9484 4672
rect 9478 4632 9484 4644
rect 9536 4632 9542 4684
rect 10490 4672 10496 4684
rect 10451 4644 10496 4672
rect 10490 4632 10496 4644
rect 10548 4632 10554 4684
rect 15090 4672 15096 4684
rect 15051 4644 15096 4672
rect 15090 4632 15096 4644
rect 15148 4632 15154 4684
rect 16194 4672 16200 4684
rect 16155 4644 16200 4672
rect 16194 4632 16200 4644
rect 16252 4632 16258 4684
rect 18589 4675 18647 4681
rect 18589 4641 18601 4675
rect 18635 4672 18647 4675
rect 18678 4672 18684 4684
rect 18635 4644 18684 4672
rect 18635 4641 18647 4644
rect 18589 4635 18647 4641
rect 18678 4632 18684 4644
rect 18736 4632 18742 4684
rect 20242 4632 20248 4684
rect 20300 4672 20306 4684
rect 20429 4675 20487 4681
rect 20429 4672 20441 4675
rect 20300 4644 20441 4672
rect 20300 4632 20306 4644
rect 20429 4641 20441 4644
rect 20475 4641 20487 4675
rect 22174 4672 22180 4684
rect 22135 4644 22180 4672
rect 20429 4635 20487 4641
rect 22174 4632 22180 4644
rect 22232 4672 22238 4684
rect 22729 4675 22787 4681
rect 22729 4672 22741 4675
rect 22232 4644 22741 4672
rect 22232 4632 22238 4644
rect 22729 4641 22741 4644
rect 22775 4641 22787 4675
rect 22729 4635 22787 4641
rect 6534 4604 6540 4616
rect 6495 4576 6540 4604
rect 6534 4564 6540 4576
rect 6592 4564 6598 4616
rect 8285 4607 8343 4613
rect 8285 4573 8297 4607
rect 8331 4604 8343 4607
rect 9110 4604 9116 4616
rect 8331 4576 9116 4604
rect 8331 4573 8343 4576
rect 8285 4567 8343 4573
rect 9110 4564 9116 4576
rect 9168 4564 9174 4616
rect 13250 4604 13256 4616
rect 13211 4576 13256 4604
rect 13250 4564 13256 4576
rect 13308 4564 13314 4616
rect 13894 4604 13900 4616
rect 13855 4576 13900 4604
rect 13894 4564 13900 4576
rect 13952 4564 13958 4616
rect 23186 4564 23192 4616
rect 23244 4604 23250 4616
rect 23557 4607 23615 4613
rect 23557 4604 23569 4607
rect 23244 4576 23569 4604
rect 23244 4564 23250 4576
rect 23557 4573 23569 4576
rect 23603 4573 23615 4607
rect 23557 4567 23615 4573
rect 24201 4607 24259 4613
rect 24201 4573 24213 4607
rect 24247 4604 24259 4607
rect 24290 4604 24296 4616
rect 24247 4576 24296 4604
rect 24247 4573 24259 4576
rect 24201 4567 24259 4573
rect 24290 4564 24296 4576
rect 24348 4564 24354 4616
rect 4651 4539 4709 4545
rect 4651 4505 4663 4539
rect 4697 4536 4709 4539
rect 4970 4536 4976 4548
rect 4697 4508 4976 4536
rect 4697 4505 4709 4508
rect 4651 4499 4709 4505
rect 4970 4496 4976 4508
rect 5028 4496 5034 4548
rect 21714 4496 21720 4548
rect 21772 4536 21778 4548
rect 22361 4539 22419 4545
rect 22361 4536 22373 4539
rect 21772 4508 22373 4536
rect 21772 4496 21778 4508
rect 22361 4505 22373 4508
rect 22407 4505 22419 4539
rect 22361 4499 22419 4505
rect 11410 4468 11416 4480
rect 11371 4440 11416 4468
rect 11410 4428 11416 4440
rect 11468 4428 11474 4480
rect 15274 4468 15280 4480
rect 15235 4440 15280 4468
rect 15274 4428 15280 4440
rect 15332 4428 15338 4480
rect 17114 4468 17120 4480
rect 17075 4440 17120 4468
rect 17114 4428 17120 4440
rect 17172 4428 17178 4480
rect 17482 4428 17488 4480
rect 17540 4468 17546 4480
rect 17577 4471 17635 4477
rect 17577 4468 17589 4471
rect 17540 4440 17589 4468
rect 17540 4428 17546 4440
rect 17577 4437 17589 4440
rect 17623 4437 17635 4471
rect 19506 4468 19512 4480
rect 19467 4440 19512 4468
rect 17577 4431 17635 4437
rect 19506 4428 19512 4440
rect 19564 4428 19570 4480
rect 632 4378 26392 4400
rect 632 4326 5176 4378
rect 5228 4326 5240 4378
rect 5292 4326 5304 4378
rect 5356 4326 5368 4378
rect 5420 4326 14510 4378
rect 14562 4326 14574 4378
rect 14626 4326 14638 4378
rect 14690 4326 14702 4378
rect 14754 4326 23843 4378
rect 23895 4326 23907 4378
rect 23959 4326 23971 4378
rect 24023 4326 24035 4378
rect 24087 4326 26392 4378
rect 632 4304 26392 4326
rect 11318 4264 11324 4276
rect 11279 4236 11324 4264
rect 11318 4224 11324 4236
rect 11376 4224 11382 4276
rect 13434 4264 13440 4276
rect 13395 4236 13440 4264
rect 13434 4224 13440 4236
rect 13492 4224 13498 4276
rect 16749 4267 16807 4273
rect 16749 4233 16761 4267
rect 16795 4264 16807 4267
rect 16930 4264 16936 4276
rect 16795 4236 16936 4264
rect 16795 4233 16807 4236
rect 16749 4227 16807 4233
rect 16930 4224 16936 4236
rect 16988 4224 16994 4276
rect 18589 4267 18647 4273
rect 18589 4233 18601 4267
rect 18635 4264 18647 4267
rect 18770 4264 18776 4276
rect 18635 4236 18776 4264
rect 18635 4233 18647 4236
rect 18589 4227 18647 4233
rect 18770 4224 18776 4236
rect 18828 4224 18834 4276
rect 20242 4224 20248 4276
rect 20300 4264 20306 4276
rect 20889 4267 20947 4273
rect 20889 4264 20901 4267
rect 20300 4236 20901 4264
rect 20300 4224 20306 4236
rect 20889 4233 20901 4236
rect 20935 4233 20947 4267
rect 21346 4264 21352 4276
rect 21307 4236 21352 4264
rect 20889 4227 20947 4233
rect 21346 4224 21352 4236
rect 21404 4224 21410 4276
rect 23646 4224 23652 4276
rect 23704 4264 23710 4276
rect 24201 4267 24259 4273
rect 24201 4264 24213 4267
rect 23704 4236 24213 4264
rect 23704 4224 23710 4236
rect 24201 4233 24213 4236
rect 24247 4233 24259 4267
rect 24201 4227 24259 4233
rect 8190 4196 8196 4208
rect 7840 4168 8196 4196
rect 7641 4131 7699 4137
rect 7641 4097 7653 4131
rect 7687 4128 7699 4131
rect 7840 4128 7868 4168
rect 8190 4156 8196 4168
rect 8248 4196 8254 4208
rect 8248 4168 9156 4196
rect 8248 4156 8254 4168
rect 7687 4100 7868 4128
rect 9128 4128 9156 4168
rect 10306 4156 10312 4208
rect 10364 4196 10370 4208
rect 10364 4168 10444 4196
rect 10364 4156 10370 4168
rect 10416 4137 10444 4168
rect 18678 4156 18684 4208
rect 18736 4196 18742 4208
rect 20613 4199 20671 4205
rect 18736 4168 18816 4196
rect 18736 4156 18742 4168
rect 10401 4131 10459 4137
rect 9128 4100 10260 4128
rect 7687 4097 7699 4100
rect 7641 4091 7699 4097
rect 3292 4063 3350 4069
rect 3292 4029 3304 4063
rect 3338 4060 3350 4063
rect 4304 4063 4362 4069
rect 3338 4032 3820 4060
rect 3338 4029 3350 4032
rect 3292 4023 3350 4029
rect 3363 3927 3421 3933
rect 3363 3893 3375 3927
rect 3409 3924 3421 3927
rect 3590 3924 3596 3936
rect 3409 3896 3596 3924
rect 3409 3893 3421 3896
rect 3363 3887 3421 3893
rect 3590 3884 3596 3896
rect 3648 3884 3654 3936
rect 3792 3933 3820 4032
rect 4304 4029 4316 4063
rect 4350 4060 4362 4063
rect 5316 4063 5374 4069
rect 4350 4032 5200 4060
rect 4350 4029 4362 4032
rect 4304 4023 4362 4029
rect 5172 4001 5200 4032
rect 5316 4029 5328 4063
rect 5362 4060 5374 4063
rect 5522 4060 5528 4072
rect 5362 4032 5528 4060
rect 5362 4029 5374 4032
rect 5316 4023 5374 4029
rect 5522 4020 5528 4032
rect 5580 4060 5586 4072
rect 6077 4063 6135 4069
rect 6077 4060 6089 4063
rect 5580 4032 6089 4060
rect 5580 4020 5586 4032
rect 6077 4029 6089 4032
rect 6123 4029 6135 4063
rect 6077 4023 6135 4029
rect 7546 4020 7552 4072
rect 7604 4060 7610 4072
rect 7733 4063 7791 4069
rect 7733 4060 7745 4063
rect 7604 4032 7745 4060
rect 7604 4020 7610 4032
rect 7733 4029 7745 4032
rect 7779 4029 7791 4063
rect 7733 4023 7791 4029
rect 8653 4063 8711 4069
rect 8653 4029 8665 4063
rect 8699 4060 8711 4063
rect 9110 4060 9116 4072
rect 8699 4032 9116 4060
rect 8699 4029 8711 4032
rect 8653 4023 8711 4029
rect 9110 4020 9116 4032
rect 9168 4020 9174 4072
rect 5157 3995 5215 4001
rect 5157 3961 5169 3995
rect 5203 3992 5215 3995
rect 5890 3992 5896 4004
rect 5203 3964 5896 3992
rect 5203 3961 5215 3964
rect 5157 3955 5215 3961
rect 5890 3952 5896 3964
rect 5948 3952 5954 4004
rect 10232 4001 10260 4100
rect 10401 4097 10413 4131
rect 10447 4097 10459 4131
rect 12422 4128 12428 4140
rect 12383 4100 12428 4128
rect 10401 4091 10459 4097
rect 12422 4088 12428 4100
rect 12480 4088 12486 4140
rect 13069 4131 13127 4137
rect 13069 4097 13081 4131
rect 13115 4128 13127 4131
rect 13342 4128 13348 4140
rect 13115 4100 13348 4128
rect 13115 4097 13127 4100
rect 13069 4091 13127 4097
rect 13342 4088 13348 4100
rect 13400 4128 13406 4140
rect 13989 4131 14047 4137
rect 13989 4128 14001 4131
rect 13400 4100 14001 4128
rect 13400 4088 13406 4100
rect 13989 4097 14001 4100
rect 14035 4128 14047 4131
rect 14170 4128 14176 4140
rect 14035 4100 14176 4128
rect 14035 4097 14047 4100
rect 13989 4091 14047 4097
rect 14170 4088 14176 4100
rect 14228 4088 14234 4140
rect 14262 4088 14268 4140
rect 14320 4128 14326 4140
rect 15550 4128 15556 4140
rect 14320 4100 14365 4128
rect 15511 4100 15556 4128
rect 14320 4088 14326 4100
rect 15550 4088 15556 4100
rect 15608 4128 15614 4140
rect 15608 4100 15780 4128
rect 15608 4088 15614 4100
rect 15752 4069 15780 4100
rect 16194 4088 16200 4140
rect 16252 4128 16258 4140
rect 17945 4131 18003 4137
rect 17945 4128 17957 4131
rect 16252 4100 17957 4128
rect 16252 4088 16258 4100
rect 17945 4097 17957 4100
rect 17991 4097 18003 4131
rect 18788 4128 18816 4168
rect 20613 4165 20625 4199
rect 20659 4196 20671 4199
rect 20794 4196 20800 4208
rect 20659 4168 20800 4196
rect 20659 4165 20671 4168
rect 20613 4159 20671 4165
rect 20794 4156 20800 4168
rect 20852 4156 20858 4208
rect 21438 4156 21444 4208
rect 21496 4156 21502 4208
rect 23186 4196 23192 4208
rect 22928 4168 23192 4196
rect 18957 4131 19015 4137
rect 18957 4128 18969 4131
rect 18788 4100 18969 4128
rect 17945 4091 18003 4097
rect 18957 4097 18969 4100
rect 19003 4097 19015 4131
rect 18957 4091 19015 4097
rect 19690 4088 19696 4140
rect 19748 4128 19754 4140
rect 19877 4131 19935 4137
rect 19877 4128 19889 4131
rect 19748 4100 19889 4128
rect 19748 4088 19754 4100
rect 19877 4097 19889 4100
rect 19923 4097 19935 4131
rect 21456 4128 21484 4156
rect 21533 4131 21591 4137
rect 21533 4128 21545 4131
rect 21456 4100 21545 4128
rect 19877 4091 19935 4097
rect 21533 4097 21545 4100
rect 21579 4097 21591 4131
rect 21533 4091 21591 4097
rect 21898 4088 21904 4140
rect 21956 4128 21962 4140
rect 22545 4131 22603 4137
rect 22545 4128 22557 4131
rect 21956 4100 22557 4128
rect 21956 4088 21962 4100
rect 22545 4097 22557 4100
rect 22591 4128 22603 4131
rect 22928 4128 22956 4168
rect 23186 4156 23192 4168
rect 23244 4156 23250 4208
rect 22591 4100 22956 4128
rect 23005 4131 23063 4137
rect 22591 4097 22603 4100
rect 22545 4091 22603 4097
rect 23005 4097 23017 4131
rect 23051 4128 23063 4131
rect 23370 4128 23376 4140
rect 23051 4100 23376 4128
rect 23051 4097 23063 4100
rect 23005 4091 23063 4097
rect 23370 4088 23376 4100
rect 23428 4088 23434 4140
rect 23462 4088 23468 4140
rect 23520 4128 23526 4140
rect 23557 4131 23615 4137
rect 23557 4128 23569 4131
rect 23520 4100 23569 4128
rect 23520 4088 23526 4100
rect 23557 4097 23569 4100
rect 23603 4097 23615 4131
rect 23557 4091 23615 4097
rect 15737 4063 15795 4069
rect 15737 4029 15749 4063
rect 15783 4029 15795 4063
rect 24750 4060 24756 4072
rect 24711 4032 24756 4060
rect 15737 4023 15795 4029
rect 24750 4020 24756 4032
rect 24808 4060 24814 4072
rect 25305 4063 25363 4069
rect 25305 4060 25317 4063
rect 24808 4032 25317 4060
rect 24808 4020 24814 4032
rect 25305 4029 25317 4032
rect 25351 4029 25363 4063
rect 25305 4023 25363 4029
rect 10217 3995 10275 4001
rect 10217 3961 10229 3995
rect 10263 3992 10275 3995
rect 10493 3995 10551 4001
rect 10493 3992 10505 3995
rect 10263 3964 10505 3992
rect 10263 3961 10275 3964
rect 10217 3955 10275 3961
rect 10493 3961 10505 3964
rect 10539 3992 10551 3995
rect 10674 3992 10680 4004
rect 10539 3964 10680 3992
rect 10539 3961 10551 3964
rect 10493 3955 10551 3961
rect 10674 3952 10680 3964
rect 10732 3952 10738 4004
rect 11045 3995 11103 4001
rect 11045 3961 11057 3995
rect 11091 3961 11103 3995
rect 12146 3992 12152 4004
rect 12107 3964 12152 3992
rect 11045 3955 11103 3961
rect 3777 3927 3835 3933
rect 3777 3893 3789 3927
rect 3823 3924 3835 3927
rect 4142 3924 4148 3936
rect 3823 3896 4148 3924
rect 3823 3893 3835 3896
rect 3777 3887 3835 3893
rect 4142 3884 4148 3896
rect 4200 3884 4206 3936
rect 4375 3927 4433 3933
rect 4375 3893 4387 3927
rect 4421 3924 4433 3927
rect 4602 3924 4608 3936
rect 4421 3896 4608 3924
rect 4421 3893 4433 3896
rect 4375 3887 4433 3893
rect 4602 3884 4608 3896
rect 4660 3884 4666 3936
rect 4786 3924 4792 3936
rect 4747 3896 4792 3924
rect 4786 3884 4792 3896
rect 4844 3884 4850 3936
rect 5387 3927 5445 3933
rect 5387 3893 5399 3927
rect 5433 3924 5445 3927
rect 5614 3924 5620 3936
rect 5433 3896 5620 3924
rect 5433 3893 5445 3896
rect 5387 3887 5445 3893
rect 5614 3884 5620 3896
rect 5672 3884 5678 3936
rect 5706 3884 5712 3936
rect 5764 3924 5770 3936
rect 6718 3924 6724 3936
rect 5764 3896 5809 3924
rect 6679 3896 6724 3924
rect 5764 3884 5770 3896
rect 6718 3884 6724 3896
rect 6776 3884 6782 3936
rect 9018 3924 9024 3936
rect 8979 3896 9024 3924
rect 9018 3884 9024 3896
rect 9076 3884 9082 3936
rect 10306 3884 10312 3936
rect 10364 3924 10370 3936
rect 11060 3924 11088 3955
rect 12146 3952 12152 3964
rect 12204 3952 12210 4004
rect 12517 3995 12575 4001
rect 12517 3961 12529 3995
rect 12563 3961 12575 3995
rect 12517 3955 12575 3961
rect 14081 3995 14139 4001
rect 14081 3961 14093 3995
rect 14127 3961 14139 3995
rect 14081 3955 14139 3961
rect 16381 3995 16439 4001
rect 16381 3961 16393 3995
rect 16427 3992 16439 3995
rect 17301 3995 17359 4001
rect 17301 3992 17313 3995
rect 16427 3964 17313 3992
rect 16427 3961 16439 3964
rect 16381 3955 16439 3961
rect 17301 3961 17313 3964
rect 17347 3961 17359 3995
rect 17301 3955 17359 3961
rect 10364 3896 11088 3924
rect 12164 3924 12192 3952
rect 12532 3924 12560 3955
rect 12164 3896 12560 3924
rect 10364 3884 10370 3896
rect 13526 3884 13532 3936
rect 13584 3924 13590 3936
rect 13713 3927 13771 3933
rect 13713 3924 13725 3927
rect 13584 3896 13725 3924
rect 13584 3884 13590 3896
rect 13713 3893 13725 3896
rect 13759 3924 13771 3927
rect 14096 3924 14124 3955
rect 13759 3896 14124 3924
rect 13759 3893 13771 3896
rect 13713 3887 13771 3893
rect 14814 3884 14820 3936
rect 14872 3924 14878 3936
rect 14909 3927 14967 3933
rect 14909 3924 14921 3927
rect 14872 3896 14921 3924
rect 14872 3884 14878 3896
rect 14909 3893 14921 3896
rect 14955 3893 14967 3927
rect 17316 3924 17344 3955
rect 17482 3952 17488 4004
rect 17540 3992 17546 4004
rect 17669 3995 17727 4001
rect 17669 3992 17681 3995
rect 17540 3964 17681 3992
rect 17540 3952 17546 3964
rect 17669 3961 17681 3964
rect 17715 3961 17727 3995
rect 17669 3955 17727 3961
rect 17761 3995 17819 4001
rect 17761 3961 17773 3995
rect 17807 3961 17819 3995
rect 17761 3955 17819 3961
rect 17776 3924 17804 3955
rect 19046 3952 19052 4004
rect 19104 3992 19110 4004
rect 19601 3995 19659 4001
rect 19601 3992 19613 3995
rect 19104 3964 19613 3992
rect 19104 3952 19110 3964
rect 19601 3961 19613 3964
rect 19647 3961 19659 3995
rect 19601 3955 19659 3961
rect 19693 3995 19751 4001
rect 19693 3961 19705 3995
rect 19739 3961 19751 3995
rect 19693 3955 19751 3961
rect 17316 3896 17804 3924
rect 19417 3927 19475 3933
rect 14909 3887 14967 3893
rect 19417 3893 19429 3927
rect 19463 3924 19475 3927
rect 19506 3924 19512 3936
rect 19463 3896 19512 3924
rect 19463 3893 19475 3896
rect 19417 3887 19475 3893
rect 19506 3884 19512 3896
rect 19564 3924 19570 3936
rect 19708 3924 19736 3955
rect 21346 3952 21352 4004
rect 21404 3992 21410 4004
rect 21625 3995 21683 4001
rect 21625 3992 21637 3995
rect 21404 3964 21637 3992
rect 21404 3952 21410 3964
rect 21625 3961 21637 3964
rect 21671 3961 21683 3995
rect 21625 3955 21683 3961
rect 22177 3995 22235 4001
rect 22177 3961 22189 3995
rect 22223 3992 22235 3995
rect 22450 3992 22456 4004
rect 22223 3964 22456 3992
rect 22223 3961 22235 3964
rect 22177 3955 22235 3961
rect 22450 3952 22456 3964
rect 22508 3952 22514 4004
rect 23281 3995 23339 4001
rect 23281 3992 23293 3995
rect 23204 3964 23293 3992
rect 23204 3936 23232 3964
rect 23281 3961 23293 3964
rect 23327 3961 23339 3995
rect 23281 3955 23339 3961
rect 23370 3952 23376 4004
rect 23428 3992 23434 4004
rect 23428 3964 23473 3992
rect 23428 3952 23434 3964
rect 20150 3924 20156 3936
rect 19564 3896 20156 3924
rect 19564 3884 19570 3896
rect 20150 3884 20156 3896
rect 20208 3884 20214 3936
rect 23186 3884 23192 3936
rect 23244 3884 23250 3936
rect 24934 3924 24940 3936
rect 24895 3896 24940 3924
rect 24934 3884 24940 3896
rect 24992 3884 24998 3936
rect 632 3834 26392 3856
rect 632 3782 9843 3834
rect 9895 3782 9907 3834
rect 9959 3782 9971 3834
rect 10023 3782 10035 3834
rect 10087 3782 19176 3834
rect 19228 3782 19240 3834
rect 19292 3782 19304 3834
rect 19356 3782 19368 3834
rect 19420 3782 26392 3834
rect 632 3760 26392 3782
rect 4050 3729 4056 3732
rect 4007 3723 4056 3729
rect 4007 3689 4019 3723
rect 4053 3689 4056 3723
rect 4007 3683 4056 3689
rect 4050 3680 4056 3683
rect 4108 3680 4114 3732
rect 6074 3729 6080 3732
rect 6031 3723 6080 3729
rect 6031 3689 6043 3723
rect 6077 3689 6080 3723
rect 6031 3683 6080 3689
rect 6074 3680 6080 3683
rect 6132 3680 6138 3732
rect 8055 3723 8113 3729
rect 8055 3689 8067 3723
rect 8101 3720 8113 3723
rect 8374 3720 8380 3732
rect 8101 3692 8380 3720
rect 8101 3689 8113 3692
rect 8055 3683 8113 3689
rect 8374 3680 8380 3692
rect 8432 3680 8438 3732
rect 10582 3680 10588 3732
rect 10640 3720 10646 3732
rect 10677 3723 10735 3729
rect 10677 3720 10689 3723
rect 10640 3692 10689 3720
rect 10640 3680 10646 3692
rect 10677 3689 10689 3692
rect 10723 3689 10735 3723
rect 12422 3720 12428 3732
rect 12383 3692 12428 3720
rect 10677 3683 10735 3689
rect 12422 3680 12428 3692
rect 12480 3680 12486 3732
rect 14170 3720 14176 3732
rect 14131 3692 14176 3720
rect 14170 3680 14176 3692
rect 14228 3680 14234 3732
rect 15090 3680 15096 3732
rect 15148 3720 15154 3732
rect 15277 3723 15335 3729
rect 15277 3720 15289 3723
rect 15148 3692 15289 3720
rect 15148 3680 15154 3692
rect 15277 3689 15289 3692
rect 15323 3689 15335 3723
rect 15277 3683 15335 3689
rect 16286 3680 16292 3732
rect 16344 3720 16350 3732
rect 16841 3723 16899 3729
rect 16841 3720 16853 3723
rect 16344 3692 16853 3720
rect 16344 3680 16350 3692
rect 16841 3689 16853 3692
rect 16887 3689 16899 3723
rect 16841 3683 16899 3689
rect 19966 3680 19972 3732
rect 20024 3720 20030 3732
rect 20426 3720 20432 3732
rect 20024 3692 20432 3720
rect 20024 3680 20030 3692
rect 20426 3680 20432 3692
rect 20484 3720 20490 3732
rect 21438 3720 21444 3732
rect 20484 3692 20656 3720
rect 21399 3692 21444 3720
rect 20484 3680 20490 3692
rect 9202 3612 9208 3664
rect 9260 3652 9266 3664
rect 9849 3655 9907 3661
rect 9849 3652 9861 3655
rect 9260 3624 9861 3652
rect 9260 3612 9266 3624
rect 9849 3621 9861 3624
rect 9895 3652 9907 3655
rect 10122 3652 10128 3664
rect 9895 3624 10128 3652
rect 9895 3621 9907 3624
rect 9849 3615 9907 3621
rect 10122 3612 10128 3624
rect 10180 3612 10186 3664
rect 11318 3612 11324 3664
rect 11376 3652 11382 3664
rect 11413 3655 11471 3661
rect 11413 3652 11425 3655
rect 11376 3624 11425 3652
rect 11376 3612 11382 3624
rect 11413 3621 11425 3624
rect 11459 3621 11471 3655
rect 11413 3615 11471 3621
rect 15550 3612 15556 3664
rect 15608 3652 15614 3664
rect 16013 3655 16071 3661
rect 16013 3652 16025 3655
rect 15608 3624 16025 3652
rect 15608 3612 15614 3624
rect 16013 3621 16025 3624
rect 16059 3621 16071 3655
rect 16013 3615 16071 3621
rect 17114 3612 17120 3664
rect 17172 3652 17178 3664
rect 17577 3655 17635 3661
rect 17577 3652 17589 3655
rect 17172 3624 17589 3652
rect 17172 3612 17178 3624
rect 17577 3621 17589 3624
rect 17623 3621 17635 3655
rect 17577 3615 17635 3621
rect 20245 3655 20303 3661
rect 20245 3621 20257 3655
rect 20291 3652 20303 3655
rect 20518 3652 20524 3664
rect 20291 3624 20524 3652
rect 20291 3621 20303 3624
rect 20245 3615 20303 3621
rect 20518 3612 20524 3624
rect 20576 3612 20582 3664
rect 20628 3661 20656 3692
rect 21438 3680 21444 3692
rect 21496 3680 21502 3732
rect 23554 3680 23560 3732
rect 23612 3680 23618 3732
rect 20613 3655 20671 3661
rect 20613 3621 20625 3655
rect 20659 3621 20671 3655
rect 22174 3652 22180 3664
rect 22135 3624 22180 3652
rect 20613 3615 20671 3621
rect 22174 3612 22180 3624
rect 22232 3612 22238 3664
rect 23572 3652 23600 3680
rect 23741 3655 23799 3661
rect 23741 3652 23753 3655
rect 23572 3624 23753 3652
rect 23741 3621 23753 3624
rect 23787 3621 23799 3655
rect 23741 3615 23799 3621
rect 3958 3593 3964 3596
rect 3936 3587 3964 3593
rect 3936 3553 3948 3587
rect 3936 3547 3964 3553
rect 3958 3544 3964 3547
rect 4016 3544 4022 3596
rect 4948 3587 5006 3593
rect 4948 3553 4960 3587
rect 4994 3584 5006 3587
rect 5062 3584 5068 3596
rect 4994 3556 5068 3584
rect 4994 3553 5006 3556
rect 4948 3547 5006 3553
rect 5062 3544 5068 3556
rect 5120 3544 5126 3596
rect 5982 3593 5988 3596
rect 5960 3587 5988 3593
rect 5960 3553 5972 3587
rect 5960 3547 5988 3553
rect 5982 3544 5988 3547
rect 6040 3544 6046 3596
rect 7984 3587 8042 3593
rect 7984 3553 7996 3587
rect 8030 3584 8042 3587
rect 8282 3584 8288 3596
rect 8030 3556 8288 3584
rect 8030 3553 8042 3556
rect 7984 3547 8042 3553
rect 8282 3544 8288 3556
rect 8340 3544 8346 3596
rect 13526 3584 13532 3596
rect 13487 3556 13532 3584
rect 13526 3544 13532 3556
rect 13584 3544 13590 3596
rect 14906 3593 14912 3596
rect 14884 3587 14912 3593
rect 14884 3553 14896 3587
rect 14884 3547 14912 3553
rect 14906 3544 14912 3547
rect 14964 3544 14970 3596
rect 18954 3584 18960 3596
rect 18915 3556 18960 3584
rect 18954 3544 18960 3556
rect 19012 3544 19018 3596
rect 6902 3516 6908 3528
rect 6863 3488 6908 3516
rect 6902 3476 6908 3488
rect 6960 3476 6966 3528
rect 9294 3476 9300 3528
rect 9352 3516 9358 3528
rect 9757 3519 9815 3525
rect 9757 3516 9769 3519
rect 9352 3488 9769 3516
rect 9352 3476 9358 3488
rect 9757 3485 9769 3488
rect 9803 3485 9815 3519
rect 10214 3516 10220 3528
rect 10175 3488 10220 3516
rect 9757 3479 9815 3485
rect 10214 3476 10220 3488
rect 10272 3476 10278 3528
rect 11137 3519 11195 3525
rect 11137 3485 11149 3519
rect 11183 3516 11195 3519
rect 11321 3519 11379 3525
rect 11321 3516 11333 3519
rect 11183 3488 11333 3516
rect 11183 3485 11195 3488
rect 11137 3479 11195 3485
rect 11321 3485 11333 3488
rect 11367 3516 11379 3519
rect 11594 3516 11600 3528
rect 11367 3488 11600 3516
rect 11367 3485 11379 3488
rect 11321 3479 11379 3485
rect 11594 3476 11600 3488
rect 11652 3476 11658 3528
rect 11965 3519 12023 3525
rect 11965 3485 11977 3519
rect 12011 3516 12023 3519
rect 12054 3516 12060 3528
rect 12011 3488 12060 3516
rect 12011 3485 12023 3488
rect 11965 3479 12023 3485
rect 12054 3476 12060 3488
rect 12112 3516 12118 3528
rect 12701 3519 12759 3525
rect 12701 3516 12713 3519
rect 12112 3488 12713 3516
rect 12112 3476 12118 3488
rect 12701 3485 12713 3488
rect 12747 3485 12759 3519
rect 12701 3479 12759 3485
rect 13894 3476 13900 3528
rect 13952 3516 13958 3528
rect 15921 3519 15979 3525
rect 15921 3516 15933 3519
rect 13952 3488 15933 3516
rect 13952 3476 13958 3488
rect 15921 3485 15933 3488
rect 15967 3485 15979 3519
rect 16194 3516 16200 3528
rect 16155 3488 16200 3516
rect 15921 3479 15979 3485
rect 15936 3448 15964 3479
rect 16194 3476 16200 3488
rect 16252 3476 16258 3528
rect 17301 3519 17359 3525
rect 17301 3485 17313 3519
rect 17347 3516 17359 3519
rect 17485 3519 17543 3525
rect 17485 3516 17497 3519
rect 17347 3488 17497 3516
rect 17347 3485 17359 3488
rect 17301 3479 17359 3485
rect 17485 3485 17497 3488
rect 17531 3516 17543 3519
rect 17574 3516 17580 3528
rect 17531 3488 17580 3516
rect 17531 3485 17543 3488
rect 17485 3479 17543 3485
rect 17574 3476 17580 3488
rect 17632 3476 17638 3528
rect 18126 3516 18132 3528
rect 17684 3488 18132 3516
rect 16286 3448 16292 3460
rect 15936 3420 16292 3448
rect 16286 3408 16292 3420
rect 16344 3448 16350 3460
rect 17684 3448 17712 3488
rect 18126 3476 18132 3488
rect 18184 3476 18190 3528
rect 20797 3519 20855 3525
rect 20797 3485 20809 3519
rect 20843 3485 20855 3519
rect 22082 3516 22088 3528
rect 22043 3488 22088 3516
rect 20797 3479 20855 3485
rect 18034 3448 18040 3460
rect 16344 3420 17712 3448
rect 17995 3420 18040 3448
rect 16344 3408 16350 3420
rect 18034 3408 18040 3420
rect 18092 3408 18098 3460
rect 19046 3408 19052 3460
rect 19104 3448 19110 3460
rect 19509 3451 19567 3457
rect 19509 3448 19521 3451
rect 19104 3420 19521 3448
rect 19104 3408 19110 3420
rect 19509 3417 19521 3420
rect 19555 3448 19567 3451
rect 20812 3448 20840 3479
rect 22082 3476 22088 3488
rect 22140 3476 22146 3528
rect 22358 3516 22364 3528
rect 22319 3488 22364 3516
rect 22358 3476 22364 3488
rect 22416 3476 22422 3528
rect 22450 3476 22456 3528
rect 22508 3516 22514 3528
rect 23646 3516 23652 3528
rect 22508 3488 23652 3516
rect 22508 3476 22514 3488
rect 23646 3476 23652 3488
rect 23704 3476 23710 3528
rect 23925 3519 23983 3525
rect 23925 3485 23937 3519
rect 23971 3485 23983 3519
rect 23925 3479 23983 3485
rect 19555 3420 20840 3448
rect 22376 3448 22404 3476
rect 23940 3448 23968 3479
rect 22376 3420 23968 3448
rect 19555 3417 19567 3420
rect 19509 3411 19567 3417
rect 4878 3340 4884 3392
rect 4936 3380 4942 3392
rect 5019 3383 5077 3389
rect 5019 3380 5031 3383
rect 4936 3352 5031 3380
rect 4936 3340 4942 3352
rect 5019 3349 5031 3352
rect 5065 3349 5077 3383
rect 5019 3343 5077 3349
rect 9386 3340 9392 3392
rect 9444 3380 9450 3392
rect 9481 3383 9539 3389
rect 9481 3380 9493 3383
rect 9444 3352 9493 3380
rect 9444 3340 9450 3352
rect 9481 3349 9493 3352
rect 9527 3349 9539 3383
rect 13618 3380 13624 3392
rect 13579 3352 13624 3380
rect 9481 3343 9539 3349
rect 13618 3340 13624 3352
rect 13676 3340 13682 3392
rect 14955 3383 15013 3389
rect 14955 3349 14967 3383
rect 15001 3380 15013 3383
rect 16010 3380 16016 3392
rect 15001 3352 16016 3380
rect 15001 3349 15013 3352
rect 14955 3343 15013 3349
rect 16010 3340 16016 3352
rect 16068 3340 16074 3392
rect 17666 3340 17672 3392
rect 17724 3380 17730 3392
rect 18405 3383 18463 3389
rect 18405 3380 18417 3383
rect 17724 3352 18417 3380
rect 17724 3340 17730 3352
rect 18405 3349 18417 3352
rect 18451 3349 18463 3383
rect 18405 3343 18463 3349
rect 18586 3340 18592 3392
rect 18644 3380 18650 3392
rect 19141 3383 19199 3389
rect 19141 3380 19153 3383
rect 18644 3352 19153 3380
rect 18644 3340 18650 3352
rect 19141 3349 19153 3352
rect 19187 3349 19199 3383
rect 23186 3380 23192 3392
rect 23147 3352 23192 3380
rect 19141 3343 19199 3349
rect 23186 3340 23192 3352
rect 23244 3340 23250 3392
rect 632 3290 26392 3312
rect 632 3238 5176 3290
rect 5228 3238 5240 3290
rect 5292 3238 5304 3290
rect 5356 3238 5368 3290
rect 5420 3238 14510 3290
rect 14562 3238 14574 3290
rect 14626 3238 14638 3290
rect 14690 3238 14702 3290
rect 14754 3238 23843 3290
rect 23895 3238 23907 3290
rect 23959 3238 23971 3290
rect 24023 3238 24035 3290
rect 24087 3238 26392 3290
rect 632 3216 26392 3238
rect 2762 3176 2768 3188
rect 2723 3148 2768 3176
rect 2762 3136 2768 3148
rect 2820 3136 2826 3188
rect 3406 3185 3412 3188
rect 3363 3179 3412 3185
rect 3363 3145 3375 3179
rect 3409 3145 3412 3179
rect 3363 3139 3412 3145
rect 3406 3136 3412 3139
rect 3464 3136 3470 3188
rect 3774 3176 3780 3188
rect 3735 3148 3780 3176
rect 3774 3136 3780 3148
rect 3832 3136 3838 3188
rect 3958 3136 3964 3188
rect 4016 3176 4022 3188
rect 4418 3185 4424 3188
rect 4053 3179 4111 3185
rect 4053 3176 4065 3179
rect 4016 3148 4065 3176
rect 4016 3136 4022 3148
rect 4053 3145 4065 3148
rect 4099 3145 4111 3179
rect 4053 3139 4111 3145
rect 4375 3179 4424 3185
rect 4375 3145 4387 3179
rect 4421 3145 4424 3179
rect 4375 3139 4424 3145
rect 4418 3136 4424 3139
rect 4476 3136 4482 3188
rect 5062 3176 5068 3188
rect 5023 3148 5068 3176
rect 5062 3136 5068 3148
rect 5120 3136 5126 3188
rect 5798 3176 5804 3188
rect 5759 3148 5804 3176
rect 5798 3136 5804 3148
rect 5856 3136 5862 3188
rect 5982 3136 5988 3188
rect 6040 3176 6046 3188
rect 6077 3179 6135 3185
rect 6077 3176 6089 3179
rect 6040 3148 6089 3176
rect 6040 3136 6046 3148
rect 6077 3145 6089 3148
rect 6123 3145 6135 3179
rect 6077 3139 6135 3145
rect 9205 3179 9263 3185
rect 9205 3145 9217 3179
rect 9251 3176 9263 3179
rect 9294 3176 9300 3188
rect 9251 3148 9300 3176
rect 9251 3145 9263 3148
rect 9205 3139 9263 3145
rect 9294 3136 9300 3148
rect 9352 3136 9358 3188
rect 10122 3176 10128 3188
rect 10083 3148 10128 3176
rect 10122 3136 10128 3148
rect 10180 3136 10186 3188
rect 10398 3136 10404 3188
rect 10456 3136 10462 3188
rect 11781 3179 11839 3185
rect 11781 3145 11793 3179
rect 11827 3176 11839 3179
rect 12238 3176 12244 3188
rect 11827 3148 12244 3176
rect 11827 3145 11839 3148
rect 11781 3139 11839 3145
rect 12238 3136 12244 3148
rect 12296 3176 12302 3188
rect 12422 3176 12428 3188
rect 12296 3148 12428 3176
rect 12296 3136 12302 3148
rect 12422 3136 12428 3148
rect 12480 3136 12486 3188
rect 13158 3176 13164 3188
rect 13119 3148 13164 3176
rect 13158 3136 13164 3148
rect 13216 3136 13222 3188
rect 13618 3176 13624 3188
rect 13579 3148 13624 3176
rect 13618 3136 13624 3148
rect 13676 3136 13682 3188
rect 15550 3136 15556 3188
rect 15608 3176 15614 3188
rect 15737 3179 15795 3185
rect 15737 3176 15749 3179
rect 15608 3148 15749 3176
rect 15608 3136 15614 3148
rect 15737 3145 15749 3148
rect 15783 3145 15795 3179
rect 15737 3139 15795 3145
rect 17025 3179 17083 3185
rect 17025 3145 17037 3179
rect 17071 3176 17083 3179
rect 17114 3176 17120 3188
rect 17071 3148 17120 3176
rect 17071 3145 17083 3148
rect 17025 3139 17083 3145
rect 2264 2975 2322 2981
rect 2264 2941 2276 2975
rect 2310 2972 2322 2975
rect 2762 2972 2768 2984
rect 2310 2944 2768 2972
rect 2310 2941 2322 2944
rect 2264 2935 2322 2941
rect 2762 2932 2768 2944
rect 2820 2932 2826 2984
rect 3292 2975 3350 2981
rect 3292 2941 3304 2975
rect 3338 2972 3350 2975
rect 3774 2972 3780 2984
rect 3338 2944 3780 2972
rect 3338 2941 3350 2944
rect 3292 2935 3350 2941
rect 3774 2932 3780 2944
rect 3832 2932 3838 2984
rect 4234 2932 4240 2984
rect 4292 2981 4298 2984
rect 4292 2975 4330 2981
rect 4318 2972 4330 2975
rect 4697 2975 4755 2981
rect 4697 2972 4709 2975
rect 4318 2944 4709 2972
rect 4318 2941 4330 2944
rect 4292 2935 4330 2941
rect 4697 2941 4709 2944
rect 4743 2941 4755 2975
rect 4697 2935 4755 2941
rect 5300 2975 5358 2981
rect 5300 2941 5312 2975
rect 5346 2972 5358 2975
rect 5816 2972 5844 3136
rect 9435 3111 9493 3117
rect 9435 3077 9447 3111
rect 9481 3108 9493 3111
rect 10416 3108 10444 3136
rect 9481 3080 10444 3108
rect 9481 3077 9493 3080
rect 9435 3071 9493 3077
rect 8834 3040 8840 3052
rect 8346 3012 8840 3040
rect 7178 2972 7184 2984
rect 5346 2944 5844 2972
rect 7139 2944 7184 2972
rect 5346 2941 5358 2944
rect 5300 2935 5358 2941
rect 4292 2932 4298 2935
rect 7178 2932 7184 2944
rect 7236 2972 7242 2984
rect 8346 2981 8374 3012
rect 8834 3000 8840 3012
rect 8892 3000 8898 3052
rect 9202 3000 9208 3052
rect 9260 3040 9266 3052
rect 10401 3043 10459 3049
rect 10401 3040 10413 3043
rect 9260 3012 10413 3040
rect 9260 3000 9266 3012
rect 10401 3009 10413 3012
rect 10447 3009 10459 3043
rect 10401 3003 10459 3009
rect 11045 3043 11103 3049
rect 11045 3009 11057 3043
rect 11091 3040 11103 3043
rect 12054 3040 12060 3052
rect 11091 3012 12060 3040
rect 11091 3009 11103 3012
rect 11045 3003 11103 3009
rect 12054 3000 12060 3012
rect 12112 3000 12118 3052
rect 12330 3040 12336 3052
rect 12291 3012 12336 3040
rect 12330 3000 12336 3012
rect 12388 3000 12394 3052
rect 7308 2975 7366 2981
rect 7308 2972 7320 2975
rect 7236 2944 7320 2972
rect 7236 2932 7242 2944
rect 7308 2941 7320 2944
rect 7354 2941 7366 2975
rect 7308 2935 7366 2941
rect 8331 2975 8389 2981
rect 8331 2941 8343 2975
rect 8377 2941 8389 2975
rect 8331 2935 8389 2941
rect 8423 2975 8481 2981
rect 8423 2941 8435 2975
rect 8469 2972 8481 2975
rect 9110 2972 9116 2984
rect 8469 2944 9116 2972
rect 8469 2941 8481 2944
rect 8423 2935 8481 2941
rect 9110 2932 9116 2944
rect 9168 2932 9174 2984
rect 9364 2975 9422 2981
rect 9364 2941 9376 2975
rect 9410 2972 9422 2975
rect 9410 2944 9892 2972
rect 9410 2941 9422 2944
rect 9364 2935 9422 2941
rect 2351 2907 2409 2913
rect 2351 2873 2363 2907
rect 2397 2904 2409 2907
rect 5387 2907 5445 2913
rect 2397 2876 3268 2904
rect 2397 2873 2409 2876
rect 2351 2867 2409 2873
rect 3240 2848 3268 2876
rect 5387 2873 5399 2907
rect 5433 2904 5445 2907
rect 5798 2904 5804 2916
rect 5433 2876 5804 2904
rect 5433 2873 5445 2876
rect 5387 2867 5445 2873
rect 5798 2864 5804 2876
rect 5856 2864 5862 2916
rect 9864 2913 9892 2944
rect 9849 2907 9907 2913
rect 9849 2873 9861 2907
rect 9895 2904 9907 2907
rect 10398 2904 10404 2916
rect 9895 2876 10404 2904
rect 9895 2873 9907 2876
rect 9849 2867 9907 2873
rect 10398 2864 10404 2876
rect 10456 2864 10462 2916
rect 10490 2864 10496 2916
rect 10548 2904 10554 2916
rect 12149 2907 12207 2913
rect 10548 2876 10593 2904
rect 10548 2864 10554 2876
rect 12149 2873 12161 2907
rect 12195 2904 12207 2907
rect 12422 2904 12428 2916
rect 12195 2876 12428 2904
rect 12195 2873 12207 2876
rect 12149 2867 12207 2873
rect 12422 2864 12428 2876
rect 12480 2864 12486 2916
rect 3222 2796 3228 2848
rect 3280 2796 3286 2848
rect 7411 2839 7469 2845
rect 7411 2805 7423 2839
rect 7457 2836 7469 2839
rect 7638 2836 7644 2848
rect 7457 2808 7644 2836
rect 7457 2805 7469 2808
rect 7411 2799 7469 2805
rect 7638 2796 7644 2808
rect 7696 2796 7702 2848
rect 8009 2839 8067 2845
rect 8009 2805 8021 2839
rect 8055 2836 8067 2839
rect 8282 2836 8288 2848
rect 8055 2808 8288 2836
rect 8055 2805 8067 2808
rect 8009 2799 8067 2805
rect 8282 2796 8288 2808
rect 8340 2796 8346 2848
rect 11318 2836 11324 2848
rect 11279 2808 11324 2836
rect 11318 2796 11324 2808
rect 11376 2796 11382 2848
rect 13636 2836 13664 3136
rect 13802 3040 13808 3052
rect 13763 3012 13808 3040
rect 13802 3000 13808 3012
rect 13860 3000 13866 3052
rect 14262 3040 14268 3052
rect 14223 3012 14268 3040
rect 14262 3000 14268 3012
rect 14320 3000 14326 3052
rect 15461 2975 15519 2981
rect 15461 2941 15473 2975
rect 15507 2972 15519 2975
rect 16473 2975 16531 2981
rect 16473 2972 16485 2975
rect 15507 2944 16485 2972
rect 15507 2941 15519 2944
rect 15461 2935 15519 2941
rect 16473 2941 16485 2944
rect 16519 2972 16531 2975
rect 17040 2972 17068 3139
rect 17114 3136 17120 3148
rect 17172 3136 17178 3188
rect 20337 3179 20395 3185
rect 20337 3145 20349 3179
rect 20383 3176 20395 3179
rect 20426 3176 20432 3188
rect 20383 3148 20432 3176
rect 20383 3145 20395 3148
rect 20337 3139 20395 3145
rect 20426 3136 20432 3148
rect 20484 3176 20490 3188
rect 23005 3179 23063 3185
rect 23005 3176 23017 3179
rect 20484 3148 23017 3176
rect 20484 3136 20490 3148
rect 23005 3145 23017 3148
rect 23051 3145 23063 3179
rect 23005 3139 23063 3145
rect 22082 3068 22088 3120
rect 22140 3108 22146 3120
rect 22361 3111 22419 3117
rect 22361 3108 22373 3111
rect 22140 3080 22373 3108
rect 22140 3068 22146 3080
rect 22361 3077 22373 3080
rect 22407 3077 22419 3111
rect 22361 3071 22419 3077
rect 17666 3040 17672 3052
rect 17627 3012 17672 3040
rect 17666 3000 17672 3012
rect 17724 3000 17730 3052
rect 18034 3040 18040 3052
rect 17995 3012 18040 3040
rect 18034 3000 18040 3012
rect 18092 3000 18098 3052
rect 19690 3040 19696 3052
rect 19651 3012 19696 3040
rect 19690 3000 19696 3012
rect 19748 3000 19754 3052
rect 21533 3043 21591 3049
rect 21533 3009 21545 3043
rect 21579 3040 21591 3043
rect 22450 3040 22456 3052
rect 21579 3012 22456 3040
rect 21579 3009 21591 3012
rect 21533 3003 21591 3009
rect 22450 3000 22456 3012
rect 22508 3000 22514 3052
rect 16519 2944 17068 2972
rect 23020 2972 23048 3139
rect 23646 3136 23652 3188
rect 23704 3176 23710 3188
rect 24569 3179 24627 3185
rect 24569 3176 24581 3179
rect 23704 3148 24581 3176
rect 23704 3136 23710 3148
rect 24569 3145 24581 3148
rect 24615 3145 24627 3179
rect 24934 3176 24940 3188
rect 24895 3148 24940 3176
rect 24569 3139 24627 3145
rect 24934 3136 24940 3148
rect 24992 3136 24998 3188
rect 23462 3068 23468 3120
rect 23520 3108 23526 3120
rect 24201 3111 24259 3117
rect 24201 3108 24213 3111
rect 23520 3080 24213 3108
rect 23520 3068 23526 3080
rect 24201 3077 24213 3080
rect 24247 3077 24259 3111
rect 24201 3071 24259 3077
rect 23281 2975 23339 2981
rect 23281 2972 23293 2975
rect 23020 2944 23293 2972
rect 16519 2941 16531 2944
rect 16473 2935 16531 2941
rect 23281 2941 23293 2944
rect 23327 2941 23339 2975
rect 23281 2935 23339 2941
rect 23554 2932 23560 2984
rect 23612 2972 23618 2984
rect 24198 2972 24204 2984
rect 23612 2944 24204 2972
rect 23612 2932 23618 2944
rect 24198 2932 24204 2944
rect 24256 2932 24262 2984
rect 24753 2975 24811 2981
rect 24753 2941 24765 2975
rect 24799 2972 24811 2975
rect 25210 2972 25216 2984
rect 24799 2944 25216 2972
rect 24799 2941 24811 2944
rect 24753 2935 24811 2941
rect 25210 2932 25216 2944
rect 25268 2972 25274 2984
rect 25305 2975 25363 2981
rect 25305 2972 25317 2975
rect 25268 2944 25317 2972
rect 25268 2932 25274 2944
rect 25305 2941 25317 2944
rect 25351 2941 25363 2975
rect 25305 2935 25363 2941
rect 13897 2907 13955 2913
rect 13897 2873 13909 2907
rect 13943 2873 13955 2907
rect 14906 2904 14912 2916
rect 14819 2876 14912 2904
rect 13897 2867 13955 2873
rect 13912 2836 13940 2867
rect 14906 2864 14912 2876
rect 14964 2904 14970 2916
rect 16562 2904 16568 2916
rect 14964 2876 16568 2904
rect 14964 2864 14970 2876
rect 16562 2864 16568 2876
rect 16620 2864 16626 2916
rect 16657 2907 16715 2913
rect 16657 2873 16669 2907
rect 16703 2904 16715 2907
rect 17301 2907 17359 2913
rect 17301 2904 17313 2907
rect 16703 2876 17313 2904
rect 16703 2873 16715 2876
rect 16657 2867 16715 2873
rect 17301 2873 17313 2876
rect 17347 2873 17359 2907
rect 17301 2867 17359 2873
rect 17761 2907 17819 2913
rect 17761 2873 17773 2907
rect 17807 2873 17819 2907
rect 17761 2867 17819 2873
rect 13636 2808 13940 2836
rect 17316 2836 17344 2867
rect 17776 2836 17804 2867
rect 18494 2864 18500 2916
rect 18552 2904 18558 2916
rect 18773 2907 18831 2913
rect 18773 2904 18785 2907
rect 18552 2876 18785 2904
rect 18552 2864 18558 2876
rect 18773 2873 18785 2876
rect 18819 2904 18831 2907
rect 19325 2907 19383 2913
rect 19325 2904 19337 2907
rect 18819 2876 19337 2904
rect 18819 2873 18831 2876
rect 18773 2867 18831 2873
rect 19325 2873 19337 2876
rect 19371 2873 19383 2907
rect 19325 2867 19383 2873
rect 19417 2907 19475 2913
rect 19417 2873 19429 2907
rect 19463 2904 19475 2907
rect 19690 2904 19696 2916
rect 19463 2876 19696 2904
rect 19463 2873 19475 2876
rect 19417 2867 19475 2873
rect 17316 2808 17804 2836
rect 19141 2839 19199 2845
rect 19141 2805 19153 2839
rect 19187 2836 19199 2839
rect 19432 2836 19460 2867
rect 19690 2864 19696 2876
rect 19748 2864 19754 2916
rect 20058 2864 20064 2916
rect 20116 2904 20122 2916
rect 20889 2907 20947 2913
rect 20889 2904 20901 2907
rect 20116 2876 20901 2904
rect 20116 2864 20122 2876
rect 20889 2873 20901 2876
rect 20935 2873 20947 2907
rect 20889 2867 20947 2873
rect 20981 2907 21039 2913
rect 20981 2873 20993 2907
rect 21027 2904 21039 2907
rect 21254 2904 21260 2916
rect 21027 2876 21260 2904
rect 21027 2873 21039 2876
rect 20981 2867 21039 2873
rect 19187 2808 19460 2836
rect 20705 2839 20763 2845
rect 19187 2805 19199 2808
rect 19141 2799 19199 2805
rect 20705 2805 20717 2839
rect 20751 2836 20763 2839
rect 20996 2836 21024 2867
rect 21254 2864 21260 2876
rect 21312 2864 21318 2916
rect 23002 2864 23008 2916
rect 23060 2904 23066 2916
rect 23189 2907 23247 2913
rect 23189 2904 23201 2907
rect 23060 2876 23201 2904
rect 23060 2864 23066 2876
rect 23189 2873 23201 2876
rect 23235 2873 23247 2907
rect 23189 2867 23247 2873
rect 20751 2808 21024 2836
rect 22085 2839 22143 2845
rect 20751 2805 20763 2808
rect 20705 2799 20763 2805
rect 22085 2805 22097 2839
rect 22131 2836 22143 2839
rect 22174 2836 22180 2848
rect 22131 2808 22180 2836
rect 22131 2805 22143 2808
rect 22085 2799 22143 2805
rect 22174 2796 22180 2808
rect 22232 2836 22238 2848
rect 22910 2836 22916 2848
rect 22232 2808 22916 2836
rect 22232 2796 22238 2808
rect 22910 2796 22916 2808
rect 22968 2796 22974 2848
rect 632 2746 26392 2768
rect 632 2694 9843 2746
rect 9895 2694 9907 2746
rect 9959 2694 9971 2746
rect 10023 2694 10035 2746
rect 10087 2694 19176 2746
rect 19228 2694 19240 2746
rect 19292 2694 19304 2746
rect 19356 2694 19368 2746
rect 19420 2694 26392 2746
rect 632 2672 26392 2694
rect 1658 2641 1664 2644
rect 1615 2635 1664 2641
rect 1615 2601 1627 2635
rect 1661 2601 1664 2635
rect 1615 2595 1664 2601
rect 1658 2592 1664 2595
rect 1716 2592 1722 2644
rect 4510 2641 4516 2644
rect 4467 2635 4516 2641
rect 4467 2601 4479 2635
rect 4513 2601 4516 2635
rect 4467 2595 4516 2601
rect 4510 2592 4516 2595
rect 4568 2592 4574 2644
rect 7270 2592 7276 2644
rect 7328 2641 7334 2644
rect 7328 2635 7377 2641
rect 7328 2601 7331 2635
rect 7365 2601 7377 2635
rect 7730 2632 7736 2644
rect 7691 2604 7736 2632
rect 7328 2595 7377 2601
rect 7328 2592 7334 2595
rect 7730 2592 7736 2604
rect 7788 2592 7794 2644
rect 8331 2635 8389 2641
rect 8331 2601 8343 2635
rect 8377 2632 8389 2635
rect 8650 2632 8656 2644
rect 8377 2604 8656 2632
rect 8377 2601 8389 2604
rect 8331 2595 8389 2601
rect 8650 2592 8656 2604
rect 8708 2592 8714 2644
rect 9619 2635 9677 2641
rect 9619 2601 9631 2635
rect 9665 2632 9677 2635
rect 10214 2632 10220 2644
rect 9665 2604 10220 2632
rect 9665 2601 9677 2604
rect 9619 2595 9677 2601
rect 10214 2592 10220 2604
rect 10272 2592 10278 2644
rect 11318 2632 11324 2644
rect 10508 2604 11324 2632
rect 1544 2499 1602 2505
rect 1544 2465 1556 2499
rect 1590 2496 1602 2499
rect 2556 2499 2614 2505
rect 1590 2468 2072 2496
rect 1590 2465 1602 2468
rect 1544 2459 1602 2465
rect 2044 2301 2072 2468
rect 2556 2465 2568 2499
rect 2602 2496 2614 2499
rect 3038 2496 3044 2508
rect 2602 2468 3044 2496
rect 2602 2465 2614 2468
rect 2556 2459 2614 2465
rect 3038 2456 3044 2468
rect 3096 2456 3102 2508
rect 4326 2456 4332 2508
rect 4384 2505 4390 2508
rect 4384 2499 4422 2505
rect 4410 2496 4422 2499
rect 4789 2499 4847 2505
rect 4789 2496 4801 2499
rect 4410 2468 4801 2496
rect 4410 2465 4422 2468
rect 4384 2459 4422 2465
rect 4789 2465 4801 2468
rect 4835 2465 4847 2499
rect 4789 2459 4847 2465
rect 7248 2499 7306 2505
rect 7248 2465 7260 2499
rect 7294 2496 7306 2499
rect 7748 2496 7776 2592
rect 9113 2567 9171 2573
rect 9113 2533 9125 2567
rect 9159 2564 9171 2567
rect 10508 2564 10536 2604
rect 9159 2536 10536 2564
rect 9159 2533 9171 2536
rect 9113 2527 9171 2533
rect 7294 2468 7776 2496
rect 8260 2499 8318 2505
rect 7294 2465 7306 2468
rect 7248 2459 7306 2465
rect 8260 2465 8272 2499
rect 8306 2496 8318 2499
rect 8742 2496 8748 2508
rect 8306 2468 8748 2496
rect 8306 2465 8318 2468
rect 8260 2459 8318 2465
rect 4384 2456 4390 2459
rect 8742 2456 8748 2468
rect 8800 2456 8806 2508
rect 10692 2505 10720 2604
rect 11318 2592 11324 2604
rect 11376 2592 11382 2644
rect 13253 2635 13311 2641
rect 13253 2601 13265 2635
rect 13299 2632 13311 2635
rect 13526 2632 13532 2644
rect 13299 2604 13532 2632
rect 13299 2601 13311 2604
rect 13253 2595 13311 2601
rect 13526 2592 13532 2604
rect 13584 2592 13590 2644
rect 14814 2632 14820 2644
rect 14775 2604 14820 2632
rect 14814 2592 14820 2604
rect 14872 2632 14878 2644
rect 16105 2635 16163 2641
rect 14872 2604 15136 2632
rect 14872 2592 14878 2604
rect 11965 2567 12023 2573
rect 11965 2533 11977 2567
rect 12011 2564 12023 2567
rect 12333 2567 12391 2573
rect 12333 2564 12345 2567
rect 12011 2536 12345 2564
rect 12011 2533 12023 2536
rect 11965 2527 12023 2533
rect 12333 2533 12345 2536
rect 12379 2564 12391 2567
rect 15001 2567 15059 2573
rect 15001 2564 15013 2567
rect 12379 2536 15013 2564
rect 12379 2533 12391 2536
rect 12333 2527 12391 2533
rect 15001 2533 15013 2536
rect 15047 2533 15059 2567
rect 15001 2527 15059 2533
rect 9548 2499 9606 2505
rect 9548 2465 9560 2499
rect 9594 2496 9606 2499
rect 10677 2499 10735 2505
rect 9594 2468 10076 2496
rect 9594 2465 9606 2468
rect 9548 2459 9606 2465
rect 5338 2428 5344 2440
rect 5299 2400 5344 2428
rect 5338 2388 5344 2400
rect 5396 2388 5402 2440
rect 2029 2295 2087 2301
rect 2029 2261 2041 2295
rect 2075 2292 2087 2295
rect 2118 2292 2124 2304
rect 2075 2264 2124 2292
rect 2075 2261 2087 2264
rect 2029 2255 2087 2261
rect 2118 2252 2124 2264
rect 2176 2252 2182 2304
rect 2627 2295 2685 2301
rect 2627 2261 2639 2295
rect 2673 2292 2685 2295
rect 2854 2292 2860 2304
rect 2673 2264 2860 2292
rect 2673 2261 2685 2264
rect 2627 2255 2685 2261
rect 2854 2252 2860 2264
rect 2912 2252 2918 2304
rect 3038 2292 3044 2304
rect 2999 2264 3044 2292
rect 3038 2252 3044 2264
rect 3096 2252 3102 2304
rect 8742 2292 8748 2304
rect 8703 2264 8748 2292
rect 8742 2252 8748 2264
rect 8800 2252 8806 2304
rect 10048 2301 10076 2468
rect 10677 2465 10689 2499
rect 10723 2465 10735 2499
rect 13802 2496 13808 2508
rect 13763 2468 13808 2496
rect 10677 2459 10735 2465
rect 13802 2456 13808 2468
rect 13860 2496 13866 2508
rect 15108 2505 15136 2604
rect 16105 2601 16117 2635
rect 16151 2632 16163 2635
rect 16286 2632 16292 2644
rect 16151 2604 16292 2632
rect 16151 2601 16163 2604
rect 16105 2595 16163 2601
rect 16286 2592 16292 2604
rect 16344 2592 16350 2644
rect 23373 2635 23431 2641
rect 23373 2601 23385 2635
rect 23419 2632 23431 2635
rect 23462 2632 23468 2644
rect 23419 2604 23468 2632
rect 23419 2601 23431 2604
rect 23373 2595 23431 2601
rect 23462 2592 23468 2604
rect 23520 2632 23526 2644
rect 23520 2604 23692 2632
rect 23520 2592 23526 2604
rect 18313 2567 18371 2573
rect 18313 2533 18325 2567
rect 18359 2564 18371 2567
rect 18589 2567 18647 2573
rect 18589 2564 18601 2567
rect 18359 2536 18601 2564
rect 18359 2533 18371 2536
rect 18313 2527 18371 2533
rect 18589 2533 18601 2536
rect 18635 2564 18647 2567
rect 18678 2564 18684 2576
rect 18635 2536 18684 2564
rect 18635 2533 18647 2536
rect 18589 2527 18647 2533
rect 18678 2524 18684 2536
rect 18736 2524 18742 2576
rect 19690 2524 19696 2576
rect 19748 2564 19754 2576
rect 20705 2567 20763 2573
rect 20705 2564 20717 2567
rect 19748 2536 20717 2564
rect 19748 2524 19754 2536
rect 20705 2533 20717 2536
rect 20751 2533 20763 2567
rect 20705 2527 20763 2533
rect 23002 2524 23008 2576
rect 23060 2564 23066 2576
rect 23557 2567 23615 2573
rect 23557 2564 23569 2567
rect 23060 2536 23569 2564
rect 23060 2524 23066 2536
rect 23557 2533 23569 2536
rect 23603 2533 23615 2567
rect 23557 2527 23615 2533
rect 14357 2499 14415 2505
rect 14357 2496 14369 2499
rect 13860 2468 14369 2496
rect 13860 2456 13866 2468
rect 14357 2465 14369 2468
rect 14403 2465 14415 2499
rect 14357 2459 14415 2465
rect 15093 2499 15151 2505
rect 15093 2465 15105 2499
rect 15139 2465 15151 2499
rect 16654 2496 16660 2508
rect 16615 2468 16660 2496
rect 15093 2459 15151 2465
rect 16654 2456 16660 2468
rect 16712 2496 16718 2508
rect 17209 2499 17267 2505
rect 17209 2496 17221 2499
rect 16712 2468 17221 2496
rect 16712 2456 16718 2468
rect 17209 2465 17221 2468
rect 17255 2465 17267 2499
rect 17209 2459 17267 2465
rect 20334 2456 20340 2508
rect 20392 2496 20398 2508
rect 20521 2499 20579 2505
rect 20521 2496 20533 2499
rect 20392 2468 20533 2496
rect 20392 2456 20398 2468
rect 20521 2465 20533 2468
rect 20567 2496 20579 2499
rect 20797 2499 20855 2505
rect 20797 2496 20809 2499
rect 20567 2468 20809 2496
rect 20567 2465 20579 2468
rect 20521 2459 20579 2465
rect 20797 2465 20809 2468
rect 20843 2465 20855 2499
rect 22266 2496 22272 2508
rect 22227 2468 22272 2496
rect 20797 2459 20855 2465
rect 22266 2456 22272 2468
rect 22324 2496 22330 2508
rect 23664 2505 23692 2604
rect 25210 2592 25216 2644
rect 25268 2641 25274 2644
rect 25268 2635 25317 2641
rect 25268 2601 25271 2635
rect 25305 2601 25317 2635
rect 25268 2595 25317 2601
rect 25268 2592 25274 2595
rect 22821 2499 22879 2505
rect 22821 2496 22833 2499
rect 22324 2468 22833 2496
rect 22324 2456 22330 2468
rect 22821 2465 22833 2468
rect 22867 2465 22879 2499
rect 22821 2459 22879 2465
rect 23649 2499 23707 2505
rect 23649 2465 23661 2499
rect 23695 2465 23707 2499
rect 23649 2459 23707 2465
rect 24382 2456 24388 2508
rect 24440 2496 24446 2508
rect 25156 2499 25214 2505
rect 25156 2496 25168 2499
rect 24440 2468 25168 2496
rect 24440 2456 24446 2468
rect 25156 2465 25168 2468
rect 25202 2496 25214 2499
rect 25581 2499 25639 2505
rect 25581 2496 25593 2499
rect 25202 2468 25593 2496
rect 25202 2465 25214 2468
rect 25156 2459 25214 2465
rect 25581 2465 25593 2468
rect 25627 2465 25639 2499
rect 25581 2459 25639 2465
rect 10401 2431 10459 2437
rect 10401 2397 10413 2431
rect 10447 2428 10459 2431
rect 10490 2428 10496 2440
rect 10447 2400 10496 2428
rect 10447 2397 10459 2400
rect 10401 2391 10459 2397
rect 10490 2388 10496 2400
rect 10548 2388 10554 2440
rect 11502 2428 11508 2440
rect 11463 2400 11508 2428
rect 11502 2388 11508 2400
rect 11560 2428 11566 2440
rect 12241 2431 12299 2437
rect 12241 2428 12253 2431
rect 11560 2400 12253 2428
rect 11560 2388 11566 2400
rect 12241 2397 12253 2400
rect 12287 2397 12299 2431
rect 12241 2391 12299 2397
rect 12330 2388 12336 2440
rect 12388 2428 12394 2440
rect 12517 2431 12575 2437
rect 12517 2428 12529 2431
rect 12388 2400 12529 2428
rect 12388 2388 12394 2400
rect 12517 2397 12529 2400
rect 12563 2397 12575 2431
rect 18497 2431 18555 2437
rect 18497 2428 18509 2431
rect 12517 2391 12575 2397
rect 17592 2400 18509 2428
rect 16841 2363 16899 2369
rect 16841 2329 16853 2363
rect 16887 2360 16899 2363
rect 17482 2360 17488 2372
rect 16887 2332 17488 2360
rect 16887 2329 16899 2332
rect 16841 2323 16899 2329
rect 17482 2320 17488 2332
rect 17540 2320 17546 2372
rect 17592 2304 17620 2400
rect 18497 2397 18509 2400
rect 18543 2397 18555 2431
rect 18497 2391 18555 2397
rect 19046 2360 19052 2372
rect 19007 2332 19052 2360
rect 19046 2320 19052 2332
rect 19104 2320 19110 2372
rect 10033 2295 10091 2301
rect 10033 2261 10045 2295
rect 10079 2292 10091 2295
rect 10306 2292 10312 2304
rect 10079 2264 10312 2292
rect 10079 2261 10091 2264
rect 10033 2255 10091 2261
rect 10306 2252 10312 2264
rect 10364 2252 10370 2304
rect 13986 2292 13992 2304
rect 13947 2264 13992 2292
rect 13986 2252 13992 2264
rect 14044 2252 14050 2304
rect 17574 2292 17580 2304
rect 17535 2264 17580 2292
rect 17574 2252 17580 2264
rect 17632 2252 17638 2304
rect 18954 2252 18960 2304
rect 19012 2292 19018 2304
rect 19414 2292 19420 2304
rect 19012 2264 19420 2292
rect 19012 2252 19018 2264
rect 19414 2252 19420 2264
rect 19472 2252 19478 2304
rect 20058 2292 20064 2304
rect 20019 2264 20064 2292
rect 20058 2252 20064 2264
rect 20116 2252 20122 2304
rect 22450 2292 22456 2304
rect 22411 2264 22456 2292
rect 22450 2252 22456 2264
rect 22508 2252 22514 2304
rect 632 2202 26392 2224
rect 632 2150 5176 2202
rect 5228 2150 5240 2202
rect 5292 2150 5304 2202
rect 5356 2150 5368 2202
rect 5420 2150 14510 2202
rect 14562 2150 14574 2202
rect 14626 2150 14638 2202
rect 14690 2150 14702 2202
rect 14754 2150 23843 2202
rect 23895 2150 23907 2202
rect 23959 2150 23971 2202
rect 24023 2150 24035 2202
rect 24087 2150 26392 2202
rect 632 2128 26392 2150
<< via1 >>
rect 3688 27412 3740 27464
rect 4792 27412 4844 27464
rect 9843 25542 9895 25594
rect 9907 25542 9959 25594
rect 9971 25542 10023 25594
rect 10035 25542 10087 25594
rect 19176 25542 19228 25594
rect 19240 25542 19292 25594
rect 19304 25542 19356 25594
rect 19368 25542 19420 25594
rect 5176 24998 5228 25050
rect 5240 24998 5292 25050
rect 5304 24998 5356 25050
rect 5368 24998 5420 25050
rect 14510 24998 14562 25050
rect 14574 24998 14626 25050
rect 14638 24998 14690 25050
rect 14702 24998 14754 25050
rect 23843 24998 23895 25050
rect 23907 24998 23959 25050
rect 23971 24998 24023 25050
rect 24035 24998 24087 25050
rect 9843 24454 9895 24506
rect 9907 24454 9959 24506
rect 9971 24454 10023 24506
rect 10035 24454 10087 24506
rect 19176 24454 19228 24506
rect 19240 24454 19292 24506
rect 19304 24454 19356 24506
rect 19368 24454 19420 24506
rect 5176 23910 5228 23962
rect 5240 23910 5292 23962
rect 5304 23910 5356 23962
rect 5368 23910 5420 23962
rect 14510 23910 14562 23962
rect 14574 23910 14626 23962
rect 14638 23910 14690 23962
rect 14702 23910 14754 23962
rect 23843 23910 23895 23962
rect 23907 23910 23959 23962
rect 23971 23910 24023 23962
rect 24035 23910 24087 23962
rect 24296 23808 24348 23860
rect 22916 23740 22968 23792
rect 24296 23604 24348 23656
rect 20340 23468 20392 23520
rect 23008 23468 23060 23520
rect 9843 23366 9895 23418
rect 9907 23366 9959 23418
rect 9971 23366 10023 23418
rect 10035 23366 10087 23418
rect 19176 23366 19228 23418
rect 19240 23366 19292 23418
rect 19304 23366 19356 23418
rect 19368 23366 19420 23418
rect 5176 22822 5228 22874
rect 5240 22822 5292 22874
rect 5304 22822 5356 22874
rect 5368 22822 5420 22874
rect 14510 22822 14562 22874
rect 14574 22822 14626 22874
rect 14638 22822 14690 22874
rect 14702 22822 14754 22874
rect 23843 22822 23895 22874
rect 23907 22822 23959 22874
rect 23971 22822 24023 22874
rect 24035 22822 24087 22874
rect 9843 22278 9895 22330
rect 9907 22278 9959 22330
rect 9971 22278 10023 22330
rect 10035 22278 10087 22330
rect 19176 22278 19228 22330
rect 19240 22278 19292 22330
rect 19304 22278 19356 22330
rect 19368 22278 19420 22330
rect 5176 21734 5228 21786
rect 5240 21734 5292 21786
rect 5304 21734 5356 21786
rect 5368 21734 5420 21786
rect 14510 21734 14562 21786
rect 14574 21734 14626 21786
rect 14638 21734 14690 21786
rect 14702 21734 14754 21786
rect 23843 21734 23895 21786
rect 23907 21734 23959 21786
rect 23971 21734 24023 21786
rect 24035 21734 24087 21786
rect 24296 21632 24348 21684
rect 24296 21428 24348 21480
rect 22364 21292 22416 21344
rect 9843 21190 9895 21242
rect 9907 21190 9959 21242
rect 9971 21190 10023 21242
rect 10035 21190 10087 21242
rect 19176 21190 19228 21242
rect 19240 21190 19292 21242
rect 19304 21190 19356 21242
rect 19368 21190 19420 21242
rect 24204 20995 24256 21004
rect 24204 20961 24222 20995
rect 24222 20961 24256 20995
rect 24204 20952 24256 20961
rect 23284 20748 23336 20800
rect 5176 20646 5228 20698
rect 5240 20646 5292 20698
rect 5304 20646 5356 20698
rect 5368 20646 5420 20698
rect 14510 20646 14562 20698
rect 14574 20646 14626 20698
rect 14638 20646 14690 20698
rect 14702 20646 14754 20698
rect 23843 20646 23895 20698
rect 23907 20646 23959 20698
rect 23971 20646 24023 20698
rect 24035 20646 24087 20698
rect 24204 20587 24256 20596
rect 24204 20553 24213 20587
rect 24213 20553 24247 20587
rect 24247 20553 24256 20587
rect 24204 20544 24256 20553
rect 9843 20102 9895 20154
rect 9907 20102 9959 20154
rect 9971 20102 10023 20154
rect 10035 20102 10087 20154
rect 19176 20102 19228 20154
rect 19240 20102 19292 20154
rect 19304 20102 19356 20154
rect 19368 20102 19420 20154
rect 25032 19864 25084 19916
rect 23008 19660 23060 19712
rect 5176 19558 5228 19610
rect 5240 19558 5292 19610
rect 5304 19558 5356 19610
rect 5368 19558 5420 19610
rect 14510 19558 14562 19610
rect 14574 19558 14626 19610
rect 14638 19558 14690 19610
rect 14702 19558 14754 19610
rect 23843 19558 23895 19610
rect 23907 19558 23959 19610
rect 23971 19558 24023 19610
rect 24035 19558 24087 19610
rect 25032 19295 25084 19304
rect 23008 19184 23060 19236
rect 25032 19261 25041 19295
rect 25041 19261 25075 19295
rect 25075 19261 25084 19295
rect 25032 19252 25084 19261
rect 25492 19116 25544 19168
rect 9843 19014 9895 19066
rect 9907 19014 9959 19066
rect 9971 19014 10023 19066
rect 10035 19014 10087 19066
rect 19176 19014 19228 19066
rect 19240 19014 19292 19066
rect 19304 19014 19356 19066
rect 19368 19014 19420 19066
rect 20524 18819 20576 18828
rect 20524 18785 20542 18819
rect 20542 18785 20576 18819
rect 20524 18776 20576 18785
rect 23468 18776 23520 18828
rect 25032 18776 25084 18828
rect 23008 18640 23060 18692
rect 20524 18572 20576 18624
rect 23100 18572 23152 18624
rect 5176 18470 5228 18522
rect 5240 18470 5292 18522
rect 5304 18470 5356 18522
rect 5368 18470 5420 18522
rect 14510 18470 14562 18522
rect 14574 18470 14626 18522
rect 14638 18470 14690 18522
rect 14702 18470 14754 18522
rect 23843 18470 23895 18522
rect 23907 18470 23959 18522
rect 23971 18470 24023 18522
rect 24035 18470 24087 18522
rect 20432 18411 20484 18420
rect 20432 18377 20441 18411
rect 20441 18377 20475 18411
rect 20475 18377 20484 18411
rect 20432 18368 20484 18377
rect 23468 18275 23520 18284
rect 23468 18241 23477 18275
rect 23477 18241 23511 18275
rect 23511 18241 23520 18275
rect 23468 18232 23520 18241
rect 24296 18232 24348 18284
rect 23652 18096 23704 18148
rect 25124 18207 25176 18216
rect 25124 18173 25168 18207
rect 25168 18173 25176 18207
rect 25124 18164 25176 18173
rect 22088 18028 22140 18080
rect 22640 18071 22692 18080
rect 22640 18037 22649 18071
rect 22649 18037 22683 18071
rect 22683 18037 22692 18071
rect 22640 18028 22692 18037
rect 23468 18028 23520 18080
rect 25032 18071 25084 18080
rect 25032 18037 25041 18071
rect 25041 18037 25075 18071
rect 25075 18037 25084 18071
rect 25032 18028 25084 18037
rect 25216 18028 25268 18080
rect 9843 17926 9895 17978
rect 9907 17926 9959 17978
rect 9971 17926 10023 17978
rect 10035 17926 10087 17978
rect 19176 17926 19228 17978
rect 19240 17926 19292 17978
rect 19304 17926 19356 17978
rect 19368 17926 19420 17978
rect 21536 17867 21588 17876
rect 21536 17833 21545 17867
rect 21545 17833 21579 17867
rect 21579 17833 21588 17867
rect 21536 17824 21588 17833
rect 20432 17688 20484 17740
rect 22732 17688 22784 17740
rect 24204 17731 24256 17740
rect 24204 17697 24222 17731
rect 24222 17697 24256 17731
rect 24204 17688 24256 17697
rect 20708 17527 20760 17536
rect 20708 17493 20717 17527
rect 20717 17493 20751 17527
rect 20751 17493 20760 17527
rect 20708 17484 20760 17493
rect 22180 17484 22232 17536
rect 23008 17484 23060 17536
rect 5176 17382 5228 17434
rect 5240 17382 5292 17434
rect 5304 17382 5356 17434
rect 5368 17382 5420 17434
rect 14510 17382 14562 17434
rect 14574 17382 14626 17434
rect 14638 17382 14690 17434
rect 14702 17382 14754 17434
rect 23843 17382 23895 17434
rect 23907 17382 23959 17434
rect 23971 17382 24023 17434
rect 24035 17382 24087 17434
rect 24204 17323 24256 17332
rect 24204 17289 24213 17323
rect 24213 17289 24247 17323
rect 24247 17289 24256 17323
rect 24204 17280 24256 17289
rect 21536 17212 21588 17264
rect 21628 17187 21680 17196
rect 21628 17153 21637 17187
rect 21637 17153 21671 17187
rect 21671 17153 21680 17187
rect 21628 17144 21680 17153
rect 16200 17076 16252 17128
rect 19972 17076 20024 17128
rect 16568 17051 16620 17060
rect 16568 17017 16577 17051
rect 16577 17017 16611 17051
rect 16611 17017 16620 17051
rect 16568 17008 16620 17017
rect 20156 16940 20208 16992
rect 20432 16940 20484 16992
rect 24388 17008 24440 17060
rect 22732 16940 22784 16992
rect 23376 16940 23428 16992
rect 24296 16940 24348 16992
rect 9843 16838 9895 16890
rect 9907 16838 9959 16890
rect 9971 16838 10023 16890
rect 10035 16838 10087 16890
rect 19176 16838 19228 16890
rect 19240 16838 19292 16890
rect 19304 16838 19356 16890
rect 19368 16838 19420 16890
rect 15648 16736 15700 16788
rect 16016 16779 16068 16788
rect 16016 16745 16025 16779
rect 16025 16745 16059 16779
rect 16059 16745 16068 16779
rect 16016 16736 16068 16745
rect 18684 16736 18736 16788
rect 16568 16668 16620 16720
rect 20708 16668 20760 16720
rect 24388 16668 24440 16720
rect 14912 16643 14964 16652
rect 14912 16609 14921 16643
rect 14921 16609 14955 16643
rect 14955 16609 14964 16643
rect 14912 16600 14964 16609
rect 15740 16600 15792 16652
rect 18224 16643 18276 16652
rect 18224 16609 18233 16643
rect 18233 16609 18267 16643
rect 18267 16609 18276 16643
rect 18224 16600 18276 16609
rect 22548 16643 22600 16652
rect 22548 16609 22557 16643
rect 22557 16609 22591 16643
rect 22591 16609 22600 16643
rect 22548 16600 22600 16609
rect 23744 16643 23796 16652
rect 23744 16609 23788 16643
rect 23788 16609 23796 16643
rect 23744 16600 23796 16609
rect 24204 16600 24256 16652
rect 25400 16600 25452 16652
rect 16660 16532 16712 16584
rect 16844 16575 16896 16584
rect 16844 16541 16853 16575
rect 16853 16541 16887 16575
rect 16887 16541 16896 16575
rect 16844 16532 16896 16541
rect 20248 16532 20300 16584
rect 21444 16532 21496 16584
rect 21628 16532 21680 16584
rect 19512 16439 19564 16448
rect 19512 16405 19521 16439
rect 19521 16405 19555 16439
rect 19555 16405 19564 16439
rect 19512 16396 19564 16405
rect 22456 16439 22508 16448
rect 22456 16405 22465 16439
rect 22465 16405 22499 16439
rect 22499 16405 22508 16439
rect 22456 16396 22508 16405
rect 5176 16294 5228 16346
rect 5240 16294 5292 16346
rect 5304 16294 5356 16346
rect 5368 16294 5420 16346
rect 14510 16294 14562 16346
rect 14574 16294 14626 16346
rect 14638 16294 14690 16346
rect 14702 16294 14754 16346
rect 23843 16294 23895 16346
rect 23907 16294 23959 16346
rect 23971 16294 24023 16346
rect 24035 16294 24087 16346
rect 16568 16235 16620 16244
rect 16568 16201 16577 16235
rect 16577 16201 16611 16235
rect 16611 16201 16620 16235
rect 16568 16192 16620 16201
rect 20432 16235 20484 16244
rect 20432 16201 20441 16235
rect 20441 16201 20475 16235
rect 20475 16201 20484 16235
rect 20432 16192 20484 16201
rect 20708 16235 20760 16244
rect 20708 16201 20717 16235
rect 20717 16201 20751 16235
rect 20751 16201 20760 16235
rect 20708 16192 20760 16201
rect 21720 16192 21772 16244
rect 22548 16235 22600 16244
rect 22548 16201 22557 16235
rect 22557 16201 22591 16235
rect 22591 16201 22600 16235
rect 22548 16192 22600 16201
rect 16660 16056 16712 16108
rect 21444 16056 21496 16108
rect 17396 16031 17448 16040
rect 17396 15997 17405 16031
rect 17405 15997 17439 16031
rect 17439 15997 17448 16031
rect 17396 15988 17448 15997
rect 19512 16031 19564 16040
rect 19512 15997 19521 16031
rect 19521 15997 19555 16031
rect 19555 15997 19564 16031
rect 19512 15988 19564 15997
rect 23284 16031 23336 16040
rect 23284 15997 23293 16031
rect 23293 15997 23327 16031
rect 23327 15997 23336 16031
rect 23284 15988 23336 15997
rect 15648 15963 15700 15972
rect 15648 15929 15657 15963
rect 15657 15929 15691 15963
rect 15691 15929 15700 15963
rect 15648 15920 15700 15929
rect 15740 15963 15792 15972
rect 15740 15929 15749 15963
rect 15749 15929 15783 15963
rect 15783 15929 15792 15963
rect 15740 15920 15792 15929
rect 17120 15920 17172 15972
rect 16752 15852 16804 15904
rect 20892 15920 20944 15972
rect 21720 15963 21772 15972
rect 21720 15929 21729 15963
rect 21729 15929 21763 15963
rect 21763 15929 21772 15963
rect 21720 15920 21772 15929
rect 22548 15920 22600 15972
rect 23744 15920 23796 15972
rect 18224 15852 18276 15904
rect 18776 15852 18828 15904
rect 23560 15852 23612 15904
rect 24756 15895 24808 15904
rect 24756 15861 24765 15895
rect 24765 15861 24799 15895
rect 24799 15861 24808 15895
rect 24756 15852 24808 15861
rect 25400 15852 25452 15904
rect 9843 15750 9895 15802
rect 9907 15750 9959 15802
rect 9971 15750 10023 15802
rect 10035 15750 10087 15802
rect 19176 15750 19228 15802
rect 19240 15750 19292 15802
rect 19304 15750 19356 15802
rect 19368 15750 19420 15802
rect 16200 15691 16252 15700
rect 16200 15657 16209 15691
rect 16209 15657 16243 15691
rect 16243 15657 16252 15691
rect 16200 15648 16252 15657
rect 17028 15648 17080 15700
rect 15924 15580 15976 15632
rect 21444 15648 21496 15700
rect 20892 15580 20944 15632
rect 22272 15623 22324 15632
rect 22272 15589 22281 15623
rect 22281 15589 22315 15623
rect 22315 15589 22324 15623
rect 22272 15580 22324 15589
rect 22456 15580 22508 15632
rect 12888 15555 12940 15564
rect 12888 15521 12897 15555
rect 12897 15521 12931 15555
rect 12931 15521 12940 15555
rect 12888 15512 12940 15521
rect 13072 15555 13124 15564
rect 13072 15521 13078 15555
rect 13078 15521 13124 15555
rect 13072 15512 13124 15521
rect 19052 15555 19104 15564
rect 19052 15521 19061 15555
rect 19061 15521 19095 15555
rect 19095 15521 19104 15555
rect 19052 15512 19104 15521
rect 19144 15512 19196 15564
rect 21720 15512 21772 15564
rect 24572 15512 24624 15564
rect 12612 15444 12664 15496
rect 13624 15444 13676 15496
rect 14820 15444 14872 15496
rect 15372 15444 15424 15496
rect 16016 15444 16068 15496
rect 17120 15487 17172 15496
rect 17120 15453 17129 15487
rect 17129 15453 17163 15487
rect 17163 15453 17172 15487
rect 17120 15444 17172 15453
rect 11784 15376 11836 15428
rect 12152 15376 12204 15428
rect 16844 15376 16896 15428
rect 20064 15444 20116 15496
rect 22548 15487 22600 15496
rect 22548 15453 22557 15487
rect 22557 15453 22591 15487
rect 22591 15453 22600 15487
rect 22548 15444 22600 15453
rect 24848 15444 24900 15496
rect 20248 15419 20300 15428
rect 20248 15385 20257 15419
rect 20257 15385 20291 15419
rect 20291 15385 20300 15419
rect 20248 15376 20300 15385
rect 13164 15351 13216 15360
rect 13164 15317 13173 15351
rect 13173 15317 13207 15351
rect 13207 15317 13216 15351
rect 13164 15308 13216 15317
rect 13532 15351 13584 15360
rect 13532 15317 13541 15351
rect 13541 15317 13575 15351
rect 13575 15317 13584 15351
rect 13532 15308 13584 15317
rect 13716 15308 13768 15360
rect 15004 15351 15056 15360
rect 15004 15317 15013 15351
rect 15013 15317 15047 15351
rect 15047 15317 15056 15351
rect 15004 15308 15056 15317
rect 5176 15206 5228 15258
rect 5240 15206 5292 15258
rect 5304 15206 5356 15258
rect 5368 15206 5420 15258
rect 14510 15206 14562 15258
rect 14574 15206 14626 15258
rect 14638 15206 14690 15258
rect 14702 15206 14754 15258
rect 23843 15206 23895 15258
rect 23907 15206 23959 15258
rect 23971 15206 24023 15258
rect 24035 15206 24087 15258
rect 12520 15104 12572 15156
rect 12888 15104 12940 15156
rect 13164 15104 13216 15156
rect 15740 15104 15792 15156
rect 16108 15104 16160 15156
rect 17028 15147 17080 15156
rect 17028 15113 17037 15147
rect 17037 15113 17071 15147
rect 17071 15113 17080 15147
rect 17028 15104 17080 15113
rect 20064 15147 20116 15156
rect 20064 15113 20073 15147
rect 20073 15113 20107 15147
rect 20107 15113 20116 15147
rect 20064 15104 20116 15113
rect 20892 15104 20944 15156
rect 22456 15104 22508 15156
rect 24940 15104 24992 15156
rect 12612 15079 12664 15088
rect 12612 15045 12621 15079
rect 12621 15045 12655 15079
rect 12655 15045 12664 15079
rect 12612 15036 12664 15045
rect 15004 14968 15056 15020
rect 19512 14968 19564 15020
rect 20340 14968 20392 15020
rect 22272 14968 22324 15020
rect 13440 14943 13492 14952
rect 13440 14909 13449 14943
rect 13449 14909 13483 14943
rect 13483 14909 13492 14943
rect 13440 14900 13492 14909
rect 13716 14943 13768 14952
rect 13716 14909 13725 14943
rect 13725 14909 13759 14943
rect 13759 14909 13768 14943
rect 13716 14900 13768 14909
rect 18592 14943 18644 14952
rect 18592 14909 18601 14943
rect 18601 14909 18635 14943
rect 18635 14909 18644 14943
rect 18592 14900 18644 14909
rect 19144 14900 19196 14952
rect 23008 14943 23060 14952
rect 23008 14909 23017 14943
rect 23017 14909 23051 14943
rect 23051 14909 23060 14943
rect 23008 14900 23060 14909
rect 24940 14900 24992 14952
rect 15924 14807 15976 14816
rect 15924 14773 15933 14807
rect 15933 14773 15967 14807
rect 15967 14773 15976 14807
rect 15924 14764 15976 14773
rect 16936 14764 16988 14816
rect 17948 14807 18000 14816
rect 17948 14773 17957 14807
rect 17957 14773 17991 14807
rect 17991 14773 18000 14807
rect 19972 14832 20024 14884
rect 20248 14832 20300 14884
rect 17948 14764 18000 14773
rect 19052 14764 19104 14816
rect 21628 14832 21680 14884
rect 23192 14875 23244 14884
rect 23192 14841 23201 14875
rect 23201 14841 23235 14875
rect 23235 14841 23244 14875
rect 23192 14832 23244 14841
rect 24572 14832 24624 14884
rect 24480 14764 24532 14816
rect 9843 14662 9895 14714
rect 9907 14662 9959 14714
rect 9971 14662 10023 14714
rect 10035 14662 10087 14714
rect 19176 14662 19228 14714
rect 19240 14662 19292 14714
rect 19304 14662 19356 14714
rect 19368 14662 19420 14714
rect 13072 14560 13124 14612
rect 16016 14560 16068 14612
rect 17856 14603 17908 14612
rect 17856 14569 17865 14603
rect 17865 14569 17899 14603
rect 17899 14569 17908 14603
rect 17856 14560 17908 14569
rect 18592 14603 18644 14612
rect 18592 14569 18601 14603
rect 18601 14569 18635 14603
rect 18635 14569 18644 14603
rect 18592 14560 18644 14569
rect 20340 14560 20392 14612
rect 21444 14560 21496 14612
rect 23008 14560 23060 14612
rect 9576 14492 9628 14544
rect 9668 14467 9720 14476
rect 9668 14433 9677 14467
rect 9677 14433 9711 14467
rect 9711 14433 9720 14467
rect 9668 14424 9720 14433
rect 14912 14492 14964 14544
rect 17120 14492 17172 14544
rect 20616 14492 20668 14544
rect 20892 14492 20944 14544
rect 21628 14535 21680 14544
rect 21628 14501 21637 14535
rect 21637 14501 21671 14535
rect 21671 14501 21680 14535
rect 21628 14492 21680 14501
rect 22640 14492 22692 14544
rect 23192 14492 23244 14544
rect 11876 14424 11928 14476
rect 13440 14467 13492 14476
rect 13440 14433 13449 14467
rect 13449 14433 13483 14467
rect 13483 14433 13492 14467
rect 13440 14424 13492 14433
rect 13808 14424 13860 14476
rect 16660 14467 16712 14476
rect 16660 14433 16669 14467
rect 16669 14433 16703 14467
rect 16703 14433 16712 14467
rect 16660 14424 16712 14433
rect 16844 14467 16896 14476
rect 16844 14433 16853 14467
rect 16853 14433 16887 14467
rect 16887 14433 16896 14467
rect 16844 14424 16896 14433
rect 19052 14467 19104 14476
rect 19052 14433 19061 14467
rect 19061 14433 19095 14467
rect 19095 14433 19104 14467
rect 19052 14424 19104 14433
rect 19696 14424 19748 14476
rect 23652 14424 23704 14476
rect 14360 14356 14412 14408
rect 14912 14399 14964 14408
rect 14912 14365 14921 14399
rect 14921 14365 14955 14399
rect 14955 14365 14964 14399
rect 14912 14356 14964 14365
rect 20892 14356 20944 14408
rect 22272 14399 22324 14408
rect 22272 14365 22281 14399
rect 22281 14365 22315 14399
rect 22315 14365 22324 14399
rect 22272 14356 22324 14365
rect 22916 14399 22968 14408
rect 22916 14365 22925 14399
rect 22925 14365 22959 14399
rect 22959 14365 22968 14399
rect 22916 14356 22968 14365
rect 23008 14356 23060 14408
rect 9300 14220 9352 14272
rect 12336 14220 12388 14272
rect 19788 14263 19840 14272
rect 19788 14229 19797 14263
rect 19797 14229 19831 14263
rect 19831 14229 19840 14263
rect 19788 14220 19840 14229
rect 23192 14263 23244 14272
rect 23192 14229 23201 14263
rect 23201 14229 23235 14263
rect 23235 14229 23244 14263
rect 23192 14220 23244 14229
rect 5176 14118 5228 14170
rect 5240 14118 5292 14170
rect 5304 14118 5356 14170
rect 5368 14118 5420 14170
rect 14510 14118 14562 14170
rect 14574 14118 14626 14170
rect 14638 14118 14690 14170
rect 14702 14118 14754 14170
rect 23843 14118 23895 14170
rect 23907 14118 23959 14170
rect 23971 14118 24023 14170
rect 24035 14118 24087 14170
rect 8932 14059 8984 14068
rect 8932 14025 8941 14059
rect 8941 14025 8975 14059
rect 8975 14025 8984 14059
rect 8932 14016 8984 14025
rect 9576 14016 9628 14068
rect 13716 14016 13768 14068
rect 11784 13948 11836 14000
rect 9668 13880 9720 13932
rect 8932 13812 8984 13864
rect 9392 13812 9444 13864
rect 10588 13812 10640 13864
rect 13808 13923 13860 13932
rect 13808 13889 13817 13923
rect 13817 13889 13851 13923
rect 13851 13889 13860 13923
rect 13808 13880 13860 13889
rect 15004 14016 15056 14068
rect 16384 14059 16436 14068
rect 16384 14025 16393 14059
rect 16393 14025 16427 14059
rect 16427 14025 16436 14059
rect 16384 14016 16436 14025
rect 16844 14016 16896 14068
rect 17396 14059 17448 14068
rect 17396 14025 17405 14059
rect 17405 14025 17439 14059
rect 17439 14025 17448 14059
rect 17396 14016 17448 14025
rect 14820 13948 14872 14000
rect 16660 13948 16712 14000
rect 19052 14016 19104 14068
rect 20248 14059 20300 14068
rect 20248 14025 20257 14059
rect 20257 14025 20291 14059
rect 20291 14025 20300 14059
rect 20248 14016 20300 14025
rect 20616 14059 20668 14068
rect 20616 14025 20625 14059
rect 20625 14025 20659 14059
rect 20659 14025 20668 14059
rect 20616 14016 20668 14025
rect 20892 14059 20944 14068
rect 20892 14025 20901 14059
rect 20901 14025 20935 14059
rect 20935 14025 20944 14059
rect 20892 14016 20944 14025
rect 21444 14059 21496 14068
rect 21444 14025 21453 14059
rect 21453 14025 21487 14059
rect 21487 14025 21496 14059
rect 21444 14016 21496 14025
rect 22640 14059 22692 14068
rect 22640 14025 22649 14059
rect 22649 14025 22683 14059
rect 22683 14025 22692 14059
rect 22640 14016 22692 14025
rect 22916 14016 22968 14068
rect 23652 14016 23704 14068
rect 14268 13880 14320 13932
rect 17948 13923 18000 13932
rect 12520 13855 12572 13864
rect 12520 13821 12529 13855
rect 12529 13821 12563 13855
rect 12563 13821 12572 13855
rect 12520 13812 12572 13821
rect 13072 13855 13124 13864
rect 13072 13821 13081 13855
rect 13081 13821 13115 13855
rect 13115 13821 13124 13855
rect 13072 13812 13124 13821
rect 13440 13855 13492 13864
rect 13440 13821 13449 13855
rect 13449 13821 13483 13855
rect 13483 13821 13492 13855
rect 13440 13812 13492 13821
rect 14820 13855 14872 13864
rect 14820 13821 14829 13855
rect 14829 13821 14863 13855
rect 14863 13821 14872 13855
rect 14820 13812 14872 13821
rect 17948 13889 17957 13923
rect 17957 13889 17991 13923
rect 17991 13889 18000 13923
rect 17948 13880 18000 13889
rect 19788 13880 19840 13932
rect 11416 13744 11468 13796
rect 15372 13787 15424 13796
rect 15372 13753 15381 13787
rect 15381 13753 15415 13787
rect 15415 13753 15424 13787
rect 15372 13744 15424 13753
rect 17672 13787 17724 13796
rect 17672 13753 17681 13787
rect 17681 13753 17715 13787
rect 17715 13753 17724 13787
rect 17672 13744 17724 13753
rect 25308 13948 25360 14000
rect 21168 13880 21220 13932
rect 21628 13923 21680 13932
rect 21628 13889 21637 13923
rect 21637 13889 21671 13923
rect 21671 13889 21680 13923
rect 21628 13880 21680 13889
rect 21444 13812 21496 13864
rect 23008 13855 23060 13864
rect 23008 13821 23017 13855
rect 23017 13821 23051 13855
rect 23051 13821 23060 13855
rect 23008 13812 23060 13821
rect 23284 13812 23336 13864
rect 24020 13812 24072 13864
rect 24388 13812 24440 13864
rect 10680 13676 10732 13728
rect 11876 13676 11928 13728
rect 16476 13719 16528 13728
rect 16476 13685 16485 13719
rect 16485 13685 16519 13719
rect 16519 13685 16528 13719
rect 16476 13676 16528 13685
rect 17396 13676 17448 13728
rect 23192 13676 23244 13728
rect 9843 13574 9895 13626
rect 9907 13574 9959 13626
rect 9971 13574 10023 13626
rect 10035 13574 10087 13626
rect 19176 13574 19228 13626
rect 19240 13574 19292 13626
rect 19304 13574 19356 13626
rect 19368 13574 19420 13626
rect 12520 13472 12572 13524
rect 14912 13472 14964 13524
rect 15096 13472 15148 13524
rect 16016 13472 16068 13524
rect 17304 13472 17356 13524
rect 15924 13447 15976 13456
rect 15924 13413 15927 13447
rect 15927 13413 15961 13447
rect 15961 13413 15976 13447
rect 15924 13404 15976 13413
rect 16292 13404 16344 13456
rect 17028 13404 17080 13456
rect 17948 13472 18000 13524
rect 18868 13472 18920 13524
rect 22272 13515 22324 13524
rect 22272 13481 22281 13515
rect 22281 13481 22315 13515
rect 22315 13481 22324 13515
rect 22272 13472 22324 13481
rect 23284 13472 23336 13524
rect 24296 13472 24348 13524
rect 17580 13404 17632 13456
rect 9392 13379 9444 13388
rect 9392 13345 9401 13379
rect 9401 13345 9435 13379
rect 9435 13345 9444 13379
rect 9392 13336 9444 13345
rect 9576 13336 9628 13388
rect 11876 13379 11928 13388
rect 11876 13345 11885 13379
rect 11885 13345 11919 13379
rect 11919 13345 11928 13379
rect 11876 13336 11928 13345
rect 13072 13379 13124 13388
rect 13072 13345 13081 13379
rect 13081 13345 13115 13379
rect 13115 13345 13124 13379
rect 13072 13336 13124 13345
rect 14360 13336 14412 13388
rect 16108 13336 16160 13388
rect 19604 13404 19656 13456
rect 20156 13404 20208 13456
rect 21168 13447 21220 13456
rect 21168 13413 21177 13447
rect 21177 13413 21211 13447
rect 21211 13413 21220 13447
rect 21168 13404 21220 13413
rect 22456 13404 22508 13456
rect 22916 13404 22968 13456
rect 18960 13336 19012 13388
rect 24204 13379 24256 13388
rect 24204 13345 24213 13379
rect 24213 13345 24247 13379
rect 24247 13345 24256 13379
rect 24204 13336 24256 13345
rect 11784 13268 11836 13320
rect 14084 13268 14136 13320
rect 20340 13268 20392 13320
rect 22548 13268 22600 13320
rect 23100 13311 23152 13320
rect 23100 13277 23109 13311
rect 23109 13277 23143 13311
rect 23143 13277 23152 13311
rect 23100 13268 23152 13277
rect 23744 13268 23796 13320
rect 17948 13243 18000 13252
rect 17948 13209 17957 13243
rect 17957 13209 17991 13243
rect 17991 13209 18000 13243
rect 17948 13200 18000 13209
rect 9208 13132 9260 13184
rect 10496 13175 10548 13184
rect 10496 13141 10505 13175
rect 10505 13141 10539 13175
rect 10539 13141 10548 13175
rect 10496 13132 10548 13141
rect 10680 13132 10732 13184
rect 11692 13175 11744 13184
rect 11692 13141 11701 13175
rect 11701 13141 11735 13175
rect 11735 13141 11744 13175
rect 11692 13132 11744 13141
rect 11784 13132 11836 13184
rect 13808 13175 13860 13184
rect 13808 13141 13817 13175
rect 13817 13141 13851 13175
rect 13851 13141 13860 13175
rect 13808 13132 13860 13141
rect 19696 13175 19748 13184
rect 19696 13141 19705 13175
rect 19705 13141 19739 13175
rect 19739 13141 19748 13175
rect 19696 13132 19748 13141
rect 21076 13132 21128 13184
rect 5176 13030 5228 13082
rect 5240 13030 5292 13082
rect 5304 13030 5356 13082
rect 5368 13030 5420 13082
rect 14510 13030 14562 13082
rect 14574 13030 14626 13082
rect 14638 13030 14690 13082
rect 14702 13030 14754 13082
rect 23843 13030 23895 13082
rect 23907 13030 23959 13082
rect 23971 13030 24023 13082
rect 24035 13030 24087 13082
rect 9300 12928 9352 12980
rect 9392 12928 9444 12980
rect 10588 12971 10640 12980
rect 10588 12937 10597 12971
rect 10597 12937 10631 12971
rect 10631 12937 10640 12971
rect 10588 12928 10640 12937
rect 9484 12903 9536 12912
rect 9484 12869 9493 12903
rect 9493 12869 9527 12903
rect 9527 12869 9536 12903
rect 9484 12860 9536 12869
rect 9576 12860 9628 12912
rect 10220 12860 10272 12912
rect 11416 12928 11468 12980
rect 12060 12928 12112 12980
rect 13624 12971 13676 12980
rect 13624 12937 13633 12971
rect 13633 12937 13667 12971
rect 13667 12937 13676 12971
rect 13624 12928 13676 12937
rect 14084 12971 14136 12980
rect 14084 12937 14093 12971
rect 14093 12937 14127 12971
rect 14127 12937 14136 12971
rect 14084 12928 14136 12937
rect 14268 12971 14320 12980
rect 14268 12937 14277 12971
rect 14277 12937 14311 12971
rect 14311 12937 14320 12971
rect 14268 12928 14320 12937
rect 16936 12971 16988 12980
rect 16936 12937 16945 12971
rect 16945 12937 16979 12971
rect 16979 12937 16988 12971
rect 16936 12928 16988 12937
rect 18960 12971 19012 12980
rect 18960 12937 18969 12971
rect 18969 12937 19003 12971
rect 19003 12937 19012 12971
rect 18960 12928 19012 12937
rect 20156 12928 20208 12980
rect 22456 12971 22508 12980
rect 22456 12937 22465 12971
rect 22465 12937 22499 12971
rect 22499 12937 22508 12971
rect 22456 12928 22508 12937
rect 24204 12971 24256 12980
rect 24204 12937 24213 12971
rect 24213 12937 24247 12971
rect 24247 12937 24256 12971
rect 24204 12928 24256 12937
rect 12152 12860 12204 12912
rect 10680 12835 10732 12844
rect 10680 12801 10689 12835
rect 10689 12801 10723 12835
rect 10723 12801 10732 12835
rect 10680 12792 10732 12801
rect 9300 12767 9352 12776
rect 9300 12733 9309 12767
rect 9309 12733 9343 12767
rect 9343 12733 9352 12767
rect 9300 12724 9352 12733
rect 9208 12656 9260 12708
rect 10496 12656 10548 12708
rect 13348 12656 13400 12708
rect 16016 12792 16068 12844
rect 17304 12903 17356 12912
rect 17304 12869 17313 12903
rect 17313 12869 17347 12903
rect 17347 12869 17356 12903
rect 17304 12860 17356 12869
rect 20708 12860 20760 12912
rect 17948 12835 18000 12844
rect 17948 12801 17957 12835
rect 17957 12801 17991 12835
rect 17991 12801 18000 12835
rect 17948 12792 18000 12801
rect 19788 12835 19840 12844
rect 19788 12801 19797 12835
rect 19797 12801 19831 12835
rect 19831 12801 19840 12835
rect 19788 12792 19840 12801
rect 20248 12792 20300 12844
rect 21076 12835 21128 12844
rect 21076 12801 21085 12835
rect 21085 12801 21119 12835
rect 21119 12801 21128 12835
rect 21076 12792 21128 12801
rect 23100 12792 23152 12844
rect 13808 12767 13860 12776
rect 13808 12733 13817 12767
rect 13817 12733 13851 12767
rect 13851 12733 13860 12767
rect 13808 12724 13860 12733
rect 14360 12724 14412 12776
rect 18500 12724 18552 12776
rect 19512 12724 19564 12776
rect 19696 12767 19748 12776
rect 19696 12733 19705 12767
rect 19705 12733 19739 12767
rect 19739 12733 19748 12767
rect 19696 12724 19748 12733
rect 20892 12767 20944 12776
rect 20892 12733 20898 12767
rect 20898 12733 20944 12767
rect 20892 12724 20944 12733
rect 21444 12767 21496 12776
rect 21444 12733 21453 12767
rect 21453 12733 21487 12767
rect 21487 12733 21496 12767
rect 21444 12724 21496 12733
rect 22640 12724 22692 12776
rect 23008 12724 23060 12776
rect 25032 12724 25084 12776
rect 14912 12656 14964 12708
rect 16292 12656 16344 12708
rect 17304 12656 17356 12708
rect 20432 12656 20484 12708
rect 10864 12588 10916 12640
rect 11324 12588 11376 12640
rect 12244 12631 12296 12640
rect 12244 12597 12253 12631
rect 12253 12597 12287 12631
rect 12287 12597 12296 12631
rect 12244 12588 12296 12597
rect 13072 12631 13124 12640
rect 13072 12597 13081 12631
rect 13081 12597 13115 12631
rect 13115 12597 13124 12631
rect 13072 12588 13124 12597
rect 16660 12631 16712 12640
rect 16660 12597 16669 12631
rect 16669 12597 16703 12631
rect 16703 12597 16712 12631
rect 16660 12588 16712 12597
rect 17580 12588 17632 12640
rect 22916 12656 22968 12708
rect 23284 12699 23336 12708
rect 23284 12665 23293 12699
rect 23293 12665 23327 12699
rect 23327 12665 23336 12699
rect 23284 12656 23336 12665
rect 23652 12656 23704 12708
rect 24296 12588 24348 12640
rect 9843 12486 9895 12538
rect 9907 12486 9959 12538
rect 9971 12486 10023 12538
rect 10035 12486 10087 12538
rect 19176 12486 19228 12538
rect 19240 12486 19292 12538
rect 19304 12486 19356 12538
rect 19368 12486 19420 12538
rect 10588 12427 10640 12436
rect 10588 12393 10597 12427
rect 10597 12393 10631 12427
rect 10631 12393 10640 12427
rect 10588 12384 10640 12393
rect 12244 12384 12296 12436
rect 13348 12384 13400 12436
rect 13808 12427 13860 12436
rect 13808 12393 13817 12427
rect 13817 12393 13851 12427
rect 13851 12393 13860 12427
rect 13808 12384 13860 12393
rect 13992 12384 14044 12436
rect 16108 12427 16160 12436
rect 16108 12393 16117 12427
rect 16117 12393 16151 12427
rect 16151 12393 16160 12427
rect 16108 12384 16160 12393
rect 16660 12384 16712 12436
rect 19512 12384 19564 12436
rect 19788 12384 19840 12436
rect 20892 12384 20944 12436
rect 22916 12384 22968 12436
rect 25032 12384 25084 12436
rect 12520 12359 12572 12368
rect 12520 12325 12529 12359
rect 12529 12325 12563 12359
rect 12563 12325 12572 12359
rect 12520 12316 12572 12325
rect 16752 12316 16804 12368
rect 17028 12359 17080 12368
rect 17028 12325 17037 12359
rect 17037 12325 17071 12359
rect 17071 12325 17080 12359
rect 17028 12316 17080 12325
rect 18960 12316 19012 12368
rect 19604 12316 19656 12368
rect 20616 12316 20668 12368
rect 23008 12316 23060 12368
rect 23836 12316 23888 12368
rect 24296 12316 24348 12368
rect 8656 12248 8708 12300
rect 10220 12248 10272 12300
rect 10496 12248 10548 12300
rect 11048 12291 11100 12300
rect 11048 12257 11057 12291
rect 11057 12257 11091 12291
rect 11091 12257 11100 12291
rect 11048 12248 11100 12257
rect 11416 12223 11468 12232
rect 11416 12189 11425 12223
rect 11425 12189 11459 12223
rect 11459 12189 11468 12223
rect 11416 12180 11468 12189
rect 18132 12248 18184 12300
rect 18316 12291 18368 12300
rect 18316 12257 18325 12291
rect 18325 12257 18359 12291
rect 18359 12257 18368 12291
rect 18316 12248 18368 12257
rect 19696 12248 19748 12300
rect 21904 12248 21956 12300
rect 23192 12248 23244 12300
rect 13440 12180 13492 12232
rect 13624 12180 13676 12232
rect 15740 12180 15792 12232
rect 16660 12180 16712 12232
rect 14544 12155 14596 12164
rect 14544 12121 14553 12155
rect 14553 12121 14587 12155
rect 14587 12121 14596 12155
rect 14544 12112 14596 12121
rect 8288 12087 8340 12096
rect 8288 12053 8297 12087
rect 8297 12053 8331 12087
rect 8331 12053 8340 12087
rect 8288 12044 8340 12053
rect 9944 12087 9996 12096
rect 9944 12053 9953 12087
rect 9953 12053 9987 12087
rect 9987 12053 9996 12087
rect 9944 12044 9996 12053
rect 11232 12087 11284 12096
rect 11232 12053 11256 12087
rect 11256 12053 11284 12087
rect 11232 12044 11284 12053
rect 11324 12087 11376 12096
rect 11324 12053 11333 12087
rect 11333 12053 11367 12087
rect 11367 12053 11376 12087
rect 11508 12087 11560 12096
rect 11324 12044 11376 12053
rect 11508 12053 11517 12087
rect 11517 12053 11551 12087
rect 11551 12053 11560 12087
rect 11508 12044 11560 12053
rect 11968 12044 12020 12096
rect 12336 12044 12388 12096
rect 13348 12087 13400 12096
rect 13348 12053 13372 12087
rect 13372 12053 13400 12087
rect 13348 12044 13400 12053
rect 14084 12044 14136 12096
rect 15832 12087 15884 12096
rect 15832 12053 15841 12087
rect 15841 12053 15875 12087
rect 15875 12053 15884 12087
rect 15832 12044 15884 12053
rect 17304 12044 17356 12096
rect 18868 12180 18920 12232
rect 20248 12180 20300 12232
rect 23468 12180 23520 12232
rect 23652 12223 23704 12232
rect 23652 12189 23661 12223
rect 23661 12189 23695 12223
rect 23695 12189 23704 12223
rect 23652 12180 23704 12189
rect 18040 12112 18092 12164
rect 18776 12112 18828 12164
rect 19604 12112 19656 12164
rect 20708 12155 20760 12164
rect 20708 12121 20717 12155
rect 20717 12121 20751 12155
rect 20751 12121 20760 12155
rect 20708 12112 20760 12121
rect 23560 12112 23612 12164
rect 24112 12112 24164 12164
rect 24848 12291 24900 12300
rect 24848 12257 24892 12291
rect 24892 12257 24900 12291
rect 24848 12248 24900 12257
rect 18224 12087 18276 12096
rect 18224 12053 18233 12087
rect 18233 12053 18267 12087
rect 18267 12053 18276 12087
rect 18224 12044 18276 12053
rect 18592 12087 18644 12096
rect 18592 12053 18601 12087
rect 18601 12053 18635 12087
rect 18635 12053 18644 12087
rect 18592 12044 18644 12053
rect 20340 12044 20392 12096
rect 22548 12087 22600 12096
rect 22548 12053 22557 12087
rect 22557 12053 22591 12087
rect 22591 12053 22600 12087
rect 22548 12044 22600 12053
rect 24296 12044 24348 12096
rect 5176 11942 5228 11994
rect 5240 11942 5292 11994
rect 5304 11942 5356 11994
rect 5368 11942 5420 11994
rect 14510 11942 14562 11994
rect 14574 11942 14626 11994
rect 14638 11942 14690 11994
rect 14702 11942 14754 11994
rect 23843 11942 23895 11994
rect 23907 11942 23959 11994
rect 23971 11942 24023 11994
rect 24035 11942 24087 11994
rect 7736 11883 7788 11892
rect 7736 11849 7745 11883
rect 7745 11849 7779 11883
rect 7779 11849 7788 11883
rect 7736 11840 7788 11849
rect 8656 11883 8708 11892
rect 8656 11849 8665 11883
rect 8665 11849 8699 11883
rect 8699 11849 8708 11883
rect 8656 11840 8708 11849
rect 9392 11883 9444 11892
rect 9392 11849 9401 11883
rect 9401 11849 9435 11883
rect 9435 11849 9444 11883
rect 9392 11840 9444 11849
rect 10220 11840 10272 11892
rect 11140 11840 11192 11892
rect 11324 11840 11376 11892
rect 13624 11840 13676 11892
rect 14176 11840 14228 11892
rect 15188 11883 15240 11892
rect 15188 11849 15197 11883
rect 15197 11849 15231 11883
rect 15231 11849 15240 11883
rect 15188 11840 15240 11849
rect 16752 11840 16804 11892
rect 17304 11883 17356 11892
rect 17304 11849 17313 11883
rect 17313 11849 17347 11883
rect 17347 11849 17356 11883
rect 17304 11840 17356 11849
rect 18684 11840 18736 11892
rect 19788 11883 19840 11892
rect 19788 11849 19797 11883
rect 19797 11849 19831 11883
rect 19831 11849 19840 11883
rect 19788 11840 19840 11849
rect 9116 11815 9168 11824
rect 9116 11781 9125 11815
rect 9125 11781 9159 11815
rect 9159 11781 9168 11815
rect 9116 11772 9168 11781
rect 12244 11815 12296 11824
rect 12244 11781 12253 11815
rect 12253 11781 12287 11815
rect 12287 11781 12296 11815
rect 12244 11772 12296 11781
rect 7736 11636 7788 11688
rect 12336 11747 12388 11756
rect 12336 11713 12345 11747
rect 12345 11713 12379 11747
rect 12379 11713 12388 11747
rect 12336 11704 12388 11713
rect 8104 11568 8156 11620
rect 9944 11636 9996 11688
rect 10220 11679 10272 11688
rect 10220 11645 10229 11679
rect 10229 11645 10263 11679
rect 10263 11645 10272 11679
rect 10220 11636 10272 11645
rect 10772 11679 10824 11688
rect 10772 11645 10781 11679
rect 10781 11645 10815 11679
rect 10815 11645 10824 11679
rect 10772 11636 10824 11645
rect 11508 11636 11560 11688
rect 12060 11636 12112 11688
rect 12428 11636 12480 11688
rect 14084 11815 14136 11824
rect 14084 11781 14093 11815
rect 14093 11781 14127 11815
rect 14127 11781 14136 11815
rect 14084 11772 14136 11781
rect 15004 11772 15056 11824
rect 18500 11772 18552 11824
rect 19604 11772 19656 11824
rect 14268 11704 14320 11756
rect 18040 11704 18092 11756
rect 18868 11704 18920 11756
rect 15188 11636 15240 11688
rect 15832 11679 15884 11688
rect 15832 11645 15841 11679
rect 15841 11645 15875 11679
rect 15875 11645 15884 11679
rect 15832 11636 15884 11645
rect 17672 11679 17724 11688
rect 17672 11645 17716 11679
rect 17716 11645 17724 11679
rect 17672 11636 17724 11645
rect 18776 11636 18828 11688
rect 20800 11840 20852 11892
rect 23008 11883 23060 11892
rect 23008 11849 23017 11883
rect 23017 11849 23051 11883
rect 23051 11849 23060 11883
rect 23008 11840 23060 11849
rect 24848 11840 24900 11892
rect 20616 11704 20668 11756
rect 21536 11704 21588 11756
rect 21352 11679 21404 11688
rect 21352 11645 21361 11679
rect 21361 11645 21395 11679
rect 21395 11645 21404 11679
rect 21352 11636 21404 11645
rect 9668 11611 9720 11620
rect 9668 11577 9677 11611
rect 9677 11577 9711 11611
rect 9711 11577 9720 11611
rect 9668 11568 9720 11577
rect 11968 11611 12020 11620
rect 11968 11577 11977 11611
rect 11977 11577 12011 11611
rect 12011 11577 12020 11611
rect 11968 11568 12020 11577
rect 13716 11568 13768 11620
rect 13992 11568 14044 11620
rect 15004 11568 15056 11620
rect 15280 11568 15332 11620
rect 18592 11568 18644 11620
rect 20892 11568 20944 11620
rect 23100 11704 23152 11756
rect 23652 11747 23704 11756
rect 23652 11713 23661 11747
rect 23661 11713 23695 11747
rect 23695 11713 23704 11747
rect 23652 11704 23704 11713
rect 24848 11679 24900 11688
rect 24848 11645 24857 11679
rect 24857 11645 24891 11679
rect 24891 11645 24900 11679
rect 24848 11636 24900 11645
rect 7368 11543 7420 11552
rect 7368 11509 7377 11543
rect 7377 11509 7411 11543
rect 7411 11509 7420 11543
rect 7368 11500 7420 11509
rect 8380 11543 8432 11552
rect 8380 11509 8389 11543
rect 8389 11509 8423 11543
rect 8423 11509 8432 11543
rect 8380 11500 8432 11509
rect 10588 11500 10640 11552
rect 11692 11543 11744 11552
rect 11692 11509 11701 11543
rect 11701 11509 11735 11543
rect 11735 11509 11744 11543
rect 11692 11500 11744 11509
rect 12612 11543 12664 11552
rect 12612 11509 12621 11543
rect 12621 11509 12655 11543
rect 12655 11509 12664 11543
rect 12612 11500 12664 11509
rect 15464 11543 15516 11552
rect 15464 11509 15473 11543
rect 15473 11509 15507 11543
rect 15507 11509 15516 11543
rect 15464 11500 15516 11509
rect 16752 11543 16804 11552
rect 16752 11509 16761 11543
rect 16761 11509 16795 11543
rect 16795 11509 16804 11543
rect 16752 11500 16804 11509
rect 18408 11500 18460 11552
rect 20708 11500 20760 11552
rect 23560 11568 23612 11620
rect 23652 11568 23704 11620
rect 24940 11568 24992 11620
rect 23744 11500 23796 11552
rect 24296 11500 24348 11552
rect 24388 11500 24440 11552
rect 9843 11398 9895 11450
rect 9907 11398 9959 11450
rect 9971 11398 10023 11450
rect 10035 11398 10087 11450
rect 19176 11398 19228 11450
rect 19240 11398 19292 11450
rect 19304 11398 19356 11450
rect 19368 11398 19420 11450
rect 9392 11296 9444 11348
rect 10220 11296 10272 11348
rect 11048 11296 11100 11348
rect 12244 11296 12296 11348
rect 12428 11339 12480 11348
rect 12428 11305 12437 11339
rect 12437 11305 12471 11339
rect 12471 11305 12480 11339
rect 12428 11296 12480 11305
rect 13440 11296 13492 11348
rect 13900 11296 13952 11348
rect 15004 11296 15056 11348
rect 16476 11339 16528 11348
rect 16476 11305 16485 11339
rect 16485 11305 16519 11339
rect 16519 11305 16528 11339
rect 16476 11296 16528 11305
rect 21352 11296 21404 11348
rect 23468 11339 23520 11348
rect 9300 11228 9352 11280
rect 8104 11203 8156 11212
rect 8104 11169 8113 11203
rect 8113 11169 8147 11203
rect 8147 11169 8156 11203
rect 8104 11160 8156 11169
rect 9668 11160 9720 11212
rect 11692 11228 11744 11280
rect 12336 11228 12388 11280
rect 14360 11228 14412 11280
rect 17672 11228 17724 11280
rect 18500 11228 18552 11280
rect 20708 11228 20760 11280
rect 21904 11271 21956 11280
rect 13072 11160 13124 11212
rect 13624 11160 13676 11212
rect 16384 11160 16436 11212
rect 16660 11203 16712 11212
rect 16660 11169 16669 11203
rect 16669 11169 16703 11203
rect 16703 11169 16712 11203
rect 16660 11160 16712 11169
rect 11416 11135 11468 11144
rect 8288 11067 8340 11076
rect 8288 11033 8297 11067
rect 8297 11033 8331 11067
rect 8331 11033 8340 11067
rect 8288 11024 8340 11033
rect 10772 11024 10824 11076
rect 11416 11101 11425 11135
rect 11425 11101 11459 11135
rect 11459 11101 11468 11135
rect 11416 11092 11468 11101
rect 11508 11135 11560 11144
rect 11508 11101 11517 11135
rect 11517 11101 11551 11135
rect 11551 11101 11560 11135
rect 15188 11135 15240 11144
rect 11508 11092 11560 11101
rect 15188 11101 15197 11135
rect 15197 11101 15231 11135
rect 15231 11101 15240 11135
rect 15188 11092 15240 11101
rect 16200 11092 16252 11144
rect 17488 11160 17540 11212
rect 18132 11203 18184 11212
rect 18132 11169 18141 11203
rect 18141 11169 18175 11203
rect 18175 11169 18184 11203
rect 18132 11160 18184 11169
rect 18776 11160 18828 11212
rect 20432 11203 20484 11212
rect 20432 11169 20441 11203
rect 20441 11169 20475 11203
rect 20475 11169 20484 11203
rect 20432 11160 20484 11169
rect 20892 11203 20944 11212
rect 20892 11169 20901 11203
rect 20901 11169 20935 11203
rect 20935 11169 20944 11203
rect 20892 11160 20944 11169
rect 18040 11092 18092 11144
rect 18960 11092 19012 11144
rect 20984 11135 21036 11144
rect 20984 11101 20993 11135
rect 20993 11101 21027 11135
rect 21027 11101 21036 11135
rect 20984 11092 21036 11101
rect 21904 11237 21913 11271
rect 21913 11237 21947 11271
rect 21947 11237 21956 11271
rect 21904 11228 21956 11237
rect 22732 11228 22784 11280
rect 23468 11305 23477 11339
rect 23477 11305 23511 11339
rect 23511 11305 23520 11339
rect 23468 11296 23520 11305
rect 24480 11203 24532 11212
rect 22640 11092 22692 11144
rect 22916 11092 22968 11144
rect 11232 11067 11284 11076
rect 11232 11033 11256 11067
rect 11256 11033 11284 11067
rect 11232 11024 11284 11033
rect 11784 11024 11836 11076
rect 13900 11024 13952 11076
rect 16108 11024 16160 11076
rect 18224 11024 18276 11076
rect 19144 11067 19196 11076
rect 11324 10999 11376 11008
rect 11324 10965 11333 10999
rect 11333 10965 11367 10999
rect 11367 10965 11376 10999
rect 11324 10956 11376 10965
rect 14912 10956 14964 11008
rect 15280 10999 15332 11008
rect 15280 10965 15289 10999
rect 15289 10965 15323 10999
rect 15323 10965 15332 10999
rect 15280 10956 15332 10965
rect 18500 10999 18552 11008
rect 18500 10965 18509 10999
rect 18509 10965 18543 10999
rect 18543 10965 18552 10999
rect 18500 10956 18552 10965
rect 18684 10956 18736 11008
rect 19144 11033 19153 11067
rect 19153 11033 19187 11067
rect 19187 11033 19196 11067
rect 19144 11024 19196 11033
rect 24480 11169 24489 11203
rect 24489 11169 24523 11203
rect 24523 11169 24532 11203
rect 24480 11160 24532 11169
rect 19420 10956 19472 11008
rect 24388 10956 24440 11008
rect 5176 10854 5228 10906
rect 5240 10854 5292 10906
rect 5304 10854 5356 10906
rect 5368 10854 5420 10906
rect 14510 10854 14562 10906
rect 14574 10854 14626 10906
rect 14638 10854 14690 10906
rect 14702 10854 14754 10906
rect 23843 10854 23895 10906
rect 23907 10854 23959 10906
rect 23971 10854 24023 10906
rect 24035 10854 24087 10906
rect 8104 10795 8156 10804
rect 8104 10761 8113 10795
rect 8113 10761 8147 10795
rect 8147 10761 8156 10795
rect 8104 10752 8156 10761
rect 9668 10752 9720 10804
rect 11324 10795 11376 10804
rect 11324 10761 11333 10795
rect 11333 10761 11367 10795
rect 11367 10761 11376 10795
rect 11324 10752 11376 10761
rect 11692 10795 11744 10804
rect 11692 10761 11701 10795
rect 11701 10761 11735 10795
rect 11735 10761 11744 10795
rect 11692 10752 11744 10761
rect 13072 10795 13124 10804
rect 13072 10761 13081 10795
rect 13081 10761 13115 10795
rect 13115 10761 13124 10795
rect 13072 10752 13124 10761
rect 13440 10795 13492 10804
rect 13440 10761 13449 10795
rect 13449 10761 13483 10795
rect 13483 10761 13492 10795
rect 13440 10752 13492 10761
rect 13808 10795 13860 10804
rect 13808 10761 13817 10795
rect 13817 10761 13851 10795
rect 13851 10761 13860 10795
rect 13808 10752 13860 10761
rect 14176 10795 14228 10804
rect 14176 10761 14200 10795
rect 14200 10761 14228 10795
rect 14176 10752 14228 10761
rect 14912 10752 14964 10804
rect 16108 10752 16160 10804
rect 17304 10752 17356 10804
rect 18684 10752 18736 10804
rect 19512 10752 19564 10804
rect 21904 10752 21956 10804
rect 22732 10752 22784 10804
rect 24480 10752 24532 10804
rect 8472 10727 8524 10736
rect 8472 10693 8481 10727
rect 8481 10693 8515 10727
rect 8515 10693 8524 10727
rect 8472 10684 8524 10693
rect 12520 10616 12572 10668
rect 10312 10591 10364 10600
rect 10312 10557 10321 10591
rect 10321 10557 10355 10591
rect 10355 10557 10364 10591
rect 10312 10548 10364 10557
rect 10772 10591 10824 10600
rect 10772 10557 10781 10591
rect 10781 10557 10815 10591
rect 10815 10557 10824 10591
rect 10772 10548 10824 10557
rect 9208 10480 9260 10532
rect 11048 10523 11100 10532
rect 11048 10489 11057 10523
rect 11057 10489 11091 10523
rect 11091 10489 11100 10523
rect 11048 10480 11100 10489
rect 11232 10480 11284 10532
rect 12152 10523 12204 10532
rect 12152 10489 12161 10523
rect 12161 10489 12195 10523
rect 12195 10489 12204 10523
rect 12152 10480 12204 10489
rect 12796 10480 12848 10532
rect 13900 10684 13952 10736
rect 19420 10727 19472 10736
rect 19420 10693 19429 10727
rect 19429 10693 19463 10727
rect 19463 10693 19472 10727
rect 19420 10684 19472 10693
rect 19696 10684 19748 10736
rect 21536 10684 21588 10736
rect 24388 10727 24440 10736
rect 15188 10616 15240 10668
rect 18960 10616 19012 10668
rect 20616 10659 20668 10668
rect 20616 10625 20625 10659
rect 20625 10625 20659 10659
rect 20659 10625 20668 10659
rect 21260 10659 21312 10668
rect 20616 10616 20668 10625
rect 13440 10548 13492 10600
rect 17580 10591 17632 10600
rect 9484 10455 9536 10464
rect 9484 10421 9493 10455
rect 9493 10421 9527 10455
rect 9527 10421 9536 10455
rect 9484 10412 9536 10421
rect 14636 10455 14688 10464
rect 14636 10421 14645 10455
rect 14645 10421 14679 10455
rect 14679 10421 14688 10455
rect 14636 10412 14688 10421
rect 15372 10455 15424 10464
rect 15372 10421 15381 10455
rect 15381 10421 15415 10455
rect 15415 10421 15424 10455
rect 17580 10557 17589 10591
rect 17589 10557 17623 10591
rect 17623 10557 17632 10591
rect 17580 10548 17632 10557
rect 18040 10591 18092 10600
rect 18040 10557 18049 10591
rect 18049 10557 18083 10591
rect 18083 10557 18092 10591
rect 18040 10548 18092 10557
rect 21260 10625 21269 10659
rect 21269 10625 21303 10659
rect 21303 10625 21312 10659
rect 21260 10616 21312 10625
rect 24388 10693 24397 10727
rect 24397 10693 24431 10727
rect 24431 10693 24440 10727
rect 24388 10684 24440 10693
rect 20892 10548 20944 10600
rect 17212 10480 17264 10532
rect 17488 10480 17540 10532
rect 18316 10523 18368 10532
rect 18316 10489 18325 10523
rect 18325 10489 18359 10523
rect 18359 10489 18368 10523
rect 18316 10480 18368 10489
rect 18500 10480 18552 10532
rect 19880 10523 19932 10532
rect 19880 10489 19889 10523
rect 19889 10489 19923 10523
rect 19923 10489 19932 10523
rect 19880 10480 19932 10489
rect 22548 10523 22600 10532
rect 22548 10489 22557 10523
rect 22557 10489 22591 10523
rect 22591 10489 22600 10523
rect 24940 10591 24992 10600
rect 24940 10557 24949 10591
rect 24949 10557 24983 10591
rect 24983 10557 24992 10591
rect 24940 10548 24992 10557
rect 22548 10480 22600 10489
rect 15372 10412 15424 10421
rect 16660 10412 16712 10464
rect 16936 10455 16988 10464
rect 16936 10421 16945 10455
rect 16945 10421 16979 10455
rect 16979 10421 16988 10455
rect 16936 10412 16988 10421
rect 24112 10455 24164 10464
rect 24112 10421 24121 10455
rect 24121 10421 24155 10455
rect 24155 10421 24164 10455
rect 24112 10412 24164 10421
rect 24480 10412 24532 10464
rect 9843 10310 9895 10362
rect 9907 10310 9959 10362
rect 9971 10310 10023 10362
rect 10035 10310 10087 10362
rect 19176 10310 19228 10362
rect 19240 10310 19292 10362
rect 19304 10310 19356 10362
rect 19368 10310 19420 10362
rect 10772 10208 10824 10260
rect 11232 10251 11284 10260
rect 11232 10217 11241 10251
rect 11241 10217 11275 10251
rect 11275 10217 11284 10251
rect 11232 10208 11284 10217
rect 11416 10208 11468 10260
rect 12060 10208 12112 10260
rect 12152 10208 12204 10260
rect 14176 10251 14228 10260
rect 14176 10217 14185 10251
rect 14185 10217 14219 10251
rect 14219 10217 14228 10251
rect 14176 10208 14228 10217
rect 14360 10208 14412 10260
rect 16200 10251 16252 10260
rect 16200 10217 16209 10251
rect 16209 10217 16243 10251
rect 16243 10217 16252 10251
rect 16200 10208 16252 10217
rect 17580 10251 17632 10260
rect 17580 10217 17589 10251
rect 17589 10217 17623 10251
rect 17623 10217 17632 10251
rect 17580 10208 17632 10217
rect 18960 10208 19012 10260
rect 19512 10251 19564 10260
rect 19512 10217 19521 10251
rect 19521 10217 19555 10251
rect 19555 10217 19564 10251
rect 19512 10208 19564 10217
rect 19696 10208 19748 10260
rect 20156 10208 20208 10260
rect 20432 10208 20484 10260
rect 21904 10251 21956 10260
rect 21904 10217 21913 10251
rect 21913 10217 21947 10251
rect 21947 10217 21956 10251
rect 21904 10208 21956 10217
rect 22640 10208 22692 10260
rect 10680 10183 10732 10192
rect 10680 10149 10683 10183
rect 10683 10149 10717 10183
rect 10717 10149 10732 10183
rect 10680 10140 10732 10149
rect 16292 10140 16344 10192
rect 16752 10183 16804 10192
rect 16752 10149 16755 10183
rect 16755 10149 16789 10183
rect 16789 10149 16804 10183
rect 16752 10140 16804 10149
rect 9208 10072 9260 10124
rect 10496 10072 10548 10124
rect 13532 10072 13584 10124
rect 13992 10072 14044 10124
rect 9484 10004 9536 10056
rect 10404 10004 10456 10056
rect 12796 10004 12848 10056
rect 12704 9979 12756 9988
rect 12704 9945 12713 9979
rect 12713 9945 12747 9979
rect 12747 9945 12756 9979
rect 12704 9936 12756 9945
rect 13900 9936 13952 9988
rect 14912 10072 14964 10124
rect 15280 10115 15332 10124
rect 15280 10081 15289 10115
rect 15289 10081 15323 10115
rect 15323 10081 15332 10115
rect 15280 10072 15332 10081
rect 16476 10072 16528 10124
rect 18500 10140 18552 10192
rect 21536 10140 21588 10192
rect 24112 10140 24164 10192
rect 16016 10004 16068 10056
rect 10312 9868 10364 9920
rect 11784 9868 11836 9920
rect 13808 9911 13860 9920
rect 13808 9877 13817 9911
rect 13817 9877 13851 9911
rect 13851 9877 13860 9911
rect 13808 9868 13860 9877
rect 16936 9936 16988 9988
rect 14912 9868 14964 9920
rect 15832 9911 15884 9920
rect 15832 9877 15841 9911
rect 15841 9877 15875 9911
rect 15875 9877 15884 9911
rect 15832 9868 15884 9877
rect 17396 9868 17448 9920
rect 17856 9868 17908 9920
rect 18684 10072 18736 10124
rect 20984 10115 21036 10124
rect 20984 10081 20993 10115
rect 20993 10081 21027 10115
rect 21027 10081 21036 10115
rect 20984 10072 21036 10081
rect 21628 10072 21680 10124
rect 23468 10072 23520 10124
rect 18960 10004 19012 10056
rect 22088 10004 22140 10056
rect 24572 10004 24624 10056
rect 24756 10047 24808 10056
rect 24756 10013 24765 10047
rect 24765 10013 24799 10047
rect 24799 10013 24808 10047
rect 24756 10004 24808 10013
rect 18408 9911 18460 9920
rect 18408 9877 18417 9911
rect 18417 9877 18451 9911
rect 18451 9877 18460 9911
rect 18408 9868 18460 9877
rect 18592 9911 18644 9920
rect 18592 9877 18601 9911
rect 18601 9877 18635 9911
rect 18635 9877 18644 9911
rect 18592 9868 18644 9877
rect 23560 9868 23612 9920
rect 5176 9766 5228 9818
rect 5240 9766 5292 9818
rect 5304 9766 5356 9818
rect 5368 9766 5420 9818
rect 14510 9766 14562 9818
rect 14574 9766 14626 9818
rect 14638 9766 14690 9818
rect 14702 9766 14754 9818
rect 23843 9766 23895 9818
rect 23907 9766 23959 9818
rect 23971 9766 24023 9818
rect 24035 9766 24087 9818
rect 7276 9664 7328 9716
rect 8196 9664 8248 9716
rect 9208 9664 9260 9716
rect 9484 9596 9536 9648
rect 10220 9596 10272 9648
rect 11232 9664 11284 9716
rect 10588 9596 10640 9648
rect 12060 9596 12112 9648
rect 13532 9664 13584 9716
rect 14912 9707 14964 9716
rect 14912 9673 14921 9707
rect 14921 9673 14955 9707
rect 14955 9673 14964 9707
rect 14912 9664 14964 9673
rect 15004 9664 15056 9716
rect 17304 9707 17356 9716
rect 17304 9673 17313 9707
rect 17313 9673 17347 9707
rect 17347 9673 17356 9707
rect 17304 9664 17356 9673
rect 18408 9664 18460 9716
rect 15924 9596 15976 9648
rect 18960 9707 19012 9716
rect 18960 9673 18969 9707
rect 18969 9673 19003 9707
rect 19003 9673 19012 9707
rect 18960 9664 19012 9673
rect 19512 9664 19564 9716
rect 21628 9664 21680 9716
rect 21812 9664 21864 9716
rect 22180 9664 22232 9716
rect 9300 9528 9352 9580
rect 10680 9528 10732 9580
rect 12796 9528 12848 9580
rect 16844 9528 16896 9580
rect 17672 9571 17724 9580
rect 17672 9537 17681 9571
rect 17681 9537 17715 9571
rect 17715 9537 17724 9571
rect 17672 9528 17724 9537
rect 9484 9460 9536 9512
rect 13716 9503 13768 9512
rect 13716 9469 13725 9503
rect 13725 9469 13759 9503
rect 13759 9469 13768 9503
rect 13716 9460 13768 9469
rect 10404 9435 10456 9444
rect 10404 9401 10413 9435
rect 10413 9401 10447 9435
rect 10447 9401 10456 9435
rect 10404 9392 10456 9401
rect 10496 9435 10548 9444
rect 10496 9401 10505 9435
rect 10505 9401 10539 9435
rect 10539 9401 10548 9435
rect 10496 9392 10548 9401
rect 13808 9392 13860 9444
rect 13992 9460 14044 9512
rect 20800 9639 20852 9648
rect 20800 9605 20809 9639
rect 20809 9605 20843 9639
rect 20843 9605 20852 9639
rect 20800 9596 20852 9605
rect 21536 9596 21588 9648
rect 21260 9571 21312 9580
rect 21260 9537 21269 9571
rect 21269 9537 21303 9571
rect 21303 9537 21312 9571
rect 21260 9528 21312 9537
rect 18960 9460 19012 9512
rect 22640 9460 22692 9512
rect 23376 9460 23428 9512
rect 15832 9392 15884 9444
rect 17396 9392 17448 9444
rect 11968 9367 12020 9376
rect 11968 9333 11977 9367
rect 11977 9333 12011 9367
rect 12011 9333 12020 9367
rect 11968 9324 12020 9333
rect 14728 9324 14780 9376
rect 16752 9324 16804 9376
rect 17856 9392 17908 9444
rect 18868 9392 18920 9444
rect 21536 9392 21588 9444
rect 23928 9392 23980 9444
rect 24848 9503 24900 9512
rect 24848 9469 24857 9503
rect 24857 9469 24891 9503
rect 24891 9469 24900 9503
rect 24848 9460 24900 9469
rect 24296 9435 24348 9444
rect 24296 9401 24305 9435
rect 24305 9401 24339 9435
rect 24339 9401 24348 9435
rect 24296 9392 24348 9401
rect 24572 9392 24624 9444
rect 18408 9324 18460 9376
rect 19788 9367 19840 9376
rect 19788 9333 19797 9367
rect 19797 9333 19831 9367
rect 19831 9333 19840 9367
rect 19788 9324 19840 9333
rect 23468 9367 23520 9376
rect 23468 9333 23477 9367
rect 23477 9333 23511 9367
rect 23511 9333 23520 9367
rect 23468 9324 23520 9333
rect 9843 9222 9895 9274
rect 9907 9222 9959 9274
rect 9971 9222 10023 9274
rect 10035 9222 10087 9274
rect 19176 9222 19228 9274
rect 19240 9222 19292 9274
rect 19304 9222 19356 9274
rect 19368 9222 19420 9274
rect 10404 9120 10456 9172
rect 12060 9163 12112 9172
rect 12060 9129 12069 9163
rect 12069 9129 12103 9163
rect 12103 9129 12112 9163
rect 12060 9120 12112 9129
rect 12520 9120 12572 9172
rect 12796 9163 12848 9172
rect 12796 9129 12805 9163
rect 12805 9129 12839 9163
rect 12839 9129 12848 9163
rect 12796 9120 12848 9129
rect 14636 9163 14688 9172
rect 14636 9129 14645 9163
rect 14645 9129 14679 9163
rect 14679 9129 14688 9163
rect 14636 9120 14688 9129
rect 16476 9163 16528 9172
rect 16476 9129 16485 9163
rect 16485 9129 16519 9163
rect 16519 9129 16528 9163
rect 16476 9120 16528 9129
rect 18684 9120 18736 9172
rect 18960 9120 19012 9172
rect 19604 9120 19656 9172
rect 20984 9120 21036 9172
rect 21352 9120 21404 9172
rect 24204 9120 24256 9172
rect 10680 9052 10732 9104
rect 11232 9052 11284 9104
rect 13072 9095 13124 9104
rect 13072 9061 13081 9095
rect 13081 9061 13115 9095
rect 13115 9061 13124 9095
rect 13072 9052 13124 9061
rect 10220 9027 10272 9036
rect 10220 8993 10229 9027
rect 10229 8993 10263 9027
rect 10263 8993 10272 9027
rect 10220 8984 10272 8993
rect 10496 8984 10548 9036
rect 11048 8984 11100 9036
rect 13716 8984 13768 9036
rect 15004 9052 15056 9104
rect 15556 9052 15608 9104
rect 16844 9095 16896 9104
rect 16844 9061 16853 9095
rect 16853 9061 16887 9095
rect 16887 9061 16896 9095
rect 16844 9052 16896 9061
rect 17580 9052 17632 9104
rect 18868 9052 18920 9104
rect 21444 9095 21496 9104
rect 21444 9061 21453 9095
rect 21453 9061 21487 9095
rect 21487 9061 21496 9095
rect 21444 9052 21496 9061
rect 22916 9095 22968 9104
rect 22916 9061 22925 9095
rect 22925 9061 22959 9095
rect 22959 9061 22968 9095
rect 22916 9052 22968 9061
rect 23376 9052 23428 9104
rect 24296 9052 24348 9104
rect 14912 8984 14964 9036
rect 19696 8984 19748 9036
rect 11968 8916 12020 8968
rect 12980 8959 13032 8968
rect 12980 8925 12989 8959
rect 12989 8925 13023 8959
rect 13023 8925 13032 8959
rect 12980 8916 13032 8925
rect 13348 8959 13400 8968
rect 13348 8925 13357 8959
rect 13357 8925 13391 8959
rect 13391 8925 13400 8959
rect 13348 8916 13400 8925
rect 13808 8916 13860 8968
rect 16936 8916 16988 8968
rect 17856 8959 17908 8968
rect 17856 8925 17865 8959
rect 17865 8925 17899 8959
rect 17899 8925 17908 8959
rect 17856 8916 17908 8925
rect 21536 8916 21588 8968
rect 23192 8959 23244 8968
rect 23192 8925 23201 8959
rect 23201 8925 23235 8959
rect 23235 8925 23244 8959
rect 23192 8916 23244 8925
rect 15648 8891 15700 8900
rect 15648 8857 15657 8891
rect 15657 8857 15691 8891
rect 15691 8857 15700 8891
rect 15648 8848 15700 8857
rect 17672 8848 17724 8900
rect 13900 8823 13952 8832
rect 13900 8789 13909 8823
rect 13909 8789 13943 8823
rect 13943 8789 13952 8823
rect 13900 8780 13952 8789
rect 20892 8823 20944 8832
rect 20892 8789 20901 8823
rect 20901 8789 20935 8823
rect 20935 8789 20944 8823
rect 20892 8780 20944 8789
rect 23468 8780 23520 8832
rect 25124 8780 25176 8832
rect 5176 8678 5228 8730
rect 5240 8678 5292 8730
rect 5304 8678 5356 8730
rect 5368 8678 5420 8730
rect 14510 8678 14562 8730
rect 14574 8678 14626 8730
rect 14638 8678 14690 8730
rect 14702 8678 14754 8730
rect 23843 8678 23895 8730
rect 23907 8678 23959 8730
rect 23971 8678 24023 8730
rect 24035 8678 24087 8730
rect 10220 8576 10272 8628
rect 11232 8619 11284 8628
rect 11232 8585 11241 8619
rect 11241 8585 11275 8619
rect 11275 8585 11284 8619
rect 11232 8576 11284 8585
rect 13440 8619 13492 8628
rect 13440 8585 13449 8619
rect 13449 8585 13483 8619
rect 13483 8585 13492 8619
rect 13440 8576 13492 8585
rect 15004 8619 15056 8628
rect 15004 8585 15013 8619
rect 15013 8585 15047 8619
rect 15047 8585 15056 8619
rect 15004 8576 15056 8585
rect 15740 8576 15792 8628
rect 16936 8619 16988 8628
rect 16936 8585 16945 8619
rect 16945 8585 16979 8619
rect 16979 8585 16988 8619
rect 16936 8576 16988 8585
rect 9392 8508 9444 8560
rect 12060 8508 12112 8560
rect 14268 8551 14320 8560
rect 14268 8517 14277 8551
rect 14277 8517 14311 8551
rect 14311 8517 14320 8551
rect 14268 8508 14320 8517
rect 10496 8483 10548 8492
rect 10496 8449 10505 8483
rect 10505 8449 10539 8483
rect 10539 8449 10548 8483
rect 10496 8440 10548 8449
rect 10404 8415 10456 8424
rect 10404 8381 10413 8415
rect 10413 8381 10447 8415
rect 10447 8381 10456 8415
rect 10404 8372 10456 8381
rect 13072 8440 13124 8492
rect 15648 8440 15700 8492
rect 16108 8440 16160 8492
rect 17580 8483 17632 8492
rect 17580 8449 17589 8483
rect 17589 8449 17623 8483
rect 17623 8449 17632 8483
rect 17580 8440 17632 8449
rect 13440 8372 13492 8424
rect 13808 8372 13860 8424
rect 16384 8415 16436 8424
rect 8932 8347 8984 8356
rect 8932 8313 8941 8347
rect 8941 8313 8975 8347
rect 8975 8313 8984 8347
rect 8932 8304 8984 8313
rect 13900 8304 13952 8356
rect 16384 8381 16393 8415
rect 16393 8381 16427 8415
rect 16427 8381 16436 8415
rect 16384 8372 16436 8381
rect 18408 8372 18460 8424
rect 18960 8372 19012 8424
rect 19972 8576 20024 8628
rect 20156 8576 20208 8628
rect 20616 8576 20668 8628
rect 19788 8415 19840 8424
rect 19788 8381 19797 8415
rect 19797 8381 19831 8415
rect 19831 8381 19840 8415
rect 19788 8372 19840 8381
rect 20248 8372 20300 8424
rect 21444 8576 21496 8628
rect 21904 8619 21956 8628
rect 21904 8585 21913 8619
rect 21913 8585 21947 8619
rect 21947 8585 21956 8619
rect 21904 8576 21956 8585
rect 22640 8619 22692 8628
rect 22640 8585 22649 8619
rect 22649 8585 22683 8619
rect 22683 8585 22692 8619
rect 22640 8576 22692 8585
rect 23008 8619 23060 8628
rect 23008 8585 23017 8619
rect 23017 8585 23051 8619
rect 23051 8585 23060 8619
rect 23008 8576 23060 8585
rect 23376 8576 23428 8628
rect 24204 8576 24256 8628
rect 24940 8619 24992 8628
rect 24940 8585 24949 8619
rect 24949 8585 24983 8619
rect 24983 8585 24992 8619
rect 24940 8576 24992 8585
rect 23192 8508 23244 8560
rect 24204 8440 24256 8492
rect 24480 8440 24532 8492
rect 20984 8372 21036 8424
rect 24756 8415 24808 8424
rect 24756 8381 24765 8415
rect 24765 8381 24799 8415
rect 24799 8381 24808 8415
rect 24756 8372 24808 8381
rect 15372 8347 15424 8356
rect 15372 8313 15381 8347
rect 15381 8313 15415 8347
rect 15415 8313 15424 8347
rect 15372 8304 15424 8313
rect 16752 8304 16804 8356
rect 20064 8347 20116 8356
rect 20064 8313 20073 8347
rect 20073 8313 20107 8347
rect 20107 8313 20116 8347
rect 20064 8304 20116 8313
rect 23284 8347 23336 8356
rect 23284 8313 23293 8347
rect 23293 8313 23327 8347
rect 23327 8313 23336 8347
rect 23284 8304 23336 8313
rect 23376 8347 23428 8356
rect 23376 8313 23385 8347
rect 23385 8313 23419 8347
rect 23419 8313 23428 8347
rect 23376 8304 23428 8313
rect 21168 8279 21220 8288
rect 21168 8245 21177 8279
rect 21177 8245 21211 8279
rect 21211 8245 21220 8279
rect 21168 8236 21220 8245
rect 9843 8134 9895 8186
rect 9907 8134 9959 8186
rect 9971 8134 10023 8186
rect 10035 8134 10087 8186
rect 19176 8134 19228 8186
rect 19240 8134 19292 8186
rect 19304 8134 19356 8186
rect 19368 8134 19420 8186
rect 10404 8032 10456 8084
rect 10588 8075 10640 8084
rect 10588 8041 10597 8075
rect 10597 8041 10631 8075
rect 10631 8041 10640 8075
rect 10588 8032 10640 8041
rect 11048 8032 11100 8084
rect 12612 8032 12664 8084
rect 12980 8075 13032 8084
rect 12980 8041 12989 8075
rect 12989 8041 13023 8075
rect 13023 8041 13032 8075
rect 12980 8032 13032 8041
rect 13808 8032 13860 8084
rect 14360 8032 14412 8084
rect 14912 8032 14964 8084
rect 15832 8032 15884 8084
rect 16108 8032 16160 8084
rect 17764 8075 17816 8084
rect 17764 8041 17773 8075
rect 17773 8041 17807 8075
rect 17807 8041 17816 8075
rect 17764 8032 17816 8041
rect 18408 8075 18460 8084
rect 18408 8041 18417 8075
rect 18417 8041 18451 8075
rect 18451 8041 18460 8075
rect 18408 8032 18460 8041
rect 19696 8032 19748 8084
rect 21628 8075 21680 8084
rect 21628 8041 21637 8075
rect 21637 8041 21671 8075
rect 21671 8041 21680 8075
rect 23284 8075 23336 8084
rect 21628 8032 21680 8041
rect 23284 8041 23293 8075
rect 23293 8041 23327 8075
rect 23327 8041 23336 8075
rect 23284 8032 23336 8041
rect 15372 7964 15424 8016
rect 16936 7964 16988 8016
rect 20800 8007 20852 8016
rect 20800 7973 20803 8007
rect 20803 7973 20837 8007
rect 20837 7973 20852 8007
rect 20800 7964 20852 7973
rect 22456 7964 22508 8016
rect 8196 7939 8248 7948
rect 8196 7905 8205 7939
rect 8205 7905 8239 7939
rect 8239 7905 8248 7939
rect 8196 7896 8248 7905
rect 9392 7896 9444 7948
rect 10772 7896 10824 7948
rect 11508 7896 11560 7948
rect 12520 7896 12572 7948
rect 13256 7939 13308 7948
rect 13256 7905 13265 7939
rect 13265 7905 13299 7939
rect 13299 7905 13308 7939
rect 13256 7896 13308 7905
rect 14636 7896 14688 7948
rect 14820 7939 14872 7948
rect 14820 7905 14829 7939
rect 14829 7905 14863 7939
rect 14863 7905 14872 7939
rect 14820 7896 14872 7905
rect 16200 7896 16252 7948
rect 17028 7896 17080 7948
rect 18960 7939 19012 7948
rect 18960 7905 18969 7939
rect 18969 7905 19003 7939
rect 19003 7905 19012 7939
rect 18960 7896 19012 7905
rect 19052 7896 19104 7948
rect 23192 7896 23244 7948
rect 8288 7871 8340 7880
rect 8288 7837 8297 7871
rect 8297 7837 8331 7871
rect 8331 7837 8340 7871
rect 8288 7828 8340 7837
rect 10404 7828 10456 7880
rect 13900 7871 13952 7880
rect 13900 7837 13909 7871
rect 13909 7837 13943 7871
rect 13943 7837 13952 7871
rect 13900 7828 13952 7837
rect 14360 7828 14412 7880
rect 20892 7828 20944 7880
rect 22364 7828 22416 7880
rect 22548 7871 22600 7880
rect 22548 7837 22557 7871
rect 22557 7837 22591 7871
rect 22591 7837 22600 7871
rect 22548 7828 22600 7837
rect 23744 7871 23796 7880
rect 23744 7837 23753 7871
rect 23753 7837 23787 7871
rect 23787 7837 23796 7871
rect 23744 7828 23796 7837
rect 12336 7760 12388 7812
rect 18132 7735 18184 7744
rect 18132 7701 18141 7735
rect 18141 7701 18175 7735
rect 18175 7701 18184 7735
rect 18132 7692 18184 7701
rect 21352 7735 21404 7744
rect 21352 7701 21361 7735
rect 21361 7701 21395 7735
rect 21395 7701 21404 7735
rect 21352 7692 21404 7701
rect 5176 7590 5228 7642
rect 5240 7590 5292 7642
rect 5304 7590 5356 7642
rect 5368 7590 5420 7642
rect 14510 7590 14562 7642
rect 14574 7590 14626 7642
rect 14638 7590 14690 7642
rect 14702 7590 14754 7642
rect 23843 7590 23895 7642
rect 23907 7590 23959 7642
rect 23971 7590 24023 7642
rect 24035 7590 24087 7642
rect 8196 7488 8248 7540
rect 10312 7488 10364 7540
rect 7736 7395 7788 7404
rect 7736 7361 7745 7395
rect 7745 7361 7779 7395
rect 7779 7361 7788 7395
rect 7736 7352 7788 7361
rect 9392 7352 9444 7404
rect 9300 7327 9352 7336
rect 9300 7293 9309 7327
rect 9309 7293 9343 7327
rect 9343 7293 9352 7327
rect 9300 7284 9352 7293
rect 10312 7327 10364 7336
rect 10312 7293 10321 7327
rect 10321 7293 10355 7327
rect 10355 7293 10364 7327
rect 10312 7284 10364 7293
rect 11508 7488 11560 7540
rect 13256 7488 13308 7540
rect 13440 7488 13492 7540
rect 15372 7531 15424 7540
rect 15372 7497 15381 7531
rect 15381 7497 15415 7531
rect 15415 7497 15424 7531
rect 15372 7488 15424 7497
rect 15832 7488 15884 7540
rect 17028 7488 17080 7540
rect 18960 7488 19012 7540
rect 14636 7463 14688 7472
rect 14636 7429 14645 7463
rect 14645 7429 14679 7463
rect 14679 7429 14688 7463
rect 14636 7420 14688 7429
rect 17856 7395 17908 7404
rect 10220 7216 10272 7268
rect 11048 7259 11100 7268
rect 11048 7225 11057 7259
rect 11057 7225 11091 7259
rect 11091 7225 11100 7259
rect 11048 7216 11100 7225
rect 12612 7284 12664 7336
rect 14360 7327 14412 7336
rect 14360 7293 14369 7327
rect 14369 7293 14403 7327
rect 14403 7293 14412 7327
rect 14360 7284 14412 7293
rect 17856 7361 17865 7395
rect 17865 7361 17899 7395
rect 17899 7361 17908 7395
rect 17856 7352 17908 7361
rect 18408 7395 18460 7404
rect 18408 7361 18417 7395
rect 18417 7361 18451 7395
rect 18451 7361 18460 7395
rect 18408 7352 18460 7361
rect 20156 7488 20208 7540
rect 20800 7488 20852 7540
rect 20156 7395 20208 7404
rect 20156 7361 20165 7395
rect 20165 7361 20199 7395
rect 20199 7361 20208 7395
rect 20156 7352 20208 7361
rect 14912 7284 14964 7336
rect 15832 7284 15884 7336
rect 19604 7327 19656 7336
rect 19604 7293 19613 7327
rect 19613 7293 19647 7327
rect 19647 7293 19656 7327
rect 19604 7284 19656 7293
rect 19788 7284 19840 7336
rect 21352 7488 21404 7540
rect 22456 7531 22508 7540
rect 22456 7497 22465 7531
rect 22465 7497 22499 7531
rect 22499 7497 22508 7531
rect 22456 7488 22508 7497
rect 21168 7395 21220 7404
rect 21168 7361 21177 7395
rect 21177 7361 21211 7395
rect 21211 7361 21220 7395
rect 21168 7352 21220 7361
rect 22548 7352 22600 7404
rect 23560 7395 23612 7404
rect 23560 7361 23569 7395
rect 23569 7361 23603 7395
rect 23603 7361 23612 7395
rect 23560 7352 23612 7361
rect 24756 7327 24808 7336
rect 16936 7259 16988 7268
rect 16936 7225 16945 7259
rect 16945 7225 16979 7259
rect 16979 7225 16988 7259
rect 16936 7216 16988 7225
rect 18132 7259 18184 7268
rect 18132 7225 18141 7259
rect 18141 7225 18175 7259
rect 18175 7225 18184 7259
rect 18132 7216 18184 7225
rect 11692 7191 11744 7200
rect 11692 7157 11701 7191
rect 11701 7157 11735 7191
rect 11735 7157 11744 7191
rect 11692 7148 11744 7157
rect 11968 7148 12020 7200
rect 16108 7191 16160 7200
rect 16108 7157 16117 7191
rect 16117 7157 16151 7191
rect 16151 7157 16160 7191
rect 16108 7148 16160 7157
rect 17856 7148 17908 7200
rect 20984 7216 21036 7268
rect 24756 7293 24765 7327
rect 24765 7293 24799 7327
rect 24799 7293 24808 7327
rect 24756 7284 24808 7293
rect 24664 7216 24716 7268
rect 23192 7148 23244 7200
rect 23744 7148 23796 7200
rect 24940 7191 24992 7200
rect 24940 7157 24949 7191
rect 24949 7157 24983 7191
rect 24983 7157 24992 7191
rect 24940 7148 24992 7157
rect 9843 7046 9895 7098
rect 9907 7046 9959 7098
rect 9971 7046 10023 7098
rect 10035 7046 10087 7098
rect 19176 7046 19228 7098
rect 19240 7046 19292 7098
rect 19304 7046 19356 7098
rect 19368 7046 19420 7098
rect 12520 6944 12572 6996
rect 14360 6944 14412 6996
rect 14820 6944 14872 6996
rect 19052 6987 19104 6996
rect 19052 6953 19061 6987
rect 19061 6953 19095 6987
rect 19095 6953 19104 6987
rect 19052 6944 19104 6953
rect 19788 6944 19840 6996
rect 20892 6987 20944 6996
rect 20892 6953 20901 6987
rect 20901 6953 20935 6987
rect 20935 6953 20944 6987
rect 20892 6944 20944 6953
rect 21168 6944 21220 6996
rect 22364 6944 22416 6996
rect 8104 6851 8156 6860
rect 8104 6817 8113 6851
rect 8113 6817 8147 6851
rect 8147 6817 8156 6851
rect 8104 6808 8156 6817
rect 9300 6876 9352 6928
rect 13348 6919 13400 6928
rect 10496 6808 10548 6860
rect 13348 6885 13357 6919
rect 13357 6885 13391 6919
rect 13391 6885 13400 6919
rect 13348 6876 13400 6885
rect 17764 6876 17816 6928
rect 21628 6919 21680 6928
rect 21628 6885 21637 6919
rect 21637 6885 21671 6919
rect 21671 6885 21680 6919
rect 21628 6876 21680 6885
rect 22548 6876 22600 6928
rect 23652 6876 23704 6928
rect 10680 6808 10732 6860
rect 10772 6808 10824 6860
rect 11692 6851 11744 6860
rect 11692 6817 11701 6851
rect 11701 6817 11735 6851
rect 11735 6817 11744 6851
rect 11692 6808 11744 6817
rect 12152 6851 12204 6860
rect 12152 6817 12161 6851
rect 12161 6817 12195 6851
rect 12195 6817 12204 6851
rect 12152 6808 12204 6817
rect 15740 6808 15792 6860
rect 16384 6851 16436 6860
rect 16384 6817 16393 6851
rect 16393 6817 16427 6851
rect 16427 6817 16436 6851
rect 16384 6808 16436 6817
rect 20432 6851 20484 6860
rect 20432 6817 20476 6851
rect 20476 6817 20484 6851
rect 20432 6808 20484 6817
rect 20616 6808 20668 6860
rect 24572 6808 24624 6860
rect 12336 6783 12388 6792
rect 12336 6749 12345 6783
rect 12345 6749 12379 6783
rect 12379 6749 12388 6783
rect 12336 6740 12388 6749
rect 13256 6783 13308 6792
rect 13256 6749 13265 6783
rect 13265 6749 13299 6783
rect 13299 6749 13308 6783
rect 13256 6740 13308 6749
rect 16016 6740 16068 6792
rect 16752 6740 16804 6792
rect 18040 6783 18092 6792
rect 18040 6749 18049 6783
rect 18049 6749 18083 6783
rect 18083 6749 18092 6783
rect 18040 6740 18092 6749
rect 18408 6783 18460 6792
rect 18408 6749 18417 6783
rect 18417 6749 18451 6783
rect 18451 6749 18460 6783
rect 18408 6740 18460 6749
rect 21352 6740 21404 6792
rect 23100 6740 23152 6792
rect 23560 6783 23612 6792
rect 23560 6749 23569 6783
rect 23569 6749 23603 6783
rect 23603 6749 23612 6783
rect 23560 6740 23612 6749
rect 10772 6647 10824 6656
rect 10772 6613 10781 6647
rect 10781 6613 10815 6647
rect 10815 6613 10824 6647
rect 10772 6604 10824 6613
rect 15096 6604 15148 6656
rect 15740 6647 15792 6656
rect 15740 6613 15749 6647
rect 15749 6613 15783 6647
rect 15783 6613 15792 6647
rect 15740 6604 15792 6613
rect 25860 6604 25912 6656
rect 5176 6502 5228 6554
rect 5240 6502 5292 6554
rect 5304 6502 5356 6554
rect 5368 6502 5420 6554
rect 14510 6502 14562 6554
rect 14574 6502 14626 6554
rect 14638 6502 14690 6554
rect 14702 6502 14754 6554
rect 23843 6502 23895 6554
rect 23907 6502 23959 6554
rect 23971 6502 24023 6554
rect 24035 6502 24087 6554
rect 6540 6400 6592 6452
rect 10404 6400 10456 6452
rect 10680 6400 10732 6452
rect 11416 6400 11468 6452
rect 8104 6307 8156 6316
rect 8104 6273 8113 6307
rect 8113 6273 8147 6307
rect 8147 6273 8156 6307
rect 8104 6264 8156 6273
rect 6172 6196 6224 6248
rect 9208 6239 9260 6248
rect 9208 6205 9217 6239
rect 9217 6205 9251 6239
rect 9251 6205 9260 6239
rect 9208 6196 9260 6205
rect 10864 6196 10916 6248
rect 7736 6128 7788 6180
rect 10404 6128 10456 6180
rect 13256 6400 13308 6452
rect 17764 6400 17816 6452
rect 19604 6443 19656 6452
rect 19604 6409 19613 6443
rect 19613 6409 19647 6443
rect 19647 6409 19656 6443
rect 19604 6400 19656 6409
rect 20984 6400 21036 6452
rect 23652 6400 23704 6452
rect 24572 6443 24624 6452
rect 24572 6409 24581 6443
rect 24581 6409 24615 6443
rect 24615 6409 24624 6443
rect 24572 6400 24624 6409
rect 15280 6332 15332 6384
rect 12060 6264 12112 6316
rect 13348 6264 13400 6316
rect 14268 6264 14320 6316
rect 16016 6307 16068 6316
rect 16016 6273 16025 6307
rect 16025 6273 16059 6307
rect 16059 6273 16068 6307
rect 16016 6264 16068 6273
rect 16292 6307 16344 6316
rect 16292 6273 16301 6307
rect 16301 6273 16335 6307
rect 16335 6273 16344 6307
rect 16292 6264 16344 6273
rect 13072 6128 13124 6180
rect 15188 6128 15240 6180
rect 8840 6103 8892 6112
rect 8840 6069 8849 6103
rect 8849 6069 8883 6103
rect 8883 6069 8892 6103
rect 8840 6060 8892 6069
rect 10680 6060 10732 6112
rect 11692 6060 11744 6112
rect 13256 6060 13308 6112
rect 16384 6128 16436 6180
rect 17672 6307 17724 6316
rect 17672 6273 17681 6307
rect 17681 6273 17715 6307
rect 17715 6273 17724 6307
rect 17672 6264 17724 6273
rect 18132 6307 18184 6316
rect 18132 6273 18141 6307
rect 18141 6273 18175 6307
rect 18175 6273 18184 6307
rect 18132 6264 18184 6273
rect 19604 6196 19656 6248
rect 19880 6196 19932 6248
rect 23192 6239 23244 6248
rect 20984 6128 21036 6180
rect 23192 6205 23201 6239
rect 23201 6205 23235 6239
rect 23235 6205 23244 6239
rect 23192 6196 23244 6205
rect 24756 6239 24808 6248
rect 24756 6205 24765 6239
rect 24765 6205 24799 6239
rect 24799 6205 24808 6239
rect 24756 6196 24808 6205
rect 20800 6060 20852 6112
rect 21904 6060 21956 6112
rect 22272 6103 22324 6112
rect 22272 6069 22281 6103
rect 22281 6069 22315 6103
rect 22315 6069 22324 6103
rect 22272 6060 22324 6069
rect 23744 6060 23796 6112
rect 9843 5958 9895 6010
rect 9907 5958 9959 6010
rect 9971 5958 10023 6010
rect 10035 5958 10087 6010
rect 19176 5958 19228 6010
rect 19240 5958 19292 6010
rect 19304 5958 19356 6010
rect 19368 5958 19420 6010
rect 10496 5899 10548 5908
rect 10496 5865 10505 5899
rect 10505 5865 10539 5899
rect 10539 5865 10548 5899
rect 10496 5856 10548 5865
rect 10864 5899 10916 5908
rect 10864 5865 10873 5899
rect 10873 5865 10907 5899
rect 10907 5865 10916 5899
rect 10864 5856 10916 5865
rect 11876 5856 11928 5908
rect 12060 5856 12112 5908
rect 14268 5899 14320 5908
rect 14268 5865 14277 5899
rect 14277 5865 14311 5899
rect 14311 5865 14320 5899
rect 14268 5856 14320 5865
rect 16016 5899 16068 5908
rect 16016 5865 16025 5899
rect 16025 5865 16059 5899
rect 16059 5865 16068 5899
rect 16016 5856 16068 5865
rect 17672 5899 17724 5908
rect 17672 5865 17681 5899
rect 17681 5865 17715 5899
rect 17715 5865 17724 5899
rect 17672 5856 17724 5865
rect 18040 5899 18092 5908
rect 18040 5865 18049 5899
rect 18049 5865 18083 5899
rect 18083 5865 18092 5899
rect 18040 5856 18092 5865
rect 18776 5856 18828 5908
rect 21628 5856 21680 5908
rect 22456 5856 22508 5908
rect 9208 5788 9260 5840
rect 10036 5788 10088 5840
rect 10772 5788 10824 5840
rect 11416 5831 11468 5840
rect 11416 5797 11419 5831
rect 11419 5797 11453 5831
rect 11453 5797 11468 5831
rect 11416 5788 11468 5797
rect 12152 5788 12204 5840
rect 13256 5788 13308 5840
rect 15188 5831 15240 5840
rect 15188 5797 15191 5831
rect 15191 5797 15225 5831
rect 15225 5797 15240 5831
rect 15188 5788 15240 5797
rect 16752 5831 16804 5840
rect 16752 5797 16761 5831
rect 16761 5797 16795 5831
rect 16795 5797 16804 5831
rect 16752 5788 16804 5797
rect 6448 5720 6500 5772
rect 7644 5720 7696 5772
rect 8196 5763 8248 5772
rect 8196 5729 8205 5763
rect 8205 5729 8239 5763
rect 8239 5729 8248 5763
rect 8196 5720 8248 5729
rect 11048 5763 11100 5772
rect 11048 5729 11057 5763
rect 11057 5729 11091 5763
rect 11091 5729 11100 5763
rect 11048 5720 11100 5729
rect 14360 5720 14412 5772
rect 14820 5763 14872 5772
rect 14820 5729 14829 5763
rect 14829 5729 14863 5763
rect 14863 5729 14872 5763
rect 14820 5720 14872 5729
rect 17856 5720 17908 5772
rect 19604 5788 19656 5840
rect 19880 5831 19932 5840
rect 19880 5797 19889 5831
rect 19889 5797 19923 5831
rect 19923 5797 19932 5831
rect 19880 5788 19932 5797
rect 20340 5788 20392 5840
rect 20616 5788 20668 5840
rect 21352 5788 21404 5840
rect 21904 5788 21956 5840
rect 23192 5831 23244 5840
rect 23192 5797 23201 5831
rect 23201 5797 23235 5831
rect 23235 5797 23244 5831
rect 23192 5788 23244 5797
rect 24480 5788 24532 5840
rect 18592 5763 18644 5772
rect 18592 5729 18601 5763
rect 18601 5729 18635 5763
rect 18635 5729 18644 5763
rect 18592 5720 18644 5729
rect 19972 5720 20024 5772
rect 20708 5720 20760 5772
rect 8932 5652 8984 5704
rect 9300 5652 9352 5704
rect 9760 5652 9812 5704
rect 13164 5652 13216 5704
rect 13348 5695 13400 5704
rect 13348 5661 13357 5695
rect 13357 5661 13391 5695
rect 13391 5661 13400 5695
rect 13348 5652 13400 5661
rect 16660 5695 16712 5704
rect 16660 5661 16669 5695
rect 16669 5661 16703 5695
rect 16703 5661 16712 5695
rect 16660 5652 16712 5661
rect 18684 5695 18736 5704
rect 7736 5584 7788 5636
rect 16292 5584 16344 5636
rect 18684 5661 18693 5695
rect 18693 5661 18727 5695
rect 18727 5661 18736 5695
rect 18684 5652 18736 5661
rect 20248 5652 20300 5704
rect 20984 5720 21036 5772
rect 23100 5720 23152 5772
rect 22088 5652 22140 5704
rect 23008 5652 23060 5704
rect 24296 5652 24348 5704
rect 24388 5627 24440 5636
rect 24388 5593 24397 5627
rect 24397 5593 24431 5627
rect 24431 5593 24440 5627
rect 24388 5584 24440 5593
rect 12244 5516 12296 5568
rect 15556 5516 15608 5568
rect 22916 5559 22968 5568
rect 22916 5525 22925 5559
rect 22925 5525 22959 5559
rect 22959 5525 22968 5559
rect 22916 5516 22968 5525
rect 5176 5414 5228 5466
rect 5240 5414 5292 5466
rect 5304 5414 5356 5466
rect 5368 5414 5420 5466
rect 14510 5414 14562 5466
rect 14574 5414 14626 5466
rect 14638 5414 14690 5466
rect 14702 5414 14754 5466
rect 23843 5414 23895 5466
rect 23907 5414 23959 5466
rect 23971 5414 24023 5466
rect 24035 5414 24087 5466
rect 6448 5312 6500 5364
rect 7644 5312 7696 5364
rect 8840 5355 8892 5364
rect 8840 5321 8849 5355
rect 8849 5321 8883 5355
rect 8883 5321 8892 5355
rect 8840 5312 8892 5321
rect 10036 5355 10088 5364
rect 10036 5321 10045 5355
rect 10045 5321 10079 5355
rect 10079 5321 10088 5355
rect 10036 5312 10088 5321
rect 11048 5312 11100 5364
rect 14360 5312 14412 5364
rect 16752 5312 16804 5364
rect 17856 5355 17908 5364
rect 17856 5321 17865 5355
rect 17865 5321 17899 5355
rect 17899 5321 17908 5355
rect 17856 5312 17908 5321
rect 18592 5312 18644 5364
rect 20248 5312 20300 5364
rect 20800 5312 20852 5364
rect 24296 5312 24348 5364
rect 24480 5355 24532 5364
rect 24480 5321 24489 5355
rect 24489 5321 24523 5355
rect 24523 5321 24532 5355
rect 24480 5312 24532 5321
rect 9300 5244 9352 5296
rect 17028 5244 17080 5296
rect 19972 5244 20024 5296
rect 6540 5176 6592 5228
rect 9760 5219 9812 5228
rect 9760 5185 9769 5219
rect 9769 5185 9803 5219
rect 9803 5185 9812 5219
rect 9760 5176 9812 5185
rect 10312 5176 10364 5228
rect 12336 5176 12388 5228
rect 15188 5176 15240 5228
rect 8104 5151 8156 5160
rect 8104 5117 8113 5151
rect 8113 5117 8147 5151
rect 8147 5117 8156 5151
rect 8104 5108 8156 5117
rect 11784 5108 11836 5160
rect 15280 5151 15332 5160
rect 15280 5117 15289 5151
rect 15289 5117 15323 5151
rect 15323 5117 15332 5151
rect 15280 5108 15332 5117
rect 8196 5083 8248 5092
rect 8196 5049 8205 5083
rect 8205 5049 8239 5083
rect 8239 5049 8248 5083
rect 8196 5040 8248 5049
rect 8472 5015 8524 5024
rect 8472 4981 8481 5015
rect 8481 4981 8515 5015
rect 8515 4981 8524 5015
rect 8472 4972 8524 4981
rect 8840 4972 8892 5024
rect 11968 5040 12020 5092
rect 11324 4972 11376 5024
rect 13072 5040 13124 5092
rect 13256 5040 13308 5092
rect 14636 5083 14688 5092
rect 14636 5049 14645 5083
rect 14645 5049 14679 5083
rect 14679 5049 14688 5083
rect 14636 5040 14688 5049
rect 13532 4972 13584 5024
rect 13716 5015 13768 5024
rect 13716 4981 13725 5015
rect 13725 4981 13759 5015
rect 13759 4981 13768 5015
rect 13716 4972 13768 4981
rect 16108 4972 16160 5024
rect 16660 5176 16712 5228
rect 18776 5176 18828 5228
rect 20248 5176 20300 5228
rect 23376 5176 23428 5228
rect 24296 5176 24348 5228
rect 19972 5108 20024 5160
rect 25032 5151 25084 5160
rect 25032 5117 25041 5151
rect 25041 5117 25075 5151
rect 25075 5117 25084 5151
rect 25032 5108 25084 5117
rect 16936 5040 16988 5092
rect 18776 5040 18828 5092
rect 20800 5040 20852 5092
rect 24296 5040 24348 5092
rect 21536 5015 21588 5024
rect 21536 4981 21545 5015
rect 21545 4981 21579 5015
rect 21579 4981 21588 5015
rect 21536 4972 21588 4981
rect 23008 5015 23060 5024
rect 23008 4981 23017 5015
rect 23017 4981 23051 5015
rect 23051 4981 23060 5015
rect 23008 4972 23060 4981
rect 25216 5015 25268 5024
rect 25216 4981 25225 5015
rect 25225 4981 25259 5015
rect 25259 4981 25268 5015
rect 25216 4972 25268 4981
rect 9843 4870 9895 4922
rect 9907 4870 9959 4922
rect 9971 4870 10023 4922
rect 10035 4870 10087 4922
rect 19176 4870 19228 4922
rect 19240 4870 19292 4922
rect 19304 4870 19356 4922
rect 19368 4870 19420 4922
rect 5804 4768 5856 4820
rect 10312 4811 10364 4820
rect 10312 4777 10321 4811
rect 10321 4777 10355 4811
rect 10355 4777 10364 4811
rect 10312 4768 10364 4777
rect 11784 4811 11836 4820
rect 11784 4777 11793 4811
rect 11793 4777 11827 4811
rect 11827 4777 11836 4811
rect 11784 4768 11836 4777
rect 12336 4768 12388 4820
rect 13164 4768 13216 4820
rect 18592 4768 18644 4820
rect 21352 4811 21404 4820
rect 21352 4777 21361 4811
rect 21361 4777 21395 4811
rect 21395 4777 21404 4811
rect 21352 4768 21404 4777
rect 22088 4811 22140 4820
rect 22088 4777 22097 4811
rect 22097 4777 22131 4811
rect 22131 4777 22140 4811
rect 22088 4768 22140 4777
rect 23376 4811 23428 4820
rect 23376 4777 23385 4811
rect 23385 4777 23419 4811
rect 23419 4777 23428 4811
rect 23376 4768 23428 4777
rect 11324 4700 11376 4752
rect 13440 4700 13492 4752
rect 14636 4700 14688 4752
rect 16936 4700 16988 4752
rect 18776 4700 18828 4752
rect 20800 4743 20852 4752
rect 20800 4709 20803 4743
rect 20803 4709 20837 4743
rect 20837 4709 20852 4743
rect 20800 4700 20852 4709
rect 23652 4743 23704 4752
rect 23652 4709 23661 4743
rect 23661 4709 23695 4743
rect 23695 4709 23704 4743
rect 23652 4700 23704 4709
rect 4792 4632 4844 4684
rect 5712 4632 5764 4684
rect 8196 4675 8248 4684
rect 8196 4641 8205 4675
rect 8205 4641 8239 4675
rect 8239 4641 8248 4675
rect 8196 4632 8248 4641
rect 9484 4675 9536 4684
rect 9484 4641 9493 4675
rect 9493 4641 9527 4675
rect 9527 4641 9536 4675
rect 9484 4632 9536 4641
rect 10496 4675 10548 4684
rect 10496 4641 10505 4675
rect 10505 4641 10539 4675
rect 10539 4641 10548 4675
rect 10496 4632 10548 4641
rect 15096 4675 15148 4684
rect 15096 4641 15105 4675
rect 15105 4641 15139 4675
rect 15139 4641 15148 4675
rect 15096 4632 15148 4641
rect 16200 4675 16252 4684
rect 16200 4641 16209 4675
rect 16209 4641 16243 4675
rect 16243 4641 16252 4675
rect 16200 4632 16252 4641
rect 18684 4632 18736 4684
rect 20248 4632 20300 4684
rect 22180 4675 22232 4684
rect 22180 4641 22189 4675
rect 22189 4641 22223 4675
rect 22223 4641 22232 4675
rect 22180 4632 22232 4641
rect 6540 4607 6592 4616
rect 6540 4573 6549 4607
rect 6549 4573 6583 4607
rect 6583 4573 6592 4607
rect 6540 4564 6592 4573
rect 9116 4564 9168 4616
rect 13256 4607 13308 4616
rect 13256 4573 13265 4607
rect 13265 4573 13299 4607
rect 13299 4573 13308 4607
rect 13256 4564 13308 4573
rect 13900 4607 13952 4616
rect 13900 4573 13909 4607
rect 13909 4573 13943 4607
rect 13943 4573 13952 4607
rect 13900 4564 13952 4573
rect 23192 4564 23244 4616
rect 24296 4564 24348 4616
rect 4976 4496 5028 4548
rect 21720 4496 21772 4548
rect 11416 4471 11468 4480
rect 11416 4437 11425 4471
rect 11425 4437 11459 4471
rect 11459 4437 11468 4471
rect 11416 4428 11468 4437
rect 15280 4471 15332 4480
rect 15280 4437 15289 4471
rect 15289 4437 15323 4471
rect 15323 4437 15332 4471
rect 15280 4428 15332 4437
rect 17120 4471 17172 4480
rect 17120 4437 17129 4471
rect 17129 4437 17163 4471
rect 17163 4437 17172 4471
rect 17120 4428 17172 4437
rect 17488 4428 17540 4480
rect 19512 4471 19564 4480
rect 19512 4437 19521 4471
rect 19521 4437 19555 4471
rect 19555 4437 19564 4471
rect 19512 4428 19564 4437
rect 5176 4326 5228 4378
rect 5240 4326 5292 4378
rect 5304 4326 5356 4378
rect 5368 4326 5420 4378
rect 14510 4326 14562 4378
rect 14574 4326 14626 4378
rect 14638 4326 14690 4378
rect 14702 4326 14754 4378
rect 23843 4326 23895 4378
rect 23907 4326 23959 4378
rect 23971 4326 24023 4378
rect 24035 4326 24087 4378
rect 11324 4267 11376 4276
rect 11324 4233 11333 4267
rect 11333 4233 11367 4267
rect 11367 4233 11376 4267
rect 11324 4224 11376 4233
rect 13440 4267 13492 4276
rect 13440 4233 13449 4267
rect 13449 4233 13483 4267
rect 13483 4233 13492 4267
rect 13440 4224 13492 4233
rect 16936 4224 16988 4276
rect 18776 4224 18828 4276
rect 20248 4224 20300 4276
rect 21352 4267 21404 4276
rect 21352 4233 21361 4267
rect 21361 4233 21395 4267
rect 21395 4233 21404 4267
rect 21352 4224 21404 4233
rect 23652 4224 23704 4276
rect 8196 4156 8248 4208
rect 10312 4156 10364 4208
rect 18684 4156 18736 4208
rect 3596 3884 3648 3936
rect 5528 4020 5580 4072
rect 7552 4020 7604 4072
rect 9116 4063 9168 4072
rect 9116 4029 9125 4063
rect 9125 4029 9159 4063
rect 9159 4029 9168 4063
rect 9116 4020 9168 4029
rect 5896 3952 5948 4004
rect 12428 4131 12480 4140
rect 12428 4097 12437 4131
rect 12437 4097 12471 4131
rect 12471 4097 12480 4131
rect 12428 4088 12480 4097
rect 13348 4088 13400 4140
rect 14176 4088 14228 4140
rect 14268 4131 14320 4140
rect 14268 4097 14277 4131
rect 14277 4097 14311 4131
rect 14311 4097 14320 4131
rect 15556 4131 15608 4140
rect 14268 4088 14320 4097
rect 15556 4097 15565 4131
rect 15565 4097 15599 4131
rect 15599 4097 15608 4131
rect 15556 4088 15608 4097
rect 16200 4088 16252 4140
rect 20800 4156 20852 4208
rect 21444 4156 21496 4208
rect 19696 4088 19748 4140
rect 21904 4088 21956 4140
rect 23192 4156 23244 4208
rect 23376 4088 23428 4140
rect 23468 4088 23520 4140
rect 24756 4063 24808 4072
rect 24756 4029 24765 4063
rect 24765 4029 24799 4063
rect 24799 4029 24808 4063
rect 24756 4020 24808 4029
rect 10680 3952 10732 4004
rect 12152 3995 12204 4004
rect 4148 3884 4200 3936
rect 4608 3884 4660 3936
rect 4792 3927 4844 3936
rect 4792 3893 4801 3927
rect 4801 3893 4835 3927
rect 4835 3893 4844 3927
rect 4792 3884 4844 3893
rect 5620 3884 5672 3936
rect 5712 3927 5764 3936
rect 5712 3893 5721 3927
rect 5721 3893 5755 3927
rect 5755 3893 5764 3927
rect 6724 3927 6776 3936
rect 5712 3884 5764 3893
rect 6724 3893 6733 3927
rect 6733 3893 6767 3927
rect 6767 3893 6776 3927
rect 6724 3884 6776 3893
rect 9024 3927 9076 3936
rect 9024 3893 9033 3927
rect 9033 3893 9067 3927
rect 9067 3893 9076 3927
rect 9024 3884 9076 3893
rect 10312 3884 10364 3936
rect 12152 3961 12161 3995
rect 12161 3961 12195 3995
rect 12195 3961 12204 3995
rect 12152 3952 12204 3961
rect 13532 3884 13584 3936
rect 14820 3884 14872 3936
rect 17488 3952 17540 4004
rect 19052 3952 19104 4004
rect 19512 3884 19564 3936
rect 21352 3952 21404 4004
rect 22456 3952 22508 4004
rect 23376 3995 23428 4004
rect 23376 3961 23385 3995
rect 23385 3961 23419 3995
rect 23419 3961 23428 3995
rect 23376 3952 23428 3961
rect 20156 3884 20208 3936
rect 23192 3884 23244 3936
rect 24940 3927 24992 3936
rect 24940 3893 24949 3927
rect 24949 3893 24983 3927
rect 24983 3893 24992 3927
rect 24940 3884 24992 3893
rect 9843 3782 9895 3834
rect 9907 3782 9959 3834
rect 9971 3782 10023 3834
rect 10035 3782 10087 3834
rect 19176 3782 19228 3834
rect 19240 3782 19292 3834
rect 19304 3782 19356 3834
rect 19368 3782 19420 3834
rect 4056 3680 4108 3732
rect 6080 3680 6132 3732
rect 8380 3680 8432 3732
rect 10588 3680 10640 3732
rect 12428 3723 12480 3732
rect 12428 3689 12437 3723
rect 12437 3689 12471 3723
rect 12471 3689 12480 3723
rect 12428 3680 12480 3689
rect 14176 3723 14228 3732
rect 14176 3689 14185 3723
rect 14185 3689 14219 3723
rect 14219 3689 14228 3723
rect 14176 3680 14228 3689
rect 15096 3680 15148 3732
rect 16292 3680 16344 3732
rect 19972 3680 20024 3732
rect 20432 3680 20484 3732
rect 21444 3723 21496 3732
rect 9208 3612 9260 3664
rect 10128 3612 10180 3664
rect 11324 3612 11376 3664
rect 15556 3612 15608 3664
rect 17120 3612 17172 3664
rect 20524 3655 20576 3664
rect 20524 3621 20533 3655
rect 20533 3621 20567 3655
rect 20567 3621 20576 3655
rect 20524 3612 20576 3621
rect 21444 3689 21453 3723
rect 21453 3689 21487 3723
rect 21487 3689 21496 3723
rect 21444 3680 21496 3689
rect 23560 3680 23612 3732
rect 22180 3655 22232 3664
rect 22180 3621 22189 3655
rect 22189 3621 22223 3655
rect 22223 3621 22232 3655
rect 22180 3612 22232 3621
rect 3964 3587 4016 3596
rect 3964 3553 3982 3587
rect 3982 3553 4016 3587
rect 3964 3544 4016 3553
rect 5068 3544 5120 3596
rect 5988 3587 6040 3596
rect 5988 3553 6006 3587
rect 6006 3553 6040 3587
rect 5988 3544 6040 3553
rect 8288 3544 8340 3596
rect 13532 3587 13584 3596
rect 13532 3553 13541 3587
rect 13541 3553 13575 3587
rect 13575 3553 13584 3587
rect 13532 3544 13584 3553
rect 14912 3587 14964 3596
rect 14912 3553 14930 3587
rect 14930 3553 14964 3587
rect 14912 3544 14964 3553
rect 18960 3587 19012 3596
rect 18960 3553 18969 3587
rect 18969 3553 19003 3587
rect 19003 3553 19012 3587
rect 18960 3544 19012 3553
rect 6908 3519 6960 3528
rect 6908 3485 6917 3519
rect 6917 3485 6951 3519
rect 6951 3485 6960 3519
rect 6908 3476 6960 3485
rect 9300 3476 9352 3528
rect 10220 3519 10272 3528
rect 10220 3485 10229 3519
rect 10229 3485 10263 3519
rect 10263 3485 10272 3519
rect 10220 3476 10272 3485
rect 11600 3476 11652 3528
rect 12060 3476 12112 3528
rect 13900 3476 13952 3528
rect 16200 3519 16252 3528
rect 16200 3485 16209 3519
rect 16209 3485 16243 3519
rect 16243 3485 16252 3519
rect 16200 3476 16252 3485
rect 17580 3476 17632 3528
rect 16292 3408 16344 3460
rect 18132 3476 18184 3528
rect 22088 3519 22140 3528
rect 18040 3451 18092 3460
rect 18040 3417 18049 3451
rect 18049 3417 18083 3451
rect 18083 3417 18092 3451
rect 18040 3408 18092 3417
rect 19052 3408 19104 3460
rect 22088 3485 22097 3519
rect 22097 3485 22131 3519
rect 22131 3485 22140 3519
rect 22088 3476 22140 3485
rect 22364 3519 22416 3528
rect 22364 3485 22373 3519
rect 22373 3485 22407 3519
rect 22407 3485 22416 3519
rect 22364 3476 22416 3485
rect 22456 3476 22508 3528
rect 23652 3519 23704 3528
rect 23652 3485 23661 3519
rect 23661 3485 23695 3519
rect 23695 3485 23704 3519
rect 23652 3476 23704 3485
rect 4884 3340 4936 3392
rect 9392 3340 9444 3392
rect 13624 3383 13676 3392
rect 13624 3349 13633 3383
rect 13633 3349 13667 3383
rect 13667 3349 13676 3383
rect 13624 3340 13676 3349
rect 16016 3340 16068 3392
rect 17672 3340 17724 3392
rect 18592 3340 18644 3392
rect 23192 3383 23244 3392
rect 23192 3349 23201 3383
rect 23201 3349 23235 3383
rect 23235 3349 23244 3383
rect 23192 3340 23244 3349
rect 5176 3238 5228 3290
rect 5240 3238 5292 3290
rect 5304 3238 5356 3290
rect 5368 3238 5420 3290
rect 14510 3238 14562 3290
rect 14574 3238 14626 3290
rect 14638 3238 14690 3290
rect 14702 3238 14754 3290
rect 23843 3238 23895 3290
rect 23907 3238 23959 3290
rect 23971 3238 24023 3290
rect 24035 3238 24087 3290
rect 2768 3179 2820 3188
rect 2768 3145 2777 3179
rect 2777 3145 2811 3179
rect 2811 3145 2820 3179
rect 2768 3136 2820 3145
rect 3412 3136 3464 3188
rect 3780 3179 3832 3188
rect 3780 3145 3789 3179
rect 3789 3145 3823 3179
rect 3823 3145 3832 3179
rect 3780 3136 3832 3145
rect 3964 3136 4016 3188
rect 4424 3136 4476 3188
rect 5068 3179 5120 3188
rect 5068 3145 5077 3179
rect 5077 3145 5111 3179
rect 5111 3145 5120 3179
rect 5068 3136 5120 3145
rect 5804 3179 5856 3188
rect 5804 3145 5813 3179
rect 5813 3145 5847 3179
rect 5847 3145 5856 3179
rect 5804 3136 5856 3145
rect 5988 3136 6040 3188
rect 9300 3136 9352 3188
rect 10128 3179 10180 3188
rect 10128 3145 10137 3179
rect 10137 3145 10171 3179
rect 10171 3145 10180 3179
rect 10128 3136 10180 3145
rect 10404 3136 10456 3188
rect 12244 3136 12296 3188
rect 12428 3136 12480 3188
rect 13164 3179 13216 3188
rect 13164 3145 13173 3179
rect 13173 3145 13207 3179
rect 13207 3145 13216 3179
rect 13164 3136 13216 3145
rect 13624 3179 13676 3188
rect 13624 3145 13633 3179
rect 13633 3145 13667 3179
rect 13667 3145 13676 3179
rect 13624 3136 13676 3145
rect 15556 3136 15608 3188
rect 2768 2932 2820 2984
rect 3780 2932 3832 2984
rect 4240 2975 4292 2984
rect 4240 2941 4284 2975
rect 4284 2941 4292 2975
rect 4240 2932 4292 2941
rect 8840 3043 8892 3052
rect 7184 2975 7236 2984
rect 7184 2941 7193 2975
rect 7193 2941 7227 2975
rect 7227 2941 7236 2975
rect 8840 3009 8849 3043
rect 8849 3009 8883 3043
rect 8883 3009 8892 3043
rect 8840 3000 8892 3009
rect 9208 3000 9260 3052
rect 12060 3043 12112 3052
rect 12060 3009 12069 3043
rect 12069 3009 12103 3043
rect 12103 3009 12112 3043
rect 12060 3000 12112 3009
rect 12336 3043 12388 3052
rect 12336 3009 12345 3043
rect 12345 3009 12379 3043
rect 12379 3009 12388 3043
rect 12336 3000 12388 3009
rect 7184 2932 7236 2941
rect 9116 2932 9168 2984
rect 5804 2864 5856 2916
rect 10404 2864 10456 2916
rect 10496 2907 10548 2916
rect 10496 2873 10505 2907
rect 10505 2873 10539 2907
rect 10539 2873 10548 2907
rect 10496 2864 10548 2873
rect 12428 2864 12480 2916
rect 3228 2796 3280 2848
rect 7644 2796 7696 2848
rect 8288 2796 8340 2848
rect 11324 2839 11376 2848
rect 11324 2805 11333 2839
rect 11333 2805 11367 2839
rect 11367 2805 11376 2839
rect 11324 2796 11376 2805
rect 13808 3043 13860 3052
rect 13808 3009 13817 3043
rect 13817 3009 13851 3043
rect 13851 3009 13860 3043
rect 13808 3000 13860 3009
rect 14268 3043 14320 3052
rect 14268 3009 14277 3043
rect 14277 3009 14311 3043
rect 14311 3009 14320 3043
rect 14268 3000 14320 3009
rect 17120 3136 17172 3188
rect 20432 3136 20484 3188
rect 22088 3068 22140 3120
rect 17672 3043 17724 3052
rect 17672 3009 17681 3043
rect 17681 3009 17715 3043
rect 17715 3009 17724 3043
rect 17672 3000 17724 3009
rect 18040 3043 18092 3052
rect 18040 3009 18049 3043
rect 18049 3009 18083 3043
rect 18083 3009 18092 3043
rect 18040 3000 18092 3009
rect 19696 3043 19748 3052
rect 19696 3009 19705 3043
rect 19705 3009 19739 3043
rect 19739 3009 19748 3043
rect 19696 3000 19748 3009
rect 22456 3000 22508 3052
rect 23652 3136 23704 3188
rect 24940 3179 24992 3188
rect 24940 3145 24949 3179
rect 24949 3145 24983 3179
rect 24983 3145 24992 3179
rect 24940 3136 24992 3145
rect 23468 3068 23520 3120
rect 23560 2932 23612 2984
rect 24204 2932 24256 2984
rect 25216 2932 25268 2984
rect 14912 2907 14964 2916
rect 14912 2873 14921 2907
rect 14921 2873 14955 2907
rect 14955 2873 14964 2907
rect 14912 2864 14964 2873
rect 16568 2864 16620 2916
rect 18500 2864 18552 2916
rect 19696 2864 19748 2916
rect 20064 2864 20116 2916
rect 21260 2864 21312 2916
rect 23008 2864 23060 2916
rect 22180 2796 22232 2848
rect 22916 2796 22968 2848
rect 9843 2694 9895 2746
rect 9907 2694 9959 2746
rect 9971 2694 10023 2746
rect 10035 2694 10087 2746
rect 19176 2694 19228 2746
rect 19240 2694 19292 2746
rect 19304 2694 19356 2746
rect 19368 2694 19420 2746
rect 1664 2592 1716 2644
rect 4516 2592 4568 2644
rect 7276 2592 7328 2644
rect 7736 2635 7788 2644
rect 7736 2601 7745 2635
rect 7745 2601 7779 2635
rect 7779 2601 7788 2635
rect 7736 2592 7788 2601
rect 8656 2592 8708 2644
rect 10220 2592 10272 2644
rect 3044 2456 3096 2508
rect 4332 2499 4384 2508
rect 4332 2465 4376 2499
rect 4376 2465 4384 2499
rect 4332 2456 4384 2465
rect 8748 2456 8800 2508
rect 11324 2592 11376 2644
rect 13532 2592 13584 2644
rect 14820 2635 14872 2644
rect 14820 2601 14829 2635
rect 14829 2601 14863 2635
rect 14863 2601 14872 2635
rect 14820 2592 14872 2601
rect 5344 2431 5396 2440
rect 5344 2397 5353 2431
rect 5353 2397 5387 2431
rect 5387 2397 5396 2431
rect 5344 2388 5396 2397
rect 2124 2252 2176 2304
rect 2860 2252 2912 2304
rect 3044 2295 3096 2304
rect 3044 2261 3053 2295
rect 3053 2261 3087 2295
rect 3087 2261 3096 2295
rect 3044 2252 3096 2261
rect 8748 2295 8800 2304
rect 8748 2261 8757 2295
rect 8757 2261 8791 2295
rect 8791 2261 8800 2295
rect 8748 2252 8800 2261
rect 13808 2499 13860 2508
rect 13808 2465 13817 2499
rect 13817 2465 13851 2499
rect 13851 2465 13860 2499
rect 16292 2592 16344 2644
rect 23468 2592 23520 2644
rect 18684 2524 18736 2576
rect 19696 2524 19748 2576
rect 23008 2524 23060 2576
rect 13808 2456 13860 2465
rect 16660 2499 16712 2508
rect 16660 2465 16669 2499
rect 16669 2465 16703 2499
rect 16703 2465 16712 2499
rect 16660 2456 16712 2465
rect 20340 2456 20392 2508
rect 22272 2499 22324 2508
rect 22272 2465 22281 2499
rect 22281 2465 22315 2499
rect 22315 2465 22324 2499
rect 25216 2592 25268 2644
rect 22272 2456 22324 2465
rect 24388 2456 24440 2508
rect 10496 2431 10548 2440
rect 10496 2397 10505 2431
rect 10505 2397 10539 2431
rect 10539 2397 10548 2431
rect 10496 2388 10548 2397
rect 11508 2431 11560 2440
rect 11508 2397 11517 2431
rect 11517 2397 11551 2431
rect 11551 2397 11560 2431
rect 11508 2388 11560 2397
rect 12336 2388 12388 2440
rect 17488 2320 17540 2372
rect 19052 2363 19104 2372
rect 19052 2329 19061 2363
rect 19061 2329 19095 2363
rect 19095 2329 19104 2363
rect 19052 2320 19104 2329
rect 10312 2252 10364 2304
rect 13992 2295 14044 2304
rect 13992 2261 14001 2295
rect 14001 2261 14035 2295
rect 14035 2261 14044 2295
rect 13992 2252 14044 2261
rect 17580 2295 17632 2304
rect 17580 2261 17589 2295
rect 17589 2261 17623 2295
rect 17623 2261 17632 2295
rect 17580 2252 17632 2261
rect 18960 2252 19012 2304
rect 19420 2295 19472 2304
rect 19420 2261 19429 2295
rect 19429 2261 19463 2295
rect 19463 2261 19472 2295
rect 19420 2252 19472 2261
rect 20064 2295 20116 2304
rect 20064 2261 20073 2295
rect 20073 2261 20107 2295
rect 20107 2261 20116 2295
rect 20064 2252 20116 2261
rect 22456 2295 22508 2304
rect 22456 2261 22465 2295
rect 22465 2261 22499 2295
rect 22499 2261 22508 2295
rect 22456 2252 22508 2261
rect 5176 2150 5228 2202
rect 5240 2150 5292 2202
rect 5304 2150 5356 2202
rect 5368 2150 5420 2202
rect 14510 2150 14562 2202
rect 14574 2150 14626 2202
rect 14638 2150 14690 2202
rect 14702 2150 14754 2202
rect 23843 2150 23895 2202
rect 23907 2150 23959 2202
rect 23971 2150 24023 2202
rect 24035 2150 24087 2202
<< metal2 >>
rect 1294 27520 1350 28000
rect 4790 27520 4846 28000
rect 8286 27520 8342 28000
rect 11782 27520 11838 28000
rect 15278 27520 15334 28000
rect 18774 27520 18830 28000
rect 22270 27520 22326 28000
rect 25766 27520 25822 28000
rect 1308 26194 1336 27520
rect 4804 27470 4832 27520
rect 3688 27464 3740 27470
rect 3688 27406 3740 27412
rect 4792 27464 4844 27470
rect 4792 27406 4844 27412
rect 1032 26166 1336 26194
rect 1032 14385 1060 26166
rect 1018 14376 1074 14385
rect 1018 14311 1074 14320
rect 3700 11257 3728 27406
rect 5150 25052 5446 25072
rect 5206 25050 5230 25052
rect 5286 25050 5310 25052
rect 5366 25050 5390 25052
rect 5228 24998 5230 25050
rect 5292 24998 5304 25050
rect 5366 24998 5368 25050
rect 5206 24996 5230 24998
rect 5286 24996 5310 24998
rect 5366 24996 5390 24998
rect 5150 24976 5446 24996
rect 5150 23964 5446 23984
rect 5206 23962 5230 23964
rect 5286 23962 5310 23964
rect 5366 23962 5390 23964
rect 5228 23910 5230 23962
rect 5292 23910 5304 23962
rect 5366 23910 5368 23962
rect 5206 23908 5230 23910
rect 5286 23908 5310 23910
rect 5366 23908 5390 23910
rect 5150 23888 5446 23908
rect 5150 22876 5446 22896
rect 5206 22874 5230 22876
rect 5286 22874 5310 22876
rect 5366 22874 5390 22876
rect 5228 22822 5230 22874
rect 5292 22822 5304 22874
rect 5366 22822 5368 22874
rect 5206 22820 5230 22822
rect 5286 22820 5310 22822
rect 5366 22820 5390 22822
rect 5150 22800 5446 22820
rect 5150 21788 5446 21808
rect 5206 21786 5230 21788
rect 5286 21786 5310 21788
rect 5366 21786 5390 21788
rect 5228 21734 5230 21786
rect 5292 21734 5304 21786
rect 5366 21734 5368 21786
rect 5206 21732 5230 21734
rect 5286 21732 5310 21734
rect 5366 21732 5390 21734
rect 5150 21712 5446 21732
rect 5150 20700 5446 20720
rect 5206 20698 5230 20700
rect 5286 20698 5310 20700
rect 5366 20698 5390 20700
rect 5228 20646 5230 20698
rect 5292 20646 5304 20698
rect 5366 20646 5368 20698
rect 5206 20644 5230 20646
rect 5286 20644 5310 20646
rect 5366 20644 5390 20646
rect 5150 20624 5446 20644
rect 5150 19612 5446 19632
rect 5206 19610 5230 19612
rect 5286 19610 5310 19612
rect 5366 19610 5390 19612
rect 5228 19558 5230 19610
rect 5292 19558 5304 19610
rect 5366 19558 5368 19610
rect 5206 19556 5230 19558
rect 5286 19556 5310 19558
rect 5366 19556 5390 19558
rect 5150 19536 5446 19556
rect 5150 18524 5446 18544
rect 5206 18522 5230 18524
rect 5286 18522 5310 18524
rect 5366 18522 5390 18524
rect 5228 18470 5230 18522
rect 5292 18470 5304 18522
rect 5366 18470 5368 18522
rect 5206 18468 5230 18470
rect 5286 18468 5310 18470
rect 5366 18468 5390 18470
rect 5150 18448 5446 18468
rect 8300 18057 8328 27520
rect 9817 25596 10113 25616
rect 9873 25594 9897 25596
rect 9953 25594 9977 25596
rect 10033 25594 10057 25596
rect 9895 25542 9897 25594
rect 9959 25542 9971 25594
rect 10033 25542 10035 25594
rect 9873 25540 9897 25542
rect 9953 25540 9977 25542
rect 10033 25540 10057 25542
rect 9817 25520 10113 25540
rect 9817 24508 10113 24528
rect 9873 24506 9897 24508
rect 9953 24506 9977 24508
rect 10033 24506 10057 24508
rect 9895 24454 9897 24506
rect 9959 24454 9971 24506
rect 10033 24454 10035 24506
rect 9873 24452 9897 24454
rect 9953 24452 9977 24454
rect 10033 24452 10057 24454
rect 9817 24432 10113 24452
rect 9817 23420 10113 23440
rect 9873 23418 9897 23420
rect 9953 23418 9977 23420
rect 10033 23418 10057 23420
rect 9895 23366 9897 23418
rect 9959 23366 9971 23418
rect 10033 23366 10035 23418
rect 9873 23364 9897 23366
rect 9953 23364 9977 23366
rect 10033 23364 10057 23366
rect 9817 23344 10113 23364
rect 9817 22332 10113 22352
rect 9873 22330 9897 22332
rect 9953 22330 9977 22332
rect 10033 22330 10057 22332
rect 9895 22278 9897 22330
rect 9959 22278 9971 22330
rect 10033 22278 10035 22330
rect 9873 22276 9897 22278
rect 9953 22276 9977 22278
rect 10033 22276 10057 22278
rect 9817 22256 10113 22276
rect 9817 21244 10113 21264
rect 9873 21242 9897 21244
rect 9953 21242 9977 21244
rect 10033 21242 10057 21244
rect 9895 21190 9897 21242
rect 9959 21190 9971 21242
rect 10033 21190 10035 21242
rect 9873 21188 9897 21190
rect 9953 21188 9977 21190
rect 10033 21188 10057 21190
rect 9817 21168 10113 21188
rect 9817 20156 10113 20176
rect 9873 20154 9897 20156
rect 9953 20154 9977 20156
rect 10033 20154 10057 20156
rect 9895 20102 9897 20154
rect 9959 20102 9971 20154
rect 10033 20102 10035 20154
rect 9873 20100 9897 20102
rect 9953 20100 9977 20102
rect 10033 20100 10057 20102
rect 9817 20080 10113 20100
rect 9817 19068 10113 19088
rect 9873 19066 9897 19068
rect 9953 19066 9977 19068
rect 10033 19066 10057 19068
rect 9895 19014 9897 19066
rect 9959 19014 9971 19066
rect 10033 19014 10035 19066
rect 9873 19012 9897 19014
rect 9953 19012 9977 19014
rect 10033 19012 10057 19014
rect 9817 18992 10113 19012
rect 10402 18728 10458 18737
rect 10402 18663 10458 18672
rect 8286 18048 8342 18057
rect 8286 17983 8342 17992
rect 9574 18048 9630 18057
rect 9574 17983 9630 17992
rect 5150 17436 5446 17456
rect 5206 17434 5230 17436
rect 5286 17434 5310 17436
rect 5366 17434 5390 17436
rect 5228 17382 5230 17434
rect 5292 17382 5304 17434
rect 5366 17382 5368 17434
rect 5206 17380 5230 17382
rect 5286 17380 5310 17382
rect 5366 17380 5390 17382
rect 5150 17360 5446 17380
rect 5150 16348 5446 16368
rect 5206 16346 5230 16348
rect 5286 16346 5310 16348
rect 5366 16346 5390 16348
rect 5228 16294 5230 16346
rect 5292 16294 5304 16346
rect 5366 16294 5368 16346
rect 5206 16292 5230 16294
rect 5286 16292 5310 16294
rect 5366 16292 5390 16294
rect 5150 16272 5446 16292
rect 5526 16144 5582 16153
rect 5526 16079 5582 16088
rect 5150 15260 5446 15280
rect 5206 15258 5230 15260
rect 5286 15258 5310 15260
rect 5366 15258 5390 15260
rect 5228 15206 5230 15258
rect 5292 15206 5304 15258
rect 5366 15206 5368 15258
rect 5206 15204 5230 15206
rect 5286 15204 5310 15206
rect 5366 15204 5390 15206
rect 5150 15184 5446 15204
rect 5150 14172 5446 14192
rect 5206 14170 5230 14172
rect 5286 14170 5310 14172
rect 5366 14170 5390 14172
rect 5228 14118 5230 14170
rect 5292 14118 5304 14170
rect 5366 14118 5368 14170
rect 5206 14116 5230 14118
rect 5286 14116 5310 14118
rect 5366 14116 5390 14118
rect 5150 14096 5446 14116
rect 5150 13084 5446 13104
rect 5206 13082 5230 13084
rect 5286 13082 5310 13084
rect 5366 13082 5390 13084
rect 5228 13030 5230 13082
rect 5292 13030 5304 13082
rect 5366 13030 5368 13082
rect 5206 13028 5230 13030
rect 5286 13028 5310 13030
rect 5366 13028 5390 13030
rect 5150 13008 5446 13028
rect 5066 12744 5122 12753
rect 5066 12679 5122 12688
rect 3686 11248 3742 11257
rect 3686 11183 3742 11192
rect 4422 10568 4478 10577
rect 4422 10503 4478 10512
rect 3318 8256 3374 8265
rect 3318 8191 3374 8200
rect 1662 7168 1718 7177
rect 1662 7103 1718 7112
rect 6 3768 62 3777
rect 6 3703 62 3712
rect 20 480 48 3703
rect 1018 2952 1074 2961
rect 1018 2887 1074 2896
rect 1032 480 1060 2887
rect 1676 2650 1704 7103
rect 2766 7032 2822 7041
rect 2766 6967 2822 6976
rect 2780 3194 2808 6967
rect 2768 3188 2820 3194
rect 2768 3130 2820 3136
rect 2780 2990 2808 3130
rect 2768 2984 2820 2990
rect 2768 2926 2820 2932
rect 3228 2848 3280 2854
rect 2030 2816 2086 2825
rect 3228 2790 3280 2796
rect 2030 2751 2086 2760
rect 1664 2644 1716 2650
rect 1664 2586 1716 2592
rect 2044 480 2072 2751
rect 3044 2508 3096 2514
rect 3044 2450 3096 2456
rect 3056 2310 3084 2450
rect 2124 2304 2176 2310
rect 2124 2246 2176 2252
rect 2860 2304 2912 2310
rect 2860 2246 2912 2252
rect 3044 2304 3096 2310
rect 3044 2246 3096 2252
rect 2136 1737 2164 2246
rect 2122 1728 2178 1737
rect 2122 1663 2178 1672
rect 2872 1465 2900 2246
rect 3056 2009 3084 2246
rect 3042 2000 3098 2009
rect 3042 1935 3098 1944
rect 3240 1737 3268 2790
rect 3226 1728 3282 1737
rect 3226 1663 3282 1672
rect 2858 1456 2914 1465
rect 3332 1442 3360 8191
rect 3778 6760 3834 6769
rect 3778 6695 3834 6704
rect 3410 4856 3466 4865
rect 3410 4791 3466 4800
rect 3424 3194 3452 4791
rect 3594 4040 3650 4049
rect 3594 3975 3650 3984
rect 3608 3942 3636 3975
rect 3596 3936 3648 3942
rect 3596 3878 3648 3884
rect 3792 3194 3820 6695
rect 4054 6488 4110 6497
rect 4054 6423 4110 6432
rect 4068 3738 4096 6423
rect 4148 3936 4200 3942
rect 4148 3878 4200 3884
rect 4056 3732 4108 3738
rect 4056 3674 4108 3680
rect 3962 3632 4018 3641
rect 3962 3567 3964 3576
rect 4016 3567 4018 3576
rect 3964 3538 4016 3544
rect 3976 3194 4004 3538
rect 3412 3188 3464 3194
rect 3412 3130 3464 3136
rect 3780 3188 3832 3194
rect 3780 3130 3832 3136
rect 3964 3188 4016 3194
rect 3964 3130 4016 3136
rect 3792 2990 3820 3130
rect 3780 2984 3832 2990
rect 3780 2926 3832 2932
rect 2858 1391 2914 1400
rect 3056 1414 3360 1442
rect 3056 480 3084 1414
rect 4160 480 4188 3878
rect 4436 3194 4464 10503
rect 4792 4684 4844 4690
rect 4792 4626 4844 4632
rect 4804 3942 4832 4626
rect 4974 4584 5030 4593
rect 4974 4519 4976 4528
rect 5028 4519 5030 4528
rect 4976 4490 5028 4496
rect 4608 3936 4660 3942
rect 4608 3878 4660 3884
rect 4792 3936 4844 3942
rect 4792 3878 4844 3884
rect 4620 3505 4648 3878
rect 4606 3496 4662 3505
rect 4606 3431 4662 3440
rect 4424 3188 4476 3194
rect 4424 3130 4476 3136
rect 4240 2984 4292 2990
rect 4238 2952 4240 2961
rect 4292 2952 4294 2961
rect 4238 2887 4294 2896
rect 4330 2816 4386 2825
rect 4330 2751 4386 2760
rect 4344 2514 4372 2751
rect 4514 2680 4570 2689
rect 4514 2615 4516 2624
rect 4568 2615 4570 2624
rect 4516 2586 4568 2592
rect 4332 2508 4384 2514
rect 4332 2450 4384 2456
rect 4804 1306 4832 3878
rect 5080 3602 5108 12679
rect 5150 11996 5446 12016
rect 5206 11994 5230 11996
rect 5286 11994 5310 11996
rect 5366 11994 5390 11996
rect 5228 11942 5230 11994
rect 5292 11942 5304 11994
rect 5366 11942 5368 11994
rect 5206 11940 5230 11942
rect 5286 11940 5310 11942
rect 5366 11940 5390 11942
rect 5150 11920 5446 11940
rect 5150 10908 5446 10928
rect 5206 10906 5230 10908
rect 5286 10906 5310 10908
rect 5366 10906 5390 10908
rect 5228 10854 5230 10906
rect 5292 10854 5304 10906
rect 5366 10854 5368 10906
rect 5206 10852 5230 10854
rect 5286 10852 5310 10854
rect 5366 10852 5390 10854
rect 5150 10832 5446 10852
rect 5150 9820 5446 9840
rect 5206 9818 5230 9820
rect 5286 9818 5310 9820
rect 5366 9818 5390 9820
rect 5228 9766 5230 9818
rect 5292 9766 5304 9818
rect 5366 9766 5368 9818
rect 5206 9764 5230 9766
rect 5286 9764 5310 9766
rect 5366 9764 5390 9766
rect 5150 9744 5446 9764
rect 5150 8732 5446 8752
rect 5206 8730 5230 8732
rect 5286 8730 5310 8732
rect 5366 8730 5390 8732
rect 5228 8678 5230 8730
rect 5292 8678 5304 8730
rect 5366 8678 5368 8730
rect 5206 8676 5230 8678
rect 5286 8676 5310 8678
rect 5366 8676 5390 8678
rect 5150 8656 5446 8676
rect 5150 7644 5446 7664
rect 5206 7642 5230 7644
rect 5286 7642 5310 7644
rect 5366 7642 5390 7644
rect 5228 7590 5230 7642
rect 5292 7590 5304 7642
rect 5366 7590 5368 7642
rect 5206 7588 5230 7590
rect 5286 7588 5310 7590
rect 5366 7588 5390 7590
rect 5150 7568 5446 7588
rect 5150 6556 5446 6576
rect 5206 6554 5230 6556
rect 5286 6554 5310 6556
rect 5366 6554 5390 6556
rect 5228 6502 5230 6554
rect 5292 6502 5304 6554
rect 5366 6502 5368 6554
rect 5206 6500 5230 6502
rect 5286 6500 5310 6502
rect 5366 6500 5390 6502
rect 5150 6480 5446 6500
rect 5150 5468 5446 5488
rect 5206 5466 5230 5468
rect 5286 5466 5310 5468
rect 5366 5466 5390 5468
rect 5228 5414 5230 5466
rect 5292 5414 5304 5466
rect 5366 5414 5368 5466
rect 5206 5412 5230 5414
rect 5286 5412 5310 5414
rect 5366 5412 5390 5414
rect 5150 5392 5446 5412
rect 5150 4380 5446 4400
rect 5206 4378 5230 4380
rect 5286 4378 5310 4380
rect 5366 4378 5390 4380
rect 5228 4326 5230 4378
rect 5292 4326 5304 4378
rect 5366 4326 5368 4378
rect 5206 4324 5230 4326
rect 5286 4324 5310 4326
rect 5366 4324 5390 4326
rect 5150 4304 5446 4324
rect 5540 4078 5568 16079
rect 8194 15464 8250 15473
rect 8194 15399 8250 15408
rect 7734 12064 7790 12073
rect 7734 11999 7790 12008
rect 7748 11898 7776 11999
rect 7736 11892 7788 11898
rect 7736 11834 7788 11840
rect 7748 11694 7776 11834
rect 7736 11688 7788 11694
rect 7736 11630 7788 11636
rect 8104 11620 8156 11626
rect 8104 11562 8156 11568
rect 7368 11552 7420 11558
rect 7368 11494 7420 11500
rect 7380 10849 7408 11494
rect 8116 11257 8144 11562
rect 8102 11248 8158 11257
rect 8102 11183 8104 11192
rect 8156 11183 8158 11192
rect 8104 11154 8156 11160
rect 7366 10840 7422 10849
rect 8116 10810 8144 11154
rect 7366 10775 7422 10784
rect 8104 10804 8156 10810
rect 8104 10746 8156 10752
rect 8208 9722 8236 15399
rect 9588 14550 9616 17983
rect 9817 17980 10113 18000
rect 9873 17978 9897 17980
rect 9953 17978 9977 17980
rect 10033 17978 10057 17980
rect 9895 17926 9897 17978
rect 9959 17926 9971 17978
rect 10033 17926 10035 17978
rect 9873 17924 9897 17926
rect 9953 17924 9977 17926
rect 10033 17924 10057 17926
rect 9817 17904 10113 17924
rect 9817 16892 10113 16912
rect 9873 16890 9897 16892
rect 9953 16890 9977 16892
rect 10033 16890 10057 16892
rect 9895 16838 9897 16890
rect 9959 16838 9971 16890
rect 10033 16838 10035 16890
rect 9873 16836 9897 16838
rect 9953 16836 9977 16838
rect 10033 16836 10057 16838
rect 9817 16816 10113 16836
rect 9817 15804 10113 15824
rect 9873 15802 9897 15804
rect 9953 15802 9977 15804
rect 10033 15802 10057 15804
rect 9895 15750 9897 15802
rect 9959 15750 9971 15802
rect 10033 15750 10035 15802
rect 9873 15748 9897 15750
rect 9953 15748 9977 15750
rect 10033 15748 10057 15750
rect 9817 15728 10113 15748
rect 9817 14716 10113 14736
rect 9873 14714 9897 14716
rect 9953 14714 9977 14716
rect 10033 14714 10057 14716
rect 9895 14662 9897 14714
rect 9959 14662 9971 14714
rect 10033 14662 10035 14714
rect 9873 14660 9897 14662
rect 9953 14660 9977 14662
rect 10033 14660 10057 14662
rect 9817 14640 10113 14660
rect 9576 14544 9628 14550
rect 9576 14486 9628 14492
rect 8930 14376 8986 14385
rect 8930 14311 8986 14320
rect 8944 14074 8972 14311
rect 9300 14272 9352 14278
rect 9300 14214 9352 14220
rect 8932 14068 8984 14074
rect 8932 14010 8984 14016
rect 8944 13870 8972 14010
rect 8932 13864 8984 13870
rect 8932 13806 8984 13812
rect 9208 13184 9260 13190
rect 9208 13126 9260 13132
rect 9220 12714 9248 13126
rect 9312 12986 9340 14214
rect 9588 14074 9616 14486
rect 9668 14476 9720 14482
rect 9668 14418 9720 14424
rect 9576 14068 9628 14074
rect 9576 14010 9628 14016
rect 9392 13864 9444 13870
rect 9392 13806 9444 13812
rect 9404 13394 9432 13806
rect 9588 13394 9616 14010
rect 9680 13938 9708 14418
rect 9668 13932 9720 13938
rect 9668 13874 9720 13880
rect 9817 13628 10113 13648
rect 9873 13626 9897 13628
rect 9953 13626 9977 13628
rect 10033 13626 10057 13628
rect 9895 13574 9897 13626
rect 9959 13574 9971 13626
rect 10033 13574 10035 13626
rect 9873 13572 9897 13574
rect 9953 13572 9977 13574
rect 10033 13572 10057 13574
rect 9817 13552 10113 13572
rect 9392 13388 9444 13394
rect 9392 13330 9444 13336
rect 9576 13388 9628 13394
rect 9576 13330 9628 13336
rect 9404 12986 9432 13330
rect 9482 13016 9538 13025
rect 9300 12980 9352 12986
rect 9300 12922 9352 12928
rect 9392 12980 9444 12986
rect 9482 12951 9538 12960
rect 9392 12922 9444 12928
rect 9312 12782 9340 12922
rect 9496 12918 9524 12951
rect 9588 12918 9616 13330
rect 9484 12912 9536 12918
rect 9484 12854 9536 12860
rect 9576 12912 9628 12918
rect 9576 12854 9628 12860
rect 10220 12912 10272 12918
rect 10220 12854 10272 12860
rect 9300 12776 9352 12782
rect 9300 12718 9352 12724
rect 9208 12708 9260 12714
rect 9208 12650 9260 12656
rect 8656 12300 8708 12306
rect 8656 12242 8708 12248
rect 8288 12096 8340 12102
rect 8288 12038 8340 12044
rect 8300 11801 8328 12038
rect 8668 11937 8696 12242
rect 8654 11928 8710 11937
rect 8654 11863 8656 11872
rect 8708 11863 8710 11872
rect 8656 11834 8708 11840
rect 8668 11803 8696 11834
rect 9116 11824 9168 11830
rect 8286 11792 8342 11801
rect 9220 11812 9248 12650
rect 9168 11784 9248 11812
rect 9116 11766 9168 11772
rect 8286 11727 8342 11736
rect 8380 11552 8432 11558
rect 8380 11494 8432 11500
rect 8286 11112 8342 11121
rect 8286 11047 8288 11056
rect 8340 11047 8342 11056
rect 8288 11018 8340 11024
rect 8392 9897 8420 11494
rect 9312 11286 9340 12718
rect 9817 12540 10113 12560
rect 9873 12538 9897 12540
rect 9953 12538 9977 12540
rect 10033 12538 10057 12540
rect 9895 12486 9897 12538
rect 9959 12486 9971 12538
rect 10033 12486 10035 12538
rect 9873 12484 9897 12486
rect 9953 12484 9977 12486
rect 10033 12484 10057 12486
rect 9817 12464 10113 12484
rect 9390 12336 9446 12345
rect 10232 12306 10260 12854
rect 9390 12271 9446 12280
rect 10220 12300 10272 12306
rect 9404 11898 9432 12271
rect 10220 12242 10272 12248
rect 9944 12096 9996 12102
rect 9944 12038 9996 12044
rect 9392 11892 9444 11898
rect 9392 11834 9444 11840
rect 9956 11694 9984 12038
rect 10232 11898 10260 12242
rect 10220 11892 10272 11898
rect 10220 11834 10272 11840
rect 9944 11688 9996 11694
rect 9944 11630 9996 11636
rect 10220 11688 10272 11694
rect 10220 11630 10272 11636
rect 9668 11620 9720 11626
rect 9668 11562 9720 11568
rect 9392 11348 9444 11354
rect 9392 11290 9444 11296
rect 9300 11280 9352 11286
rect 9300 11222 9352 11228
rect 8472 10736 8524 10742
rect 8470 10704 8472 10713
rect 8524 10704 8526 10713
rect 8470 10639 8526 10648
rect 9208 10532 9260 10538
rect 9208 10474 9260 10480
rect 9220 10130 9248 10474
rect 9208 10124 9260 10130
rect 9208 10066 9260 10072
rect 8378 9888 8434 9897
rect 8378 9823 8434 9832
rect 9220 9722 9248 10066
rect 7276 9716 7328 9722
rect 7276 9658 7328 9664
rect 8196 9716 8248 9722
rect 8196 9658 8248 9664
rect 9208 9716 9260 9722
rect 9208 9658 9260 9664
rect 6446 9072 6502 9081
rect 6446 9007 6502 9016
rect 5986 8936 6042 8945
rect 5986 8871 6042 8880
rect 5802 8800 5858 8809
rect 5802 8735 5858 8744
rect 5816 4826 5844 8735
rect 5804 4820 5856 4826
rect 5804 4762 5856 4768
rect 5712 4684 5764 4690
rect 5712 4626 5764 4632
rect 5528 4072 5580 4078
rect 5528 4014 5580 4020
rect 5724 3942 5752 4626
rect 5896 4004 5948 4010
rect 5896 3946 5948 3952
rect 5620 3936 5672 3942
rect 5620 3878 5672 3884
rect 5712 3936 5764 3942
rect 5712 3878 5764 3884
rect 5068 3596 5120 3602
rect 5068 3538 5120 3544
rect 4884 3392 4936 3398
rect 4884 3334 4936 3340
rect 4896 3097 4924 3334
rect 5080 3194 5108 3538
rect 5150 3292 5446 3312
rect 5206 3290 5230 3292
rect 5286 3290 5310 3292
rect 5366 3290 5390 3292
rect 5228 3238 5230 3290
rect 5292 3238 5304 3290
rect 5366 3238 5368 3290
rect 5206 3236 5230 3238
rect 5286 3236 5310 3238
rect 5366 3236 5390 3238
rect 5150 3216 5446 3236
rect 5068 3188 5120 3194
rect 5068 3130 5120 3136
rect 4882 3088 4938 3097
rect 4882 3023 4938 3032
rect 5344 2440 5396 2446
rect 5342 2408 5344 2417
rect 5396 2408 5398 2417
rect 5342 2343 5398 2352
rect 5150 2204 5446 2224
rect 5206 2202 5230 2204
rect 5286 2202 5310 2204
rect 5366 2202 5390 2204
rect 5228 2150 5230 2202
rect 5292 2150 5304 2202
rect 5366 2150 5368 2202
rect 5206 2148 5230 2150
rect 5286 2148 5310 2150
rect 5366 2148 5390 2150
rect 5150 2128 5446 2148
rect 4804 1278 5200 1306
rect 5172 480 5200 1278
rect 5632 1057 5660 3878
rect 5724 3777 5752 3878
rect 5710 3768 5766 3777
rect 5710 3703 5766 3712
rect 5802 3224 5858 3233
rect 5802 3159 5804 3168
rect 5856 3159 5858 3168
rect 5804 3130 5856 3136
rect 5804 2916 5856 2922
rect 5804 2858 5856 2864
rect 5816 1873 5844 2858
rect 5908 2825 5936 3946
rect 6000 3602 6028 8871
rect 6460 7041 6488 9007
rect 6446 7032 6502 7041
rect 6446 6967 6502 6976
rect 6538 6488 6594 6497
rect 6538 6423 6540 6432
rect 6592 6423 6594 6432
rect 6540 6394 6592 6400
rect 6172 6248 6224 6254
rect 6172 6190 6224 6196
rect 6078 3768 6134 3777
rect 6078 3703 6080 3712
rect 6132 3703 6134 3712
rect 6080 3674 6132 3680
rect 5988 3596 6040 3602
rect 5988 3538 6040 3544
rect 6000 3194 6028 3538
rect 5988 3188 6040 3194
rect 5988 3130 6040 3136
rect 5894 2816 5950 2825
rect 5894 2751 5950 2760
rect 5802 1864 5858 1873
rect 5802 1799 5858 1808
rect 5618 1048 5674 1057
rect 5618 983 5674 992
rect 6184 480 6212 6190
rect 6448 5772 6500 5778
rect 6448 5714 6500 5720
rect 6460 5409 6488 5714
rect 6446 5400 6502 5409
rect 6446 5335 6448 5344
rect 6500 5335 6502 5344
rect 6448 5306 6500 5312
rect 6460 5275 6488 5306
rect 6538 5264 6594 5273
rect 6538 5199 6540 5208
rect 6592 5199 6594 5208
rect 6540 5170 6592 5176
rect 6540 4616 6592 4622
rect 6540 4558 6592 4564
rect 6552 4185 6580 4558
rect 6538 4176 6594 4185
rect 6538 4111 6594 4120
rect 6724 3936 6776 3942
rect 6724 3878 6776 3884
rect 6736 2553 6764 3878
rect 6908 3528 6960 3534
rect 6908 3470 6960 3476
rect 6920 3369 6948 3470
rect 6906 3360 6962 3369
rect 6906 3295 6962 3304
rect 7184 2984 7236 2990
rect 7182 2952 7184 2961
rect 7236 2952 7238 2961
rect 7182 2887 7238 2896
rect 7182 2816 7238 2825
rect 7182 2751 7238 2760
rect 6722 2544 6778 2553
rect 6722 2479 6778 2488
rect 7196 480 7224 2751
rect 7288 2650 7316 9658
rect 8378 9616 8434 9625
rect 9300 9580 9352 9586
rect 8378 9551 8434 9560
rect 7826 9480 7882 9489
rect 7826 9415 7882 9424
rect 7734 7848 7790 7857
rect 7734 7783 7790 7792
rect 7748 7410 7776 7783
rect 7736 7404 7788 7410
rect 7736 7346 7788 7352
rect 7840 7177 7868 9415
rect 8194 7984 8250 7993
rect 8194 7919 8196 7928
rect 8248 7919 8250 7928
rect 8196 7890 8248 7896
rect 8208 7546 8236 7890
rect 8288 7880 8340 7886
rect 8286 7848 8288 7857
rect 8340 7848 8342 7857
rect 8286 7783 8342 7792
rect 8196 7540 8248 7546
rect 8196 7482 8248 7488
rect 8102 7304 8158 7313
rect 8102 7239 8158 7248
rect 7826 7168 7882 7177
rect 7826 7103 7882 7112
rect 8116 6866 8144 7239
rect 8104 6860 8156 6866
rect 8104 6802 8156 6808
rect 8102 6352 8158 6361
rect 8102 6287 8104 6296
rect 8156 6287 8158 6296
rect 8104 6258 8156 6264
rect 7734 6216 7790 6225
rect 7734 6151 7736 6160
rect 7788 6151 7790 6160
rect 7736 6122 7788 6128
rect 8194 5808 8250 5817
rect 7644 5772 7696 5778
rect 8194 5743 8196 5752
rect 7644 5714 7696 5720
rect 8248 5743 8250 5752
rect 8196 5714 8248 5720
rect 7656 5370 7684 5714
rect 7734 5672 7790 5681
rect 7734 5607 7736 5616
rect 7788 5607 7790 5616
rect 7736 5578 7788 5584
rect 7644 5364 7696 5370
rect 7644 5306 7696 5312
rect 8104 5160 8156 5166
rect 8104 5102 8156 5108
rect 8194 5128 8250 5137
rect 8116 4457 8144 5102
rect 8194 5063 8196 5072
rect 8248 5063 8250 5072
rect 8196 5034 8248 5040
rect 8196 4684 8248 4690
rect 8196 4626 8248 4632
rect 8102 4448 8158 4457
rect 8102 4383 8158 4392
rect 8208 4214 8236 4626
rect 8196 4208 8248 4214
rect 8196 4150 8248 4156
rect 7552 4072 7604 4078
rect 7552 4014 7604 4020
rect 7276 2644 7328 2650
rect 7276 2586 7328 2592
rect 7564 1601 7592 4014
rect 8392 3738 8420 9551
rect 9220 9540 9300 9568
rect 8930 8392 8986 8401
rect 8930 8327 8932 8336
rect 8984 8327 8986 8336
rect 8932 8298 8984 8304
rect 8654 7712 8710 7721
rect 8654 7647 8710 7656
rect 8472 5024 8524 5030
rect 8472 4966 8524 4972
rect 8484 4049 8512 4966
rect 8470 4040 8526 4049
rect 8470 3975 8526 3984
rect 8380 3732 8432 3738
rect 8380 3674 8432 3680
rect 8288 3596 8340 3602
rect 8288 3538 8340 3544
rect 8300 2854 8328 3538
rect 7644 2848 7696 2854
rect 8288 2848 8340 2854
rect 7644 2790 7696 2796
rect 7734 2816 7790 2825
rect 7550 1592 7606 1601
rect 7550 1527 7606 1536
rect 7656 921 7684 2790
rect 8288 2790 8340 2796
rect 7734 2751 7790 2760
rect 7748 2650 7776 2751
rect 7736 2644 7788 2650
rect 7736 2586 7788 2592
rect 7642 912 7698 921
rect 7642 847 7698 856
rect 8300 480 8328 2790
rect 8668 2650 8696 7647
rect 9220 6338 9248 9540
rect 9300 9522 9352 9528
rect 9404 8566 9432 11290
rect 9680 11218 9708 11562
rect 9817 11452 10113 11472
rect 9873 11450 9897 11452
rect 9953 11450 9977 11452
rect 10033 11450 10057 11452
rect 9895 11398 9897 11450
rect 9959 11398 9971 11450
rect 10033 11398 10035 11450
rect 9873 11396 9897 11398
rect 9953 11396 9977 11398
rect 10033 11396 10057 11398
rect 9817 11376 10113 11396
rect 10232 11354 10260 11630
rect 10220 11348 10272 11354
rect 10220 11290 10272 11296
rect 9668 11212 9720 11218
rect 9668 11154 9720 11160
rect 9680 10810 9708 11154
rect 9668 10804 9720 10810
rect 9668 10746 9720 10752
rect 9484 10464 9536 10470
rect 9484 10406 9536 10412
rect 9496 10169 9524 10406
rect 9482 10160 9538 10169
rect 9482 10095 9538 10104
rect 9484 10056 9536 10062
rect 9680 10033 9708 10746
rect 10312 10600 10364 10606
rect 10312 10542 10364 10548
rect 9817 10364 10113 10384
rect 9873 10362 9897 10364
rect 9953 10362 9977 10364
rect 10033 10362 10057 10364
rect 9895 10310 9897 10362
rect 9959 10310 9971 10362
rect 10033 10310 10035 10362
rect 9873 10308 9897 10310
rect 9953 10308 9977 10310
rect 10033 10308 10057 10310
rect 9817 10288 10113 10308
rect 9484 9998 9536 10004
rect 9666 10024 9722 10033
rect 9496 9654 9524 9998
rect 9666 9959 9722 9968
rect 10324 9926 10352 10542
rect 10416 10062 10444 18663
rect 11598 17096 11654 17105
rect 11598 17031 11654 17040
rect 10588 13864 10640 13870
rect 10588 13806 10640 13812
rect 10496 13184 10548 13190
rect 10496 13126 10548 13132
rect 10508 12714 10536 13126
rect 10600 12986 10628 13806
rect 11416 13796 11468 13802
rect 11416 13738 11468 13744
rect 10680 13728 10732 13734
rect 10680 13670 10732 13676
rect 10692 13190 10720 13670
rect 10680 13184 10732 13190
rect 10680 13126 10732 13132
rect 10588 12980 10640 12986
rect 10588 12922 10640 12928
rect 10496 12708 10548 12714
rect 10496 12650 10548 12656
rect 10508 12306 10536 12650
rect 10600 12442 10628 12922
rect 10692 12850 10720 13126
rect 11428 12986 11456 13738
rect 11416 12980 11468 12986
rect 11416 12922 11468 12928
rect 10680 12844 10732 12850
rect 10680 12786 10732 12792
rect 10864 12640 10916 12646
rect 10864 12582 10916 12588
rect 11324 12640 11376 12646
rect 11324 12582 11376 12588
rect 10588 12436 10640 12442
rect 10588 12378 10640 12384
rect 10496 12300 10548 12306
rect 10496 12242 10548 12248
rect 10772 11688 10824 11694
rect 10772 11630 10824 11636
rect 10588 11552 10640 11558
rect 10588 11494 10640 11500
rect 10678 11520 10734 11529
rect 10600 10146 10628 11494
rect 10678 11455 10734 11464
rect 10692 10577 10720 11455
rect 10784 11082 10812 11630
rect 10772 11076 10824 11082
rect 10772 11018 10824 11024
rect 10784 10606 10812 11018
rect 10772 10600 10824 10606
rect 10678 10568 10734 10577
rect 10772 10542 10824 10548
rect 10678 10503 10734 10512
rect 10784 10266 10812 10542
rect 10772 10260 10824 10266
rect 10772 10202 10824 10208
rect 10508 10130 10628 10146
rect 10680 10192 10732 10198
rect 10680 10134 10732 10140
rect 10496 10124 10628 10130
rect 10548 10118 10628 10124
rect 10496 10066 10548 10072
rect 10404 10056 10456 10062
rect 10404 9998 10456 10004
rect 10312 9920 10364 9926
rect 10312 9862 10364 9868
rect 9666 9752 9722 9761
rect 9666 9687 9722 9696
rect 9484 9648 9536 9654
rect 9484 9590 9536 9596
rect 9484 9512 9536 9518
rect 9484 9454 9536 9460
rect 9392 8560 9444 8566
rect 9392 8502 9444 8508
rect 9404 7954 9432 8502
rect 9496 8265 9524 9454
rect 9482 8256 9538 8265
rect 9482 8191 9538 8200
rect 9392 7948 9444 7954
rect 9392 7890 9444 7896
rect 9298 7440 9354 7449
rect 9404 7410 9432 7890
rect 9298 7375 9354 7384
rect 9392 7404 9444 7410
rect 9312 7342 9340 7375
rect 9392 7346 9444 7352
rect 9300 7336 9352 7342
rect 9300 7278 9352 7284
rect 9312 6934 9340 7278
rect 9300 6928 9352 6934
rect 9300 6870 9352 6876
rect 9220 6310 9340 6338
rect 9208 6248 9260 6254
rect 9208 6190 9260 6196
rect 8840 6112 8892 6118
rect 8840 6054 8892 6060
rect 8852 5370 8880 6054
rect 9220 5846 9248 6190
rect 9208 5840 9260 5846
rect 9208 5782 9260 5788
rect 9312 5710 9340 6310
rect 8932 5704 8984 5710
rect 8932 5646 8984 5652
rect 9300 5704 9352 5710
rect 9300 5646 9352 5652
rect 8840 5364 8892 5370
rect 8840 5306 8892 5312
rect 8852 5030 8880 5306
rect 8840 5024 8892 5030
rect 8840 4966 8892 4972
rect 8838 3088 8894 3097
rect 8838 3023 8840 3032
rect 8892 3023 8894 3032
rect 8840 2994 8892 3000
rect 8656 2644 8708 2650
rect 8656 2586 8708 2592
rect 8748 2508 8800 2514
rect 8748 2450 8800 2456
rect 8760 2310 8788 2450
rect 8748 2304 8800 2310
rect 8746 2272 8748 2281
rect 8800 2272 8802 2281
rect 8746 2207 8802 2216
rect 8944 1329 8972 5646
rect 9312 5302 9340 5646
rect 9300 5296 9352 5302
rect 9300 5238 9352 5244
rect 9574 4856 9630 4865
rect 9574 4791 9630 4800
rect 9482 4720 9538 4729
rect 9482 4655 9484 4664
rect 9536 4655 9538 4664
rect 9484 4626 9536 4632
rect 9116 4616 9168 4622
rect 9116 4558 9168 4564
rect 9128 4434 9156 4558
rect 9128 4406 9248 4434
rect 9114 4312 9170 4321
rect 9114 4247 9170 4256
rect 9128 4078 9156 4247
rect 9116 4072 9168 4078
rect 9022 4040 9078 4049
rect 9116 4014 9168 4020
rect 9022 3975 9078 3984
rect 9036 3942 9064 3975
rect 9024 3936 9076 3942
rect 9024 3878 9076 3884
rect 9220 3670 9248 4406
rect 9588 4185 9616 4791
rect 9298 4176 9354 4185
rect 9298 4111 9354 4120
rect 9574 4176 9630 4185
rect 9574 4111 9630 4120
rect 9208 3664 9260 3670
rect 9208 3606 9260 3612
rect 9312 3534 9340 4111
rect 9300 3528 9352 3534
rect 9300 3470 9352 3476
rect 9312 3194 9340 3470
rect 9392 3392 9444 3398
rect 9392 3334 9444 3340
rect 9300 3188 9352 3194
rect 9300 3130 9352 3136
rect 9208 3052 9260 3058
rect 9404 3040 9432 3334
rect 9680 3074 9708 9687
rect 10220 9648 10272 9654
rect 10220 9590 10272 9596
rect 9817 9276 10113 9296
rect 9873 9274 9897 9276
rect 9953 9274 9977 9276
rect 10033 9274 10057 9276
rect 9895 9222 9897 9274
rect 9959 9222 9971 9274
rect 10033 9222 10035 9274
rect 9873 9220 9897 9222
rect 9953 9220 9977 9222
rect 10033 9220 10057 9222
rect 9817 9200 10113 9220
rect 10232 9042 10260 9590
rect 10220 9036 10272 9042
rect 10220 8978 10272 8984
rect 10232 8634 10260 8978
rect 10220 8628 10272 8634
rect 10220 8570 10272 8576
rect 9817 8188 10113 8208
rect 9873 8186 9897 8188
rect 9953 8186 9977 8188
rect 10033 8186 10057 8188
rect 9895 8134 9897 8186
rect 9959 8134 9971 8186
rect 10033 8134 10035 8186
rect 9873 8132 9897 8134
rect 9953 8132 9977 8134
rect 10033 8132 10057 8134
rect 9817 8112 10113 8132
rect 10218 8120 10274 8129
rect 10218 8055 10274 8064
rect 10232 7721 10260 8055
rect 10218 7712 10274 7721
rect 10218 7647 10274 7656
rect 10324 7546 10352 9862
rect 10600 9654 10628 10118
rect 10588 9648 10640 9654
rect 10588 9590 10640 9596
rect 10692 9586 10720 10134
rect 10680 9580 10732 9586
rect 10680 9522 10732 9528
rect 10404 9444 10456 9450
rect 10404 9386 10456 9392
rect 10496 9444 10548 9450
rect 10496 9386 10548 9392
rect 10416 9178 10444 9386
rect 10404 9172 10456 9178
rect 10404 9114 10456 9120
rect 10508 9042 10536 9386
rect 10692 9110 10720 9522
rect 10680 9104 10732 9110
rect 10680 9046 10732 9052
rect 10496 9036 10548 9042
rect 10496 8978 10548 8984
rect 10402 8664 10458 8673
rect 10402 8599 10458 8608
rect 10416 8430 10444 8599
rect 10496 8492 10548 8498
rect 10496 8434 10548 8440
rect 10404 8424 10456 8430
rect 10404 8366 10456 8372
rect 10416 8090 10444 8366
rect 10404 8084 10456 8090
rect 10404 8026 10456 8032
rect 10404 7880 10456 7886
rect 10404 7822 10456 7828
rect 10312 7540 10364 7546
rect 10312 7482 10364 7488
rect 10324 7342 10352 7482
rect 10312 7336 10364 7342
rect 10312 7278 10364 7284
rect 10220 7268 10272 7274
rect 10220 7210 10272 7216
rect 9817 7100 10113 7120
rect 9873 7098 9897 7100
rect 9953 7098 9977 7100
rect 10033 7098 10057 7100
rect 9895 7046 9897 7098
rect 9959 7046 9971 7098
rect 10033 7046 10035 7098
rect 9873 7044 9897 7046
rect 9953 7044 9977 7046
rect 10033 7044 10057 7046
rect 9817 7024 10113 7044
rect 10232 7041 10260 7210
rect 10416 7177 10444 7822
rect 10402 7168 10458 7177
rect 10402 7103 10458 7112
rect 10218 7032 10274 7041
rect 10218 6967 10274 6976
rect 10508 6866 10536 8434
rect 10588 8084 10640 8090
rect 10588 8026 10640 8032
rect 10496 6860 10548 6866
rect 10496 6802 10548 6808
rect 10404 6452 10456 6458
rect 10404 6394 10456 6400
rect 10416 6186 10444 6394
rect 10404 6180 10456 6186
rect 10404 6122 10456 6128
rect 10402 6080 10458 6089
rect 9817 6012 10113 6032
rect 10402 6015 10458 6024
rect 9873 6010 9897 6012
rect 9953 6010 9977 6012
rect 10033 6010 10057 6012
rect 9895 5958 9897 6010
rect 9959 5958 9971 6010
rect 10033 5958 10035 6010
rect 9873 5956 9897 5958
rect 9953 5956 9977 5958
rect 10033 5956 10057 5958
rect 9817 5936 10113 5956
rect 10036 5840 10088 5846
rect 10036 5782 10088 5788
rect 9760 5704 9812 5710
rect 9760 5646 9812 5652
rect 9772 5234 9800 5646
rect 10048 5370 10076 5782
rect 10218 5400 10274 5409
rect 10036 5364 10088 5370
rect 10218 5335 10274 5344
rect 10036 5306 10088 5312
rect 9760 5228 9812 5234
rect 9760 5170 9812 5176
rect 9817 4924 10113 4944
rect 9873 4922 9897 4924
rect 9953 4922 9977 4924
rect 10033 4922 10057 4924
rect 9895 4870 9897 4922
rect 9959 4870 9971 4922
rect 10033 4870 10035 4922
rect 9873 4868 9897 4870
rect 9953 4868 9977 4870
rect 10033 4868 10057 4870
rect 9817 4848 10113 4868
rect 10232 3890 10260 5335
rect 10312 5228 10364 5234
rect 10312 5170 10364 5176
rect 10324 4826 10352 5170
rect 10312 4820 10364 4826
rect 10312 4762 10364 4768
rect 10324 4214 10352 4762
rect 10312 4208 10364 4214
rect 10312 4150 10364 4156
rect 10312 3936 10364 3942
rect 10232 3884 10312 3890
rect 10232 3878 10364 3884
rect 10232 3862 10352 3878
rect 9817 3836 10113 3856
rect 9873 3834 9897 3836
rect 9953 3834 9977 3836
rect 10033 3834 10057 3836
rect 9895 3782 9897 3834
rect 9959 3782 9971 3834
rect 10033 3782 10035 3834
rect 9873 3780 9897 3782
rect 9953 3780 9977 3782
rect 10033 3780 10057 3782
rect 9817 3760 10113 3780
rect 10128 3664 10180 3670
rect 10128 3606 10180 3612
rect 10140 3194 10168 3606
rect 10232 3534 10260 3862
rect 10220 3528 10272 3534
rect 10220 3470 10272 3476
rect 10416 3194 10444 6015
rect 10508 5914 10536 6802
rect 10496 5908 10548 5914
rect 10496 5850 10548 5856
rect 10600 5080 10628 8026
rect 10692 6866 10720 9046
rect 10770 8256 10826 8265
rect 10770 8191 10826 8200
rect 10784 7954 10812 8191
rect 10772 7948 10824 7954
rect 10772 7890 10824 7896
rect 10784 6866 10812 7890
rect 10876 7449 10904 12582
rect 11048 12300 11100 12306
rect 11048 12242 11100 12248
rect 11060 11354 11088 12242
rect 11336 12102 11364 12582
rect 11416 12232 11468 12238
rect 11414 12200 11416 12209
rect 11468 12200 11470 12209
rect 11414 12135 11470 12144
rect 11232 12096 11284 12102
rect 11232 12038 11284 12044
rect 11324 12096 11376 12102
rect 11324 12038 11376 12044
rect 11138 11928 11194 11937
rect 11138 11863 11140 11872
rect 11192 11863 11194 11872
rect 11140 11834 11192 11840
rect 11048 11348 11100 11354
rect 11048 11290 11100 11296
rect 11244 11082 11272 12038
rect 11336 11898 11364 12038
rect 11324 11892 11376 11898
rect 11324 11834 11376 11840
rect 11232 11076 11284 11082
rect 11232 11018 11284 11024
rect 11336 11014 11364 11834
rect 11428 11150 11456 12135
rect 11508 12096 11560 12102
rect 11508 12038 11560 12044
rect 11520 11694 11548 12038
rect 11508 11688 11560 11694
rect 11508 11630 11560 11636
rect 11416 11144 11468 11150
rect 11416 11086 11468 11092
rect 11508 11144 11560 11150
rect 11508 11086 11560 11092
rect 11324 11008 11376 11014
rect 11324 10950 11376 10956
rect 11336 10810 11364 10950
rect 11324 10804 11376 10810
rect 11324 10746 11376 10752
rect 11048 10532 11100 10538
rect 11048 10474 11100 10480
rect 11232 10532 11284 10538
rect 11232 10474 11284 10480
rect 11060 9042 11088 10474
rect 11244 10266 11272 10474
rect 11428 10266 11456 11086
rect 11232 10260 11284 10266
rect 11232 10202 11284 10208
rect 11416 10260 11468 10266
rect 11416 10202 11468 10208
rect 11244 9722 11272 10202
rect 11232 9716 11284 9722
rect 11232 9658 11284 9664
rect 11232 9104 11284 9110
rect 11232 9046 11284 9052
rect 11048 9036 11100 9042
rect 11048 8978 11100 8984
rect 11060 8090 11088 8978
rect 11244 8634 11272 9046
rect 11232 8628 11284 8634
rect 11232 8570 11284 8576
rect 11048 8084 11100 8090
rect 11048 8026 11100 8032
rect 11520 7954 11548 11086
rect 11508 7948 11560 7954
rect 11508 7890 11560 7896
rect 11520 7546 11548 7890
rect 11508 7540 11560 7546
rect 11508 7482 11560 7488
rect 10862 7440 10918 7449
rect 10862 7375 10918 7384
rect 11048 7268 11100 7274
rect 11048 7210 11100 7216
rect 10680 6860 10732 6866
rect 10680 6802 10732 6808
rect 10772 6860 10824 6866
rect 10772 6802 10824 6808
rect 10692 6458 10720 6802
rect 10862 6760 10918 6769
rect 10862 6695 10918 6704
rect 10772 6656 10824 6662
rect 10772 6598 10824 6604
rect 10680 6452 10732 6458
rect 10680 6394 10732 6400
rect 10680 6112 10732 6118
rect 10680 6054 10732 6060
rect 10508 5052 10628 5080
rect 10508 4690 10536 5052
rect 10496 4684 10548 4690
rect 10496 4626 10548 4632
rect 10508 4162 10536 4626
rect 10508 4134 10628 4162
rect 10600 3738 10628 4134
rect 10692 4010 10720 6054
rect 10784 5846 10812 6598
rect 10876 6361 10904 6695
rect 10862 6352 10918 6361
rect 10862 6287 10918 6296
rect 10864 6248 10916 6254
rect 10864 6190 10916 6196
rect 10876 5914 10904 6190
rect 10864 5908 10916 5914
rect 10864 5850 10916 5856
rect 10772 5840 10824 5846
rect 10772 5782 10824 5788
rect 11060 5778 11088 7210
rect 11416 6452 11468 6458
rect 11416 6394 11468 6400
rect 11428 5846 11456 6394
rect 11416 5840 11468 5846
rect 11416 5782 11468 5788
rect 11048 5772 11100 5778
rect 11048 5714 11100 5720
rect 11060 5370 11088 5714
rect 11048 5364 11100 5370
rect 11048 5306 11100 5312
rect 11324 5024 11376 5030
rect 11324 4966 11376 4972
rect 11336 4758 11364 4966
rect 11324 4752 11376 4758
rect 11324 4694 11376 4700
rect 11336 4282 11364 4694
rect 11416 4480 11468 4486
rect 11416 4422 11468 4428
rect 11324 4276 11376 4282
rect 11324 4218 11376 4224
rect 10680 4004 10732 4010
rect 10680 3946 10732 3952
rect 10588 3732 10640 3738
rect 10588 3674 10640 3680
rect 11324 3664 11376 3670
rect 11428 3652 11456 4422
rect 11376 3624 11456 3652
rect 11324 3606 11376 3612
rect 10128 3188 10180 3194
rect 10128 3130 10180 3136
rect 10404 3188 10456 3194
rect 10404 3130 10456 3136
rect 9680 3046 10260 3074
rect 9260 3012 9432 3040
rect 9208 2994 9260 3000
rect 9116 2984 9168 2990
rect 9116 2926 9168 2932
rect 8930 1320 8986 1329
rect 8930 1255 8986 1264
rect 9128 1193 9156 2926
rect 9298 2816 9354 2825
rect 9298 2751 9354 2760
rect 9114 1184 9170 1193
rect 9114 1119 9170 1128
rect 9312 480 9340 2751
rect 9404 2689 9432 3012
rect 9817 2748 10113 2768
rect 9873 2746 9897 2748
rect 9953 2746 9977 2748
rect 10033 2746 10057 2748
rect 9895 2694 9897 2746
rect 9959 2694 9971 2746
rect 10033 2694 10035 2746
rect 9873 2692 9897 2694
rect 9953 2692 9977 2694
rect 10033 2692 10057 2694
rect 9390 2680 9446 2689
rect 9817 2672 10113 2692
rect 10232 2650 10260 3046
rect 10404 2916 10456 2922
rect 10404 2858 10456 2864
rect 10496 2916 10548 2922
rect 10496 2858 10548 2864
rect 10416 2825 10444 2858
rect 10402 2816 10458 2825
rect 10402 2751 10458 2760
rect 9390 2615 9446 2624
rect 10220 2644 10272 2650
rect 10220 2586 10272 2592
rect 10508 2446 10536 2858
rect 11336 2854 11364 3606
rect 11612 3534 11640 17031
rect 11796 15434 11824 27520
rect 15292 27418 15320 27520
rect 14924 27390 15320 27418
rect 14484 25052 14780 25072
rect 14540 25050 14564 25052
rect 14620 25050 14644 25052
rect 14700 25050 14724 25052
rect 14562 24998 14564 25050
rect 14626 24998 14638 25050
rect 14700 24998 14702 25050
rect 14540 24996 14564 24998
rect 14620 24996 14644 24998
rect 14700 24996 14724 24998
rect 14484 24976 14780 24996
rect 14484 23964 14780 23984
rect 14540 23962 14564 23964
rect 14620 23962 14644 23964
rect 14700 23962 14724 23964
rect 14562 23910 14564 23962
rect 14626 23910 14638 23962
rect 14700 23910 14702 23962
rect 14540 23908 14564 23910
rect 14620 23908 14644 23910
rect 14700 23908 14724 23910
rect 14484 23888 14780 23908
rect 14484 22876 14780 22896
rect 14540 22874 14564 22876
rect 14620 22874 14644 22876
rect 14700 22874 14724 22876
rect 14562 22822 14564 22874
rect 14626 22822 14638 22874
rect 14700 22822 14702 22874
rect 14540 22820 14564 22822
rect 14620 22820 14644 22822
rect 14700 22820 14724 22822
rect 14484 22800 14780 22820
rect 14484 21788 14780 21808
rect 14540 21786 14564 21788
rect 14620 21786 14644 21788
rect 14700 21786 14724 21788
rect 14562 21734 14564 21786
rect 14626 21734 14638 21786
rect 14700 21734 14702 21786
rect 14540 21732 14564 21734
rect 14620 21732 14644 21734
rect 14700 21732 14724 21734
rect 14484 21712 14780 21732
rect 14484 20700 14780 20720
rect 14540 20698 14564 20700
rect 14620 20698 14644 20700
rect 14700 20698 14724 20700
rect 14562 20646 14564 20698
rect 14626 20646 14638 20698
rect 14700 20646 14702 20698
rect 14540 20644 14564 20646
rect 14620 20644 14644 20646
rect 14700 20644 14724 20646
rect 14484 20624 14780 20644
rect 14484 19612 14780 19632
rect 14540 19610 14564 19612
rect 14620 19610 14644 19612
rect 14700 19610 14724 19612
rect 14562 19558 14564 19610
rect 14626 19558 14638 19610
rect 14700 19558 14702 19610
rect 14540 19556 14564 19558
rect 14620 19556 14644 19558
rect 14700 19556 14724 19558
rect 14484 19536 14780 19556
rect 13254 19272 13310 19281
rect 13254 19207 13310 19216
rect 12426 16688 12482 16697
rect 12426 16623 12482 16632
rect 11784 15428 11836 15434
rect 11784 15370 11836 15376
rect 12152 15428 12204 15434
rect 12152 15370 12204 15376
rect 11876 14476 11928 14482
rect 11876 14418 11928 14424
rect 11784 14000 11836 14006
rect 11784 13942 11836 13948
rect 11796 13326 11824 13942
rect 11888 13734 11916 14418
rect 11876 13728 11928 13734
rect 11928 13676 12008 13682
rect 11876 13670 12008 13676
rect 11888 13654 12008 13670
rect 11876 13388 11928 13394
rect 11876 13330 11928 13336
rect 11784 13320 11836 13326
rect 11784 13262 11836 13268
rect 11692 13184 11744 13190
rect 11692 13126 11744 13132
rect 11784 13184 11836 13190
rect 11784 13126 11836 13132
rect 11704 12889 11732 13126
rect 11690 12880 11746 12889
rect 11690 12815 11746 12824
rect 11692 11552 11744 11558
rect 11796 11540 11824 13126
rect 11888 12481 11916 13330
rect 11874 12472 11930 12481
rect 11874 12407 11930 12416
rect 11980 12102 12008 13654
rect 12060 12980 12112 12986
rect 12060 12922 12112 12928
rect 11968 12096 12020 12102
rect 11968 12038 12020 12044
rect 12072 11694 12100 12922
rect 12164 12918 12192 15370
rect 12336 14272 12388 14278
rect 12336 14214 12388 14220
rect 12152 12912 12204 12918
rect 12152 12854 12204 12860
rect 12244 12640 12296 12646
rect 12244 12582 12296 12588
rect 12256 12442 12284 12582
rect 12244 12436 12296 12442
rect 12244 12378 12296 12384
rect 12256 11830 12284 12378
rect 12348 12209 12376 14214
rect 12334 12200 12390 12209
rect 12334 12135 12390 12144
rect 12336 12096 12388 12102
rect 12336 12038 12388 12044
rect 12244 11824 12296 11830
rect 12244 11766 12296 11772
rect 12060 11688 12112 11694
rect 12060 11630 12112 11636
rect 11968 11620 12020 11626
rect 11888 11580 11968 11608
rect 11888 11540 11916 11580
rect 11968 11562 12020 11568
rect 11744 11512 11916 11540
rect 11692 11494 11744 11500
rect 11704 11286 11732 11494
rect 12256 11354 12284 11766
rect 12348 11762 12376 12038
rect 12440 11778 12468 16623
rect 13070 15600 13126 15609
rect 12888 15564 12940 15570
rect 13070 15535 13072 15544
rect 12888 15506 12940 15512
rect 13124 15535 13126 15544
rect 13072 15506 13124 15512
rect 12612 15496 12664 15502
rect 12612 15438 12664 15444
rect 12520 15156 12572 15162
rect 12520 15098 12572 15104
rect 12532 13870 12560 15098
rect 12624 15094 12652 15438
rect 12900 15162 12928 15506
rect 12888 15156 12940 15162
rect 12888 15098 12940 15104
rect 12612 15088 12664 15094
rect 12612 15030 12664 15036
rect 13084 14618 13112 15506
rect 13164 15360 13216 15366
rect 13164 15302 13216 15308
rect 13176 15162 13204 15302
rect 13164 15156 13216 15162
rect 13164 15098 13216 15104
rect 13072 14612 13124 14618
rect 13072 14554 13124 14560
rect 13084 13870 13112 14554
rect 12520 13864 12572 13870
rect 12520 13806 12572 13812
rect 13072 13864 13124 13870
rect 13072 13806 13124 13812
rect 12532 13530 12560 13806
rect 12520 13524 12572 13530
rect 12520 13466 12572 13472
rect 13072 13388 13124 13394
rect 13072 13330 13124 13336
rect 13084 12646 13112 13330
rect 13072 12640 13124 12646
rect 13070 12608 13072 12617
rect 13124 12608 13126 12617
rect 13070 12543 13126 12552
rect 12518 12472 12574 12481
rect 13268 12424 13296 19207
rect 14484 18524 14780 18544
rect 14540 18522 14564 18524
rect 14620 18522 14644 18524
rect 14700 18522 14724 18524
rect 14562 18470 14564 18522
rect 14626 18470 14638 18522
rect 14700 18470 14702 18522
rect 14540 18468 14564 18470
rect 14620 18468 14644 18470
rect 14700 18468 14724 18470
rect 14484 18448 14780 18468
rect 14484 17436 14780 17456
rect 14540 17434 14564 17436
rect 14620 17434 14644 17436
rect 14700 17434 14724 17436
rect 14562 17382 14564 17434
rect 14626 17382 14638 17434
rect 14700 17382 14702 17434
rect 14540 17380 14564 17382
rect 14620 17380 14644 17382
rect 14700 17380 14724 17382
rect 14484 17360 14780 17380
rect 14924 16776 14952 27390
rect 16014 18320 16070 18329
rect 16014 18255 16070 18264
rect 16028 16794 16056 18255
rect 17854 17368 17910 17377
rect 17854 17303 17910 17312
rect 16200 17128 16252 17134
rect 16200 17070 16252 17076
rect 14832 16748 14952 16776
rect 15648 16788 15700 16794
rect 14484 16348 14780 16368
rect 14540 16346 14564 16348
rect 14620 16346 14644 16348
rect 14700 16346 14724 16348
rect 14562 16294 14564 16346
rect 14626 16294 14638 16346
rect 14700 16294 14702 16346
rect 14540 16292 14564 16294
rect 14620 16292 14644 16294
rect 14700 16292 14724 16294
rect 14484 16272 14780 16292
rect 14832 15502 14860 16748
rect 15648 16730 15700 16736
rect 16016 16788 16068 16794
rect 16016 16730 16068 16736
rect 14912 16652 14964 16658
rect 14912 16594 14964 16600
rect 13624 15496 13676 15502
rect 13624 15438 13676 15444
rect 14820 15496 14872 15502
rect 14820 15438 14872 15444
rect 13532 15360 13584 15366
rect 13532 15302 13584 15308
rect 13440 14952 13492 14958
rect 13440 14894 13492 14900
rect 13452 14482 13480 14894
rect 13440 14476 13492 14482
rect 13440 14418 13492 14424
rect 13452 13870 13480 14418
rect 13440 13864 13492 13870
rect 13440 13806 13492 13812
rect 13348 12708 13400 12714
rect 13348 12650 13400 12656
rect 13360 12442 13388 12650
rect 12518 12407 12574 12416
rect 12532 12374 12560 12407
rect 13176 12396 13296 12424
rect 13348 12436 13400 12442
rect 12520 12368 12572 12374
rect 12520 12310 12572 12316
rect 12336 11756 12388 11762
rect 12440 11750 12560 11778
rect 12336 11698 12388 11704
rect 12244 11348 12296 11354
rect 12244 11290 12296 11296
rect 12348 11286 12376 11698
rect 12428 11688 12480 11694
rect 12428 11630 12480 11636
rect 12440 11354 12468 11630
rect 12428 11348 12480 11354
rect 12428 11290 12480 11296
rect 11692 11280 11744 11286
rect 11692 11222 11744 11228
rect 12336 11280 12388 11286
rect 12336 11222 12388 11228
rect 11704 10810 11732 11222
rect 11784 11076 11836 11082
rect 11784 11018 11836 11024
rect 11692 10804 11744 10810
rect 11692 10746 11744 10752
rect 11796 9926 11824 11018
rect 12532 10674 12560 11750
rect 12612 11552 12664 11558
rect 12612 11494 12664 11500
rect 12520 10668 12572 10674
rect 12520 10610 12572 10616
rect 12152 10532 12204 10538
rect 12152 10474 12204 10480
rect 12164 10266 12192 10474
rect 12060 10260 12112 10266
rect 12060 10202 12112 10208
rect 12152 10260 12204 10266
rect 12152 10202 12204 10208
rect 11784 9920 11836 9926
rect 11784 9862 11836 9868
rect 12072 9654 12100 10202
rect 12060 9648 12112 9654
rect 12060 9590 12112 9596
rect 11968 9376 12020 9382
rect 11968 9318 12020 9324
rect 11980 8974 12008 9318
rect 12072 9178 12100 9590
rect 12532 9178 12560 10610
rect 12060 9172 12112 9178
rect 12060 9114 12112 9120
rect 12520 9172 12572 9178
rect 12520 9114 12572 9120
rect 11968 8968 12020 8974
rect 11968 8910 12020 8916
rect 12072 8566 12100 9114
rect 12624 8673 12652 11494
rect 13072 11212 13124 11218
rect 13072 11154 13124 11160
rect 13084 10810 13112 11154
rect 13072 10804 13124 10810
rect 13072 10746 13124 10752
rect 12796 10532 12848 10538
rect 12796 10474 12848 10480
rect 12808 10062 12836 10474
rect 12796 10056 12848 10062
rect 12796 9998 12848 10004
rect 12704 9988 12756 9994
rect 12704 9930 12756 9936
rect 12716 8945 12744 9930
rect 12808 9586 12836 9998
rect 12796 9580 12848 9586
rect 12796 9522 12848 9528
rect 12808 9178 12836 9522
rect 12796 9172 12848 9178
rect 12796 9114 12848 9120
rect 13072 9104 13124 9110
rect 13072 9046 13124 9052
rect 12980 8968 13032 8974
rect 12702 8936 12758 8945
rect 12980 8910 13032 8916
rect 12702 8871 12758 8880
rect 12610 8664 12666 8673
rect 12610 8599 12666 8608
rect 12060 8560 12112 8566
rect 12060 8502 12112 8508
rect 12334 8528 12390 8537
rect 12334 8463 12390 8472
rect 12348 7818 12376 8463
rect 12624 8090 12652 8599
rect 12992 8090 13020 8910
rect 13084 8498 13112 9046
rect 13072 8492 13124 8498
rect 13072 8434 13124 8440
rect 12612 8084 12664 8090
rect 12612 8026 12664 8032
rect 12980 8084 13032 8090
rect 12980 8026 13032 8032
rect 12520 7948 12572 7954
rect 12520 7890 12572 7896
rect 12336 7812 12388 7818
rect 12336 7754 12388 7760
rect 12150 7440 12206 7449
rect 12150 7375 12206 7384
rect 11692 7200 11744 7206
rect 11692 7142 11744 7148
rect 11968 7200 12020 7206
rect 11968 7142 12020 7148
rect 11704 6866 11732 7142
rect 11692 6860 11744 6866
rect 11692 6802 11744 6808
rect 11704 6118 11732 6802
rect 11782 6760 11838 6769
rect 11782 6695 11838 6704
rect 11692 6112 11744 6118
rect 11692 6054 11744 6060
rect 11796 5166 11824 6695
rect 11980 5930 12008 7142
rect 12058 7032 12114 7041
rect 12058 6967 12114 6976
rect 12072 6322 12100 6967
rect 12164 6866 12192 7375
rect 12532 7177 12560 7890
rect 12624 7342 12652 8026
rect 12612 7336 12664 7342
rect 12612 7278 12664 7284
rect 12518 7168 12574 7177
rect 12518 7103 12574 7112
rect 12532 7002 12560 7103
rect 12520 6996 12572 7002
rect 12520 6938 12572 6944
rect 12152 6860 12204 6866
rect 12152 6802 12204 6808
rect 12060 6316 12112 6322
rect 12060 6258 12112 6264
rect 11888 5914 12008 5930
rect 12072 5914 12100 6258
rect 11876 5908 12008 5914
rect 11928 5902 12008 5908
rect 12060 5908 12112 5914
rect 11876 5850 11928 5856
rect 12060 5850 12112 5856
rect 12164 5846 12192 6802
rect 12336 6792 12388 6798
rect 12336 6734 12388 6740
rect 12152 5840 12204 5846
rect 12152 5782 12204 5788
rect 12244 5568 12296 5574
rect 12244 5510 12296 5516
rect 11784 5160 11836 5166
rect 11784 5102 11836 5108
rect 11796 4826 11824 5102
rect 11968 5092 12020 5098
rect 11968 5034 12020 5040
rect 11784 4820 11836 4826
rect 11784 4762 11836 4768
rect 11980 3777 12008 5034
rect 12150 4040 12206 4049
rect 12150 3975 12152 3984
rect 12204 3975 12206 3984
rect 12152 3946 12204 3952
rect 11966 3768 12022 3777
rect 11966 3703 12022 3712
rect 11600 3528 11652 3534
rect 11600 3470 11652 3476
rect 12060 3528 12112 3534
rect 12060 3470 12112 3476
rect 12072 3058 12100 3470
rect 12256 3194 12284 5510
rect 12348 5234 12376 6734
rect 13072 6180 13124 6186
rect 13072 6122 13124 6128
rect 12336 5228 12388 5234
rect 12336 5170 12388 5176
rect 12348 4826 12376 5170
rect 13084 5098 13112 6122
rect 13176 5710 13204 12396
rect 13348 12378 13400 12384
rect 13360 12102 13388 12378
rect 13452 12345 13480 13806
rect 13438 12336 13494 12345
rect 13438 12271 13494 12280
rect 13440 12232 13492 12238
rect 13440 12174 13492 12180
rect 13348 12096 13400 12102
rect 13348 12038 13400 12044
rect 13452 11354 13480 12174
rect 13440 11348 13492 11354
rect 13440 11290 13492 11296
rect 13254 11248 13310 11257
rect 13254 11183 13310 11192
rect 13268 9625 13296 11183
rect 13452 10810 13480 11290
rect 13440 10804 13492 10810
rect 13440 10746 13492 10752
rect 13452 10606 13480 10746
rect 13440 10600 13492 10606
rect 13346 10568 13402 10577
rect 13440 10542 13492 10548
rect 13346 10503 13402 10512
rect 13360 9874 13388 10503
rect 13544 10130 13572 15302
rect 13636 12986 13664 15438
rect 13716 15360 13768 15366
rect 13716 15302 13768 15308
rect 13728 14958 13756 15302
rect 14484 15260 14780 15280
rect 14540 15258 14564 15260
rect 14620 15258 14644 15260
rect 14700 15258 14724 15260
rect 14562 15206 14564 15258
rect 14626 15206 14638 15258
rect 14700 15206 14702 15258
rect 14540 15204 14564 15206
rect 14620 15204 14644 15206
rect 14700 15204 14724 15206
rect 14484 15184 14780 15204
rect 13716 14952 13768 14958
rect 13716 14894 13768 14900
rect 13728 14074 13756 14894
rect 14174 14784 14230 14793
rect 14174 14719 14230 14728
rect 13808 14476 13860 14482
rect 13808 14418 13860 14424
rect 13716 14068 13768 14074
rect 13716 14010 13768 14016
rect 13820 13977 13848 14418
rect 13806 13968 13862 13977
rect 13728 13912 13806 13920
rect 13728 13892 13808 13912
rect 13624 12980 13676 12986
rect 13624 12922 13676 12928
rect 13636 12238 13664 12922
rect 13728 12594 13756 13892
rect 13860 13903 13862 13912
rect 13808 13874 13860 13880
rect 14084 13320 14136 13326
rect 14084 13262 14136 13268
rect 13808 13184 13860 13190
rect 13808 13126 13860 13132
rect 13820 12782 13848 13126
rect 13990 13016 14046 13025
rect 14096 12986 14124 13262
rect 13990 12951 14046 12960
rect 14084 12980 14136 12986
rect 13808 12776 13860 12782
rect 13808 12718 13860 12724
rect 13728 12566 13848 12594
rect 13820 12442 13848 12566
rect 14004 12442 14032 12951
rect 14084 12922 14136 12928
rect 13808 12436 13860 12442
rect 13808 12378 13860 12384
rect 13992 12436 14044 12442
rect 13992 12378 14044 12384
rect 13624 12232 13676 12238
rect 13624 12174 13676 12180
rect 13636 12073 13664 12174
rect 13622 12064 13678 12073
rect 13622 11999 13678 12008
rect 13636 11898 13664 11999
rect 13624 11892 13676 11898
rect 13624 11834 13676 11840
rect 13636 11218 13664 11834
rect 13898 11792 13954 11801
rect 13898 11727 13954 11736
rect 13716 11620 13768 11626
rect 13716 11562 13768 11568
rect 13624 11212 13676 11218
rect 13624 11154 13676 11160
rect 13532 10124 13584 10130
rect 13532 10066 13584 10072
rect 13438 9888 13494 9897
rect 13360 9846 13438 9874
rect 13438 9823 13494 9832
rect 13254 9616 13310 9625
rect 13254 9551 13310 9560
rect 13348 8968 13400 8974
rect 13346 8936 13348 8945
rect 13400 8936 13402 8945
rect 13346 8871 13402 8880
rect 13452 8634 13480 9823
rect 13544 9722 13572 10066
rect 13532 9716 13584 9722
rect 13532 9658 13584 9664
rect 13728 9518 13756 11562
rect 13912 11354 13940 11727
rect 14004 11626 14032 12378
rect 14096 12102 14124 12922
rect 14084 12096 14136 12102
rect 14084 12038 14136 12044
rect 14096 11830 14124 12038
rect 14188 11898 14216 14719
rect 14924 14550 14952 16594
rect 15660 15978 15688 16730
rect 15740 16652 15792 16658
rect 15740 16594 15792 16600
rect 15752 15978 15780 16594
rect 15648 15972 15700 15978
rect 15648 15914 15700 15920
rect 15740 15972 15792 15978
rect 15740 15914 15792 15920
rect 15372 15496 15424 15502
rect 15372 15438 15424 15444
rect 15004 15360 15056 15366
rect 15004 15302 15056 15308
rect 15016 15026 15044 15302
rect 15004 15020 15056 15026
rect 15004 14962 15056 14968
rect 14912 14544 14964 14550
rect 14964 14492 15044 14498
rect 14912 14486 15044 14492
rect 14924 14470 15044 14486
rect 14360 14408 14412 14414
rect 14360 14350 14412 14356
rect 14912 14408 14964 14414
rect 14912 14350 14964 14356
rect 14268 13932 14320 13938
rect 14268 13874 14320 13880
rect 14280 12986 14308 13874
rect 14372 13394 14400 14350
rect 14484 14172 14780 14192
rect 14540 14170 14564 14172
rect 14620 14170 14644 14172
rect 14700 14170 14724 14172
rect 14562 14118 14564 14170
rect 14626 14118 14638 14170
rect 14700 14118 14702 14170
rect 14540 14116 14564 14118
rect 14620 14116 14644 14118
rect 14700 14116 14724 14118
rect 14484 14096 14780 14116
rect 14820 14000 14872 14006
rect 14820 13942 14872 13948
rect 14832 13870 14860 13942
rect 14820 13864 14872 13870
rect 14820 13806 14872 13812
rect 14924 13530 14952 14350
rect 15016 14074 15044 14470
rect 15004 14068 15056 14074
rect 15004 14010 15056 14016
rect 15384 13802 15412 15438
rect 15752 15162 15780 15914
rect 16212 15706 16240 17070
rect 16568 17060 16620 17066
rect 16568 17002 16620 17008
rect 16580 16726 16608 17002
rect 16568 16720 16620 16726
rect 16568 16662 16620 16668
rect 16580 16250 16608 16662
rect 16660 16584 16712 16590
rect 16660 16526 16712 16532
rect 16844 16584 16896 16590
rect 16844 16526 16896 16532
rect 16568 16244 16620 16250
rect 16568 16186 16620 16192
rect 16672 16114 16700 16526
rect 16856 16153 16884 16526
rect 16842 16144 16898 16153
rect 16660 16108 16712 16114
rect 16842 16079 16898 16088
rect 16660 16050 16712 16056
rect 16752 15904 16804 15910
rect 16752 15846 16804 15852
rect 16200 15700 16252 15706
rect 16200 15642 16252 15648
rect 15924 15632 15976 15638
rect 15924 15574 15976 15580
rect 15740 15156 15792 15162
rect 15740 15098 15792 15104
rect 15936 14822 15964 15574
rect 16016 15496 16068 15502
rect 16016 15438 16068 15444
rect 16028 15178 16056 15438
rect 16028 15162 16148 15178
rect 16028 15156 16160 15162
rect 16028 15150 16108 15156
rect 16108 15098 16160 15104
rect 15924 14816 15976 14822
rect 15924 14758 15976 14764
rect 15372 13796 15424 13802
rect 15372 13738 15424 13744
rect 14912 13524 14964 13530
rect 14912 13466 14964 13472
rect 15096 13524 15148 13530
rect 15096 13466 15148 13472
rect 14360 13388 14412 13394
rect 14360 13330 14412 13336
rect 14484 13084 14780 13104
rect 14540 13082 14564 13084
rect 14620 13082 14644 13084
rect 14700 13082 14724 13084
rect 14562 13030 14564 13082
rect 14626 13030 14638 13082
rect 14700 13030 14702 13082
rect 14540 13028 14564 13030
rect 14620 13028 14644 13030
rect 14700 13028 14724 13030
rect 14484 13008 14780 13028
rect 14268 12980 14320 12986
rect 14268 12922 14320 12928
rect 14360 12776 14412 12782
rect 14360 12718 14412 12724
rect 14266 12200 14322 12209
rect 14266 12135 14322 12144
rect 14176 11892 14228 11898
rect 14176 11834 14228 11840
rect 14084 11824 14136 11830
rect 14084 11766 14136 11772
rect 14280 11762 14308 12135
rect 14268 11756 14320 11762
rect 14268 11698 14320 11704
rect 13992 11620 14044 11626
rect 13992 11562 14044 11568
rect 13900 11348 13952 11354
rect 13900 11290 13952 11296
rect 13912 11082 13940 11290
rect 14372 11286 14400 12718
rect 14912 12708 14964 12714
rect 14912 12650 14964 12656
rect 14542 12200 14598 12209
rect 14542 12135 14544 12144
rect 14596 12135 14598 12144
rect 14544 12106 14596 12112
rect 14484 11996 14780 12016
rect 14540 11994 14564 11996
rect 14620 11994 14644 11996
rect 14700 11994 14724 11996
rect 14562 11942 14564 11994
rect 14626 11942 14638 11994
rect 14700 11942 14702 11994
rect 14540 11940 14564 11942
rect 14620 11940 14644 11942
rect 14700 11940 14724 11942
rect 14484 11920 14780 11940
rect 14360 11280 14412 11286
rect 14360 11222 14412 11228
rect 13900 11076 13952 11082
rect 13900 11018 13952 11024
rect 13806 10840 13862 10849
rect 13806 10775 13808 10784
rect 13860 10775 13862 10784
rect 13808 10746 13860 10752
rect 13912 10742 13940 11018
rect 14176 10804 14228 10810
rect 14176 10746 14228 10752
rect 13900 10736 13952 10742
rect 13900 10678 13952 10684
rect 14188 10266 14216 10746
rect 14372 10266 14400 11222
rect 14924 11014 14952 12650
rect 15004 11824 15056 11830
rect 15004 11766 15056 11772
rect 15016 11665 15044 11766
rect 15002 11656 15058 11665
rect 15002 11591 15004 11600
rect 15056 11591 15058 11600
rect 15004 11562 15056 11568
rect 15016 11354 15044 11562
rect 15004 11348 15056 11354
rect 15004 11290 15056 11296
rect 14912 11008 14964 11014
rect 14912 10950 14964 10956
rect 14484 10908 14780 10928
rect 14540 10906 14564 10908
rect 14620 10906 14644 10908
rect 14700 10906 14724 10908
rect 14562 10854 14564 10906
rect 14626 10854 14638 10906
rect 14700 10854 14702 10906
rect 14540 10852 14564 10854
rect 14620 10852 14644 10854
rect 14700 10852 14724 10854
rect 14484 10832 14780 10852
rect 14924 10810 14952 10950
rect 14912 10804 14964 10810
rect 14964 10764 15044 10792
rect 14912 10746 14964 10752
rect 14636 10464 14688 10470
rect 14636 10406 14688 10412
rect 14648 10305 14676 10406
rect 14634 10296 14690 10305
rect 14176 10260 14228 10266
rect 14176 10202 14228 10208
rect 14360 10260 14412 10266
rect 14634 10231 14690 10240
rect 14360 10202 14412 10208
rect 13990 10160 14046 10169
rect 13990 10095 13992 10104
rect 14044 10095 14046 10104
rect 14912 10124 14964 10130
rect 13992 10066 14044 10072
rect 14912 10066 14964 10072
rect 14924 10010 14952 10066
rect 13900 9988 13952 9994
rect 13900 9930 13952 9936
rect 14832 9982 14952 10010
rect 13808 9920 13860 9926
rect 13808 9862 13860 9868
rect 13716 9512 13768 9518
rect 13716 9454 13768 9460
rect 13728 9042 13756 9454
rect 13820 9450 13848 9862
rect 13912 9466 13940 9930
rect 14484 9820 14780 9840
rect 14540 9818 14564 9820
rect 14620 9818 14644 9820
rect 14700 9818 14724 9820
rect 14562 9766 14564 9818
rect 14626 9766 14638 9818
rect 14700 9766 14702 9818
rect 14540 9764 14564 9766
rect 14620 9764 14644 9766
rect 14700 9764 14724 9766
rect 14484 9744 14780 9764
rect 14832 9602 14860 9982
rect 14912 9920 14964 9926
rect 14912 9862 14964 9868
rect 14924 9722 14952 9862
rect 15016 9722 15044 10764
rect 14912 9716 14964 9722
rect 14912 9658 14964 9664
rect 15004 9716 15056 9722
rect 15004 9658 15056 9664
rect 14648 9574 14860 9602
rect 13992 9512 14044 9518
rect 13912 9460 13992 9466
rect 13912 9454 14044 9460
rect 13808 9444 13860 9450
rect 13808 9386 13860 9392
rect 13912 9438 14032 9454
rect 13716 9036 13768 9042
rect 13716 8978 13768 8984
rect 13820 8974 13848 9386
rect 13808 8968 13860 8974
rect 13808 8910 13860 8916
rect 13440 8628 13492 8634
rect 13440 8570 13492 8576
rect 13452 8430 13480 8570
rect 13820 8430 13848 8910
rect 13912 8838 13940 9438
rect 14648 9178 14676 9574
rect 14728 9376 14780 9382
rect 14728 9318 14780 9324
rect 14636 9172 14688 9178
rect 14636 9114 14688 9120
rect 14740 8922 14768 9318
rect 15004 9104 15056 9110
rect 15004 9046 15056 9052
rect 14912 9036 14964 9042
rect 14912 8978 14964 8984
rect 14740 8894 14860 8922
rect 13900 8832 13952 8838
rect 13900 8774 13952 8780
rect 13440 8424 13492 8430
rect 13440 8366 13492 8372
rect 13808 8424 13860 8430
rect 13808 8366 13860 8372
rect 13256 7948 13308 7954
rect 13256 7890 13308 7896
rect 13268 7546 13296 7890
rect 13452 7546 13480 8366
rect 13820 8090 13848 8366
rect 13912 8362 13940 8774
rect 14484 8732 14780 8752
rect 14540 8730 14564 8732
rect 14620 8730 14644 8732
rect 14700 8730 14724 8732
rect 14562 8678 14564 8730
rect 14626 8678 14638 8730
rect 14700 8678 14702 8730
rect 14540 8676 14564 8678
rect 14620 8676 14644 8678
rect 14700 8676 14724 8678
rect 14484 8656 14780 8676
rect 14268 8560 14320 8566
rect 14268 8502 14320 8508
rect 13900 8356 13952 8362
rect 13900 8298 13952 8304
rect 13912 8265 13940 8298
rect 13898 8256 13954 8265
rect 13898 8191 13954 8200
rect 13808 8084 13860 8090
rect 13808 8026 13860 8032
rect 13900 7880 13952 7886
rect 13900 7822 13952 7828
rect 13256 7540 13308 7546
rect 13256 7482 13308 7488
rect 13440 7540 13492 7546
rect 13440 7482 13492 7488
rect 13912 7449 13940 7822
rect 13898 7440 13954 7449
rect 13898 7375 13954 7384
rect 13348 6928 13400 6934
rect 13346 6896 13348 6905
rect 13400 6896 13402 6905
rect 13346 6831 13402 6840
rect 13256 6792 13308 6798
rect 13256 6734 13308 6740
rect 13268 6497 13296 6734
rect 13254 6488 13310 6497
rect 13254 6423 13256 6432
rect 13308 6423 13310 6432
rect 13256 6394 13308 6400
rect 13268 6363 13296 6394
rect 13360 6322 13388 6831
rect 14280 6322 14308 8502
rect 14634 8256 14690 8265
rect 14634 8191 14690 8200
rect 14360 8084 14412 8090
rect 14360 8026 14412 8032
rect 14372 7886 14400 8026
rect 14648 7954 14676 8191
rect 14832 7954 14860 8894
rect 14924 8090 14952 8978
rect 15016 8634 15044 9046
rect 15108 8945 15136 13466
rect 15936 13462 15964 14758
rect 16016 14612 16068 14618
rect 16016 14554 16068 14560
rect 16028 13530 16056 14554
rect 16660 14476 16712 14482
rect 16660 14418 16712 14424
rect 16384 14068 16436 14074
rect 16384 14010 16436 14016
rect 16396 13977 16424 14010
rect 16672 14006 16700 14418
rect 16660 14000 16712 14006
rect 16382 13968 16438 13977
rect 16382 13903 16438 13912
rect 16488 13960 16660 13988
rect 16488 13818 16516 13960
rect 16660 13942 16712 13948
rect 16396 13790 16516 13818
rect 16016 13524 16068 13530
rect 16016 13466 16068 13472
rect 15924 13456 15976 13462
rect 15924 13398 15976 13404
rect 16028 12850 16056 13466
rect 16292 13456 16344 13462
rect 16292 13398 16344 13404
rect 16108 13388 16160 13394
rect 16108 13330 16160 13336
rect 16016 12844 16068 12850
rect 16016 12786 16068 12792
rect 16120 12442 16148 13330
rect 16304 12714 16332 13398
rect 16292 12708 16344 12714
rect 16292 12650 16344 12656
rect 16108 12436 16160 12442
rect 16108 12378 16160 12384
rect 15186 12336 15242 12345
rect 15186 12271 15242 12280
rect 15200 11898 15228 12271
rect 15740 12232 15792 12238
rect 15740 12174 15792 12180
rect 15188 11892 15240 11898
rect 15188 11834 15240 11840
rect 15200 11694 15228 11834
rect 15188 11688 15240 11694
rect 15188 11630 15240 11636
rect 15280 11620 15332 11626
rect 15280 11562 15332 11568
rect 15188 11144 15240 11150
rect 15188 11086 15240 11092
rect 15200 10674 15228 11086
rect 15292 11014 15320 11562
rect 15464 11552 15516 11558
rect 15464 11494 15516 11500
rect 15280 11008 15332 11014
rect 15280 10950 15332 10956
rect 15188 10668 15240 10674
rect 15188 10610 15240 10616
rect 15292 10130 15320 10950
rect 15372 10464 15424 10470
rect 15372 10406 15424 10412
rect 15384 10169 15412 10406
rect 15370 10160 15426 10169
rect 15280 10124 15332 10130
rect 15370 10095 15426 10104
rect 15280 10066 15332 10072
rect 15094 8936 15150 8945
rect 15094 8871 15150 8880
rect 15004 8628 15056 8634
rect 15004 8570 15056 8576
rect 15372 8356 15424 8362
rect 15372 8298 15424 8304
rect 14912 8084 14964 8090
rect 14912 8026 14964 8032
rect 14636 7948 14688 7954
rect 14636 7890 14688 7896
rect 14820 7948 14872 7954
rect 14820 7890 14872 7896
rect 14360 7880 14412 7886
rect 14360 7822 14412 7828
rect 14372 7342 14400 7822
rect 14484 7644 14780 7664
rect 14540 7642 14564 7644
rect 14620 7642 14644 7644
rect 14700 7642 14724 7644
rect 14562 7590 14564 7642
rect 14626 7590 14638 7642
rect 14700 7590 14702 7642
rect 14540 7588 14564 7590
rect 14620 7588 14644 7590
rect 14700 7588 14724 7590
rect 14484 7568 14780 7588
rect 14636 7472 14688 7478
rect 14636 7414 14688 7420
rect 14360 7336 14412 7342
rect 14360 7278 14412 7284
rect 14372 7002 14400 7278
rect 14360 6996 14412 7002
rect 14360 6938 14412 6944
rect 14648 6746 14676 7414
rect 14832 7002 14860 7890
rect 14924 7342 14952 8026
rect 15384 8022 15412 8298
rect 15372 8016 15424 8022
rect 15372 7958 15424 7964
rect 15384 7546 15412 7958
rect 15372 7540 15424 7546
rect 15372 7482 15424 7488
rect 14912 7336 14964 7342
rect 14912 7278 14964 7284
rect 14820 6996 14872 7002
rect 14820 6938 14872 6944
rect 14648 6718 14860 6746
rect 14484 6556 14780 6576
rect 14540 6554 14564 6556
rect 14620 6554 14644 6556
rect 14700 6554 14724 6556
rect 14562 6502 14564 6554
rect 14626 6502 14638 6554
rect 14700 6502 14702 6554
rect 14540 6500 14564 6502
rect 14620 6500 14644 6502
rect 14700 6500 14724 6502
rect 14484 6480 14780 6500
rect 13348 6316 13400 6322
rect 13348 6258 13400 6264
rect 14268 6316 14320 6322
rect 14268 6258 14320 6264
rect 13256 6112 13308 6118
rect 13256 6054 13308 6060
rect 13268 5846 13296 6054
rect 14280 5914 14308 6258
rect 14268 5908 14320 5914
rect 14268 5850 14320 5856
rect 13256 5840 13308 5846
rect 13256 5782 13308 5788
rect 13164 5704 13216 5710
rect 13164 5646 13216 5652
rect 13072 5092 13124 5098
rect 13072 5034 13124 5040
rect 13176 4826 13204 5646
rect 13268 5098 13296 5782
rect 14832 5778 14860 6718
rect 15096 6656 15148 6662
rect 15096 6598 15148 6604
rect 14360 5772 14412 5778
rect 14360 5714 14412 5720
rect 14820 5772 14872 5778
rect 14820 5714 14872 5720
rect 13348 5704 13400 5710
rect 13348 5646 13400 5652
rect 13256 5092 13308 5098
rect 13256 5034 13308 5040
rect 12336 4820 12388 4826
rect 12336 4762 12388 4768
rect 13164 4820 13216 4826
rect 13164 4762 13216 4768
rect 13256 4616 13308 4622
rect 12426 4584 12482 4593
rect 13256 4558 13308 4564
rect 12426 4519 12482 4528
rect 12440 4146 12468 4519
rect 12428 4140 12480 4146
rect 12428 4082 12480 4088
rect 12440 3738 12468 4082
rect 12428 3732 12480 3738
rect 12428 3674 12480 3680
rect 13268 3505 13296 4558
rect 13360 4146 13388 5646
rect 14372 5370 14400 5714
rect 14484 5468 14780 5488
rect 14540 5466 14564 5468
rect 14620 5466 14644 5468
rect 14700 5466 14724 5468
rect 14562 5414 14564 5466
rect 14626 5414 14638 5466
rect 14700 5414 14702 5466
rect 14540 5412 14564 5414
rect 14620 5412 14644 5414
rect 14700 5412 14724 5414
rect 14484 5392 14780 5412
rect 14360 5364 14412 5370
rect 14360 5306 14412 5312
rect 14636 5092 14688 5098
rect 14636 5034 14688 5040
rect 13532 5024 13584 5030
rect 13532 4966 13584 4972
rect 13716 5024 13768 5030
rect 13716 4966 13768 4972
rect 13440 4752 13492 4758
rect 13440 4694 13492 4700
rect 13452 4282 13480 4694
rect 13440 4276 13492 4282
rect 13440 4218 13492 4224
rect 13348 4140 13400 4146
rect 13348 4082 13400 4088
rect 13544 3942 13572 4966
rect 13728 4321 13756 4966
rect 14266 4856 14322 4865
rect 14266 4791 14322 4800
rect 13900 4616 13952 4622
rect 13900 4558 13952 4564
rect 13714 4312 13770 4321
rect 13714 4247 13770 4256
rect 13532 3936 13584 3942
rect 13532 3878 13584 3884
rect 13544 3602 13572 3878
rect 13532 3596 13584 3602
rect 13532 3538 13584 3544
rect 13254 3496 13310 3505
rect 13254 3431 13310 3440
rect 13162 3360 13218 3369
rect 13162 3295 13218 3304
rect 12334 3224 12390 3233
rect 12244 3188 12296 3194
rect 13176 3194 13204 3295
rect 12334 3159 12390 3168
rect 12428 3188 12480 3194
rect 12244 3130 12296 3136
rect 12348 3058 12376 3159
rect 12428 3130 12480 3136
rect 13164 3188 13216 3194
rect 13164 3130 13216 3136
rect 12060 3052 12112 3058
rect 12060 2994 12112 3000
rect 12336 3052 12388 3058
rect 12336 2994 12388 3000
rect 11324 2848 11376 2854
rect 11324 2790 11376 2796
rect 12242 2816 12298 2825
rect 11336 2650 11364 2790
rect 12242 2751 12298 2760
rect 11324 2644 11376 2650
rect 11324 2586 11376 2592
rect 10496 2440 10548 2446
rect 11508 2440 11560 2446
rect 10496 2382 10548 2388
rect 11506 2408 11508 2417
rect 11560 2408 11562 2417
rect 11506 2343 11562 2352
rect 10312 2304 10364 2310
rect 10312 2246 10364 2252
rect 11322 2272 11378 2281
rect 10324 480 10352 2246
rect 12256 2258 12284 2751
rect 12348 2446 12376 2994
rect 12440 2922 12468 3130
rect 13438 3088 13494 3097
rect 13438 3023 13494 3032
rect 12428 2916 12480 2922
rect 12428 2858 12480 2864
rect 12440 2825 12468 2858
rect 12426 2816 12482 2825
rect 12426 2751 12482 2760
rect 12336 2440 12388 2446
rect 12336 2382 12388 2388
rect 12256 2230 12468 2258
rect 11322 2207 11378 2216
rect 11336 480 11364 2207
rect 12440 480 12468 2230
rect 13452 480 13480 3023
rect 13544 2650 13572 3538
rect 13912 3534 13940 4558
rect 14280 4146 14308 4791
rect 14648 4758 14676 5034
rect 14636 4752 14688 4758
rect 14636 4694 14688 4700
rect 15108 4690 15136 6598
rect 15280 6384 15332 6390
rect 15280 6326 15332 6332
rect 15188 6180 15240 6186
rect 15188 6122 15240 6128
rect 15200 5846 15228 6122
rect 15188 5840 15240 5846
rect 15188 5782 15240 5788
rect 15200 5234 15228 5782
rect 15188 5228 15240 5234
rect 15188 5170 15240 5176
rect 15292 5166 15320 6326
rect 15476 5681 15504 11494
rect 15554 9888 15610 9897
rect 15554 9823 15610 9832
rect 15568 9110 15596 9823
rect 15556 9104 15608 9110
rect 15556 9046 15608 9052
rect 15648 8900 15700 8906
rect 15648 8842 15700 8848
rect 15660 8498 15688 8842
rect 15752 8634 15780 12174
rect 15832 12096 15884 12102
rect 15832 12038 15884 12044
rect 15844 11694 15872 12038
rect 15832 11688 15884 11694
rect 15832 11630 15884 11636
rect 16200 11144 16252 11150
rect 16200 11086 16252 11092
rect 16108 11076 16160 11082
rect 16108 11018 16160 11024
rect 16120 10810 16148 11018
rect 16108 10804 16160 10810
rect 16108 10746 16160 10752
rect 16212 10305 16240 11086
rect 16198 10296 16254 10305
rect 16198 10231 16200 10240
rect 16252 10231 16254 10240
rect 16200 10202 16252 10208
rect 16304 10198 16332 12650
rect 16396 11218 16424 13790
rect 16476 13728 16528 13734
rect 16476 13670 16528 13676
rect 16488 13433 16516 13670
rect 16474 13424 16530 13433
rect 16474 13359 16530 13368
rect 16660 12640 16712 12646
rect 16660 12582 16712 12588
rect 16672 12481 16700 12582
rect 16658 12472 16714 12481
rect 16658 12407 16660 12416
rect 16712 12407 16714 12416
rect 16660 12378 16712 12384
rect 16764 12374 16792 15846
rect 16856 15434 16884 16079
rect 17396 16040 17448 16046
rect 17396 15982 17448 15988
rect 17120 15972 17172 15978
rect 17120 15914 17172 15920
rect 17028 15700 17080 15706
rect 17028 15642 17080 15648
rect 16844 15428 16896 15434
rect 16844 15370 16896 15376
rect 17040 15162 17068 15642
rect 17132 15502 17160 15914
rect 17120 15496 17172 15502
rect 17120 15438 17172 15444
rect 17028 15156 17080 15162
rect 17028 15098 17080 15104
rect 16936 14816 16988 14822
rect 16936 14758 16988 14764
rect 16844 14476 16896 14482
rect 16844 14418 16896 14424
rect 16856 14074 16884 14418
rect 16844 14068 16896 14074
rect 16844 14010 16896 14016
rect 16948 12986 16976 14758
rect 17132 14550 17160 15438
rect 17120 14544 17172 14550
rect 17120 14486 17172 14492
rect 17408 14074 17436 15982
rect 17868 14618 17896 17303
rect 18684 16788 18736 16794
rect 18684 16730 18736 16736
rect 18224 16652 18276 16658
rect 18224 16594 18276 16600
rect 18236 15910 18264 16594
rect 18224 15904 18276 15910
rect 18224 15846 18276 15852
rect 18038 15328 18094 15337
rect 18038 15263 18094 15272
rect 17948 14816 18000 14822
rect 17946 14784 17948 14793
rect 18000 14784 18002 14793
rect 17946 14719 18002 14728
rect 17856 14612 17908 14618
rect 17856 14554 17908 14560
rect 17396 14068 17448 14074
rect 17396 14010 17448 14016
rect 17408 13734 17436 14010
rect 17868 13818 17896 14554
rect 17948 13932 18000 13938
rect 17948 13874 18000 13880
rect 17684 13802 17896 13818
rect 17672 13796 17896 13802
rect 17724 13790 17896 13796
rect 17672 13738 17724 13744
rect 17396 13728 17448 13734
rect 17316 13688 17396 13716
rect 17316 13530 17344 13688
rect 17396 13670 17448 13676
rect 17960 13530 17988 13874
rect 17304 13524 17356 13530
rect 17304 13466 17356 13472
rect 17948 13524 18000 13530
rect 17948 13466 18000 13472
rect 17028 13456 17080 13462
rect 17028 13398 17080 13404
rect 17580 13456 17632 13462
rect 17580 13398 17632 13404
rect 16936 12980 16988 12986
rect 16936 12922 16988 12928
rect 17040 12374 17068 13398
rect 17304 12912 17356 12918
rect 17302 12880 17304 12889
rect 17356 12880 17358 12889
rect 17302 12815 17358 12824
rect 17316 12714 17344 12815
rect 17304 12708 17356 12714
rect 17304 12650 17356 12656
rect 17592 12646 17620 13398
rect 17948 13252 18000 13258
rect 17948 13194 18000 13200
rect 17960 12850 17988 13194
rect 17948 12844 18000 12850
rect 17948 12786 18000 12792
rect 17960 12753 17988 12786
rect 17946 12744 18002 12753
rect 17946 12679 18002 12688
rect 17580 12640 17632 12646
rect 17580 12582 17632 12588
rect 18052 12458 18080 15263
rect 18592 14952 18644 14958
rect 18592 14894 18644 14900
rect 18604 14618 18632 14894
rect 18592 14612 18644 14618
rect 18592 14554 18644 14560
rect 18604 13376 18632 14554
rect 18512 13348 18632 13376
rect 18512 12782 18540 13348
rect 18500 12776 18552 12782
rect 18314 12744 18370 12753
rect 18500 12718 18552 12724
rect 18314 12679 18370 12688
rect 17776 12430 18080 12458
rect 16752 12368 16804 12374
rect 16752 12310 16804 12316
rect 17028 12368 17080 12374
rect 17028 12310 17080 12316
rect 17578 12336 17634 12345
rect 16660 12232 16712 12238
rect 16660 12174 16712 12180
rect 16672 11778 16700 12174
rect 16764 11898 16792 12310
rect 17578 12271 17634 12280
rect 17302 12200 17358 12209
rect 17302 12135 17358 12144
rect 17316 12102 17344 12135
rect 17304 12096 17356 12102
rect 17304 12038 17356 12044
rect 17316 11898 17344 12038
rect 16752 11892 16804 11898
rect 16752 11834 16804 11840
rect 17304 11892 17356 11898
rect 17304 11834 17356 11840
rect 16672 11750 16792 11778
rect 16764 11558 16792 11750
rect 16752 11552 16804 11558
rect 16750 11520 16752 11529
rect 16804 11520 16806 11529
rect 16750 11455 16806 11464
rect 16476 11348 16528 11354
rect 16476 11290 16528 11296
rect 16384 11212 16436 11218
rect 16384 11154 16436 11160
rect 16292 10192 16344 10198
rect 16292 10134 16344 10140
rect 16488 10130 16516 11290
rect 16660 11212 16712 11218
rect 16660 11154 16712 11160
rect 17488 11212 17540 11218
rect 17488 11154 17540 11160
rect 16672 10470 16700 11154
rect 17304 10804 17356 10810
rect 17304 10746 17356 10752
rect 17210 10568 17266 10577
rect 17210 10503 17212 10512
rect 17264 10503 17266 10512
rect 17212 10474 17264 10480
rect 16660 10464 16712 10470
rect 16660 10406 16712 10412
rect 16936 10464 16988 10470
rect 16936 10406 16988 10412
rect 16752 10192 16804 10198
rect 16752 10134 16804 10140
rect 16476 10124 16528 10130
rect 16476 10066 16528 10072
rect 16016 10056 16068 10062
rect 16016 9998 16068 10004
rect 15832 9920 15884 9926
rect 15832 9862 15884 9868
rect 15844 9450 15872 9862
rect 15924 9648 15976 9654
rect 15924 9590 15976 9596
rect 15832 9444 15884 9450
rect 15832 9386 15884 9392
rect 15740 8628 15792 8634
rect 15740 8570 15792 8576
rect 15648 8492 15700 8498
rect 15648 8434 15700 8440
rect 15844 8090 15872 9386
rect 15832 8084 15884 8090
rect 15832 8026 15884 8032
rect 15844 7546 15872 8026
rect 15832 7540 15884 7546
rect 15832 7482 15884 7488
rect 15844 7342 15872 7482
rect 15832 7336 15884 7342
rect 15832 7278 15884 7284
rect 15936 7018 15964 9590
rect 16028 8616 16056 9998
rect 16488 9178 16516 10066
rect 16764 9382 16792 10134
rect 16948 9994 16976 10406
rect 16936 9988 16988 9994
rect 16936 9930 16988 9936
rect 17316 9722 17344 10746
rect 17500 10538 17528 11154
rect 17592 10606 17620 12271
rect 17670 11792 17726 11801
rect 17670 11727 17726 11736
rect 17684 11694 17712 11727
rect 17672 11688 17724 11694
rect 17672 11630 17724 11636
rect 17684 11286 17712 11630
rect 17672 11280 17724 11286
rect 17672 11222 17724 11228
rect 17580 10600 17632 10606
rect 17580 10542 17632 10548
rect 17488 10532 17540 10538
rect 17488 10474 17540 10480
rect 17592 10266 17620 10542
rect 17580 10260 17632 10266
rect 17580 10202 17632 10208
rect 17396 9920 17448 9926
rect 17396 9862 17448 9868
rect 17304 9716 17356 9722
rect 17304 9658 17356 9664
rect 16844 9580 16896 9586
rect 16844 9522 16896 9528
rect 16752 9376 16804 9382
rect 16752 9318 16804 9324
rect 16476 9172 16528 9178
rect 16476 9114 16528 9120
rect 16028 8588 16240 8616
rect 16108 8492 16160 8498
rect 16108 8434 16160 8440
rect 16120 8090 16148 8434
rect 16108 8084 16160 8090
rect 16108 8026 16160 8032
rect 16212 7954 16240 8588
rect 16384 8424 16436 8430
rect 16384 8366 16436 8372
rect 16200 7948 16252 7954
rect 16200 7890 16252 7896
rect 16108 7200 16160 7206
rect 16108 7142 16160 7148
rect 15936 6990 16056 7018
rect 15740 6860 15792 6866
rect 15740 6802 15792 6808
rect 15752 6662 15780 6802
rect 16028 6798 16056 6990
rect 16120 6905 16148 7142
rect 16106 6896 16162 6905
rect 16396 6866 16424 8366
rect 16764 8362 16792 9318
rect 16856 9110 16884 9522
rect 17408 9450 17436 9862
rect 17670 9616 17726 9625
rect 17670 9551 17672 9560
rect 17724 9551 17726 9560
rect 17672 9522 17724 9528
rect 17396 9444 17448 9450
rect 17396 9386 17448 9392
rect 16844 9104 16896 9110
rect 16842 9072 16844 9081
rect 17580 9104 17632 9110
rect 16896 9072 16898 9081
rect 17580 9046 17632 9052
rect 16842 9007 16898 9016
rect 16936 8968 16988 8974
rect 16936 8910 16988 8916
rect 16948 8634 16976 8910
rect 16936 8628 16988 8634
rect 16936 8570 16988 8576
rect 17592 8498 17620 9046
rect 17684 8906 17712 9522
rect 17672 8900 17724 8906
rect 17672 8842 17724 8848
rect 17580 8492 17632 8498
rect 17580 8434 17632 8440
rect 16752 8356 16804 8362
rect 17776 8344 17804 12430
rect 18328 12306 18356 12679
rect 18512 12345 18540 12718
rect 18498 12336 18554 12345
rect 18132 12300 18184 12306
rect 18132 12242 18184 12248
rect 18316 12300 18368 12306
rect 18498 12271 18554 12280
rect 18316 12242 18368 12248
rect 18040 12164 18092 12170
rect 18040 12106 18092 12112
rect 18052 11762 18080 12106
rect 18040 11756 18092 11762
rect 18040 11698 18092 11704
rect 18144 11218 18172 12242
rect 18328 12158 18632 12186
rect 18224 12096 18276 12102
rect 18328 12084 18356 12158
rect 18604 12102 18632 12158
rect 18276 12056 18356 12084
rect 18592 12096 18644 12102
rect 18224 12038 18276 12044
rect 18592 12038 18644 12044
rect 18236 11665 18264 12038
rect 18696 11898 18724 16730
rect 18788 16402 18816 27520
rect 19150 25596 19446 25616
rect 19206 25594 19230 25596
rect 19286 25594 19310 25596
rect 19366 25594 19390 25596
rect 19228 25542 19230 25594
rect 19292 25542 19304 25594
rect 19366 25542 19368 25594
rect 19206 25540 19230 25542
rect 19286 25540 19310 25542
rect 19366 25540 19390 25542
rect 19150 25520 19446 25540
rect 19150 24508 19446 24528
rect 19206 24506 19230 24508
rect 19286 24506 19310 24508
rect 19366 24506 19390 24508
rect 19228 24454 19230 24506
rect 19292 24454 19304 24506
rect 19366 24454 19368 24506
rect 19206 24452 19230 24454
rect 19286 24452 19310 24454
rect 19366 24452 19390 24454
rect 19150 24432 19446 24452
rect 20890 23624 20946 23633
rect 20890 23559 20946 23568
rect 20340 23520 20392 23526
rect 20340 23462 20392 23468
rect 19150 23420 19446 23440
rect 19206 23418 19230 23420
rect 19286 23418 19310 23420
rect 19366 23418 19390 23420
rect 19228 23366 19230 23418
rect 19292 23366 19304 23418
rect 19366 23366 19368 23418
rect 19206 23364 19230 23366
rect 19286 23364 19310 23366
rect 19366 23364 19390 23366
rect 19150 23344 19446 23364
rect 19150 22332 19446 22352
rect 19206 22330 19230 22332
rect 19286 22330 19310 22332
rect 19366 22330 19390 22332
rect 19228 22278 19230 22330
rect 19292 22278 19304 22330
rect 19366 22278 19368 22330
rect 19206 22276 19230 22278
rect 19286 22276 19310 22278
rect 19366 22276 19390 22278
rect 19150 22256 19446 22276
rect 19150 21244 19446 21264
rect 19206 21242 19230 21244
rect 19286 21242 19310 21244
rect 19366 21242 19390 21244
rect 19228 21190 19230 21242
rect 19292 21190 19304 21242
rect 19366 21190 19368 21242
rect 19206 21188 19230 21190
rect 19286 21188 19310 21190
rect 19366 21188 19390 21190
rect 19150 21168 19446 21188
rect 19150 20156 19446 20176
rect 19206 20154 19230 20156
rect 19286 20154 19310 20156
rect 19366 20154 19390 20156
rect 19228 20102 19230 20154
rect 19292 20102 19304 20154
rect 19366 20102 19368 20154
rect 19206 20100 19230 20102
rect 19286 20100 19310 20102
rect 19366 20100 19390 20102
rect 19150 20080 19446 20100
rect 19150 19068 19446 19088
rect 19206 19066 19230 19068
rect 19286 19066 19310 19068
rect 19366 19066 19390 19068
rect 19228 19014 19230 19066
rect 19292 19014 19304 19066
rect 19366 19014 19368 19066
rect 19206 19012 19230 19014
rect 19286 19012 19310 19014
rect 19366 19012 19390 19014
rect 19150 18992 19446 19012
rect 19150 17980 19446 18000
rect 19206 17978 19230 17980
rect 19286 17978 19310 17980
rect 19366 17978 19390 17980
rect 19228 17926 19230 17978
rect 19292 17926 19304 17978
rect 19366 17926 19368 17978
rect 19206 17924 19230 17926
rect 19286 17924 19310 17926
rect 19366 17924 19390 17926
rect 19150 17904 19446 17924
rect 19972 17128 20024 17134
rect 19972 17070 20024 17076
rect 19150 16892 19446 16912
rect 19206 16890 19230 16892
rect 19286 16890 19310 16892
rect 19366 16890 19390 16892
rect 19228 16838 19230 16890
rect 19292 16838 19304 16890
rect 19366 16838 19368 16890
rect 19206 16836 19230 16838
rect 19286 16836 19310 16838
rect 19366 16836 19390 16838
rect 19150 16816 19446 16836
rect 19512 16448 19564 16454
rect 18788 16374 19000 16402
rect 19512 16390 19564 16396
rect 18776 15904 18828 15910
rect 18776 15846 18828 15852
rect 18788 13512 18816 15846
rect 18972 15609 19000 16374
rect 19524 16046 19552 16390
rect 19512 16040 19564 16046
rect 19512 15982 19564 15988
rect 19150 15804 19446 15824
rect 19206 15802 19230 15804
rect 19286 15802 19310 15804
rect 19366 15802 19390 15804
rect 19228 15750 19230 15802
rect 19292 15750 19304 15802
rect 19366 15750 19368 15802
rect 19206 15748 19230 15750
rect 19286 15748 19310 15750
rect 19366 15748 19390 15750
rect 19150 15728 19446 15748
rect 18958 15600 19014 15609
rect 18958 15535 19014 15544
rect 19052 15564 19104 15570
rect 18868 13524 18920 13530
rect 18788 13484 18868 13512
rect 18788 12170 18816 13484
rect 18868 13466 18920 13472
rect 18972 13394 19000 15535
rect 19052 15506 19104 15512
rect 19144 15564 19196 15570
rect 19144 15506 19196 15512
rect 19064 14822 19092 15506
rect 19156 14958 19184 15506
rect 19524 15026 19552 15982
rect 19512 15020 19564 15026
rect 19512 14962 19564 14968
rect 19144 14952 19196 14958
rect 19144 14894 19196 14900
rect 19984 14890 20012 17070
rect 20156 16992 20208 16998
rect 20156 16934 20208 16940
rect 20064 15496 20116 15502
rect 20064 15438 20116 15444
rect 20076 15162 20104 15438
rect 20064 15156 20116 15162
rect 20064 15098 20116 15104
rect 19972 14884 20024 14890
rect 19972 14826 20024 14832
rect 19052 14816 19104 14822
rect 19052 14758 19104 14764
rect 19064 14482 19092 14758
rect 19150 14716 19446 14736
rect 19206 14714 19230 14716
rect 19286 14714 19310 14716
rect 19366 14714 19390 14716
rect 19228 14662 19230 14714
rect 19292 14662 19304 14714
rect 19366 14662 19368 14714
rect 19206 14660 19230 14662
rect 19286 14660 19310 14662
rect 19366 14660 19390 14662
rect 19150 14640 19446 14660
rect 19052 14476 19104 14482
rect 19052 14418 19104 14424
rect 19696 14476 19748 14482
rect 19696 14418 19748 14424
rect 19064 14074 19092 14418
rect 19052 14068 19104 14074
rect 19052 14010 19104 14016
rect 19150 13628 19446 13648
rect 19206 13626 19230 13628
rect 19286 13626 19310 13628
rect 19366 13626 19390 13628
rect 19228 13574 19230 13626
rect 19292 13574 19304 13626
rect 19366 13574 19368 13626
rect 19206 13572 19230 13574
rect 19286 13572 19310 13574
rect 19366 13572 19390 13574
rect 19150 13552 19446 13572
rect 19602 13560 19658 13569
rect 19602 13495 19658 13504
rect 19616 13462 19644 13495
rect 19604 13456 19656 13462
rect 19604 13398 19656 13404
rect 18960 13388 19012 13394
rect 18960 13330 19012 13336
rect 18972 12986 19000 13330
rect 18960 12980 19012 12986
rect 18960 12922 19012 12928
rect 19512 12776 19564 12782
rect 19512 12718 19564 12724
rect 18958 12608 19014 12617
rect 18958 12543 19014 12552
rect 18972 12374 19000 12543
rect 19150 12540 19446 12560
rect 19206 12538 19230 12540
rect 19286 12538 19310 12540
rect 19366 12538 19390 12540
rect 19228 12486 19230 12538
rect 19292 12486 19304 12538
rect 19366 12486 19368 12538
rect 19206 12484 19230 12486
rect 19286 12484 19310 12486
rect 19366 12484 19390 12486
rect 19150 12464 19446 12484
rect 19524 12442 19552 12718
rect 19512 12436 19564 12442
rect 19512 12378 19564 12384
rect 19616 12374 19644 13398
rect 19708 13190 19736 14418
rect 19788 14272 19840 14278
rect 19788 14214 19840 14220
rect 19800 13938 19828 14214
rect 19788 13932 19840 13938
rect 19788 13874 19840 13880
rect 19696 13184 19748 13190
rect 19696 13126 19748 13132
rect 19708 12782 19736 13126
rect 19800 12850 19828 13874
rect 20168 13462 20196 16934
rect 20248 16584 20300 16590
rect 20248 16526 20300 16532
rect 20260 15473 20288 16526
rect 20246 15464 20302 15473
rect 20246 15399 20248 15408
rect 20300 15399 20302 15408
rect 20248 15370 20300 15376
rect 20352 15026 20380 23462
rect 20798 20768 20854 20777
rect 20798 20703 20854 20712
rect 20522 20088 20578 20097
rect 20522 20023 20578 20032
rect 20536 18834 20564 20023
rect 20524 18828 20576 18834
rect 20524 18770 20576 18776
rect 20536 18714 20564 18770
rect 20444 18686 20564 18714
rect 20444 18426 20472 18686
rect 20524 18624 20576 18630
rect 20524 18566 20576 18572
rect 20432 18420 20484 18426
rect 20432 18362 20484 18368
rect 20432 17740 20484 17746
rect 20432 17682 20484 17688
rect 20444 16998 20472 17682
rect 20432 16992 20484 16998
rect 20432 16934 20484 16940
rect 20444 16250 20472 16934
rect 20432 16244 20484 16250
rect 20432 16186 20484 16192
rect 20340 15020 20392 15026
rect 20340 14962 20392 14968
rect 20248 14884 20300 14890
rect 20248 14826 20300 14832
rect 20260 14074 20288 14826
rect 20352 14618 20380 14962
rect 20340 14612 20392 14618
rect 20340 14554 20392 14560
rect 20248 14068 20300 14074
rect 20248 14010 20300 14016
rect 20156 13456 20208 13462
rect 20156 13398 20208 13404
rect 20168 12986 20196 13398
rect 20340 13320 20392 13326
rect 20340 13262 20392 13268
rect 20156 12980 20208 12986
rect 20156 12922 20208 12928
rect 19788 12844 19840 12850
rect 19788 12786 19840 12792
rect 20248 12844 20300 12850
rect 20248 12786 20300 12792
rect 19696 12776 19748 12782
rect 19696 12718 19748 12724
rect 18960 12368 19012 12374
rect 18960 12310 19012 12316
rect 19604 12368 19656 12374
rect 19604 12310 19656 12316
rect 19708 12306 19736 12718
rect 19788 12436 19840 12442
rect 19788 12378 19840 12384
rect 19696 12300 19748 12306
rect 19696 12242 19748 12248
rect 18868 12232 18920 12238
rect 18868 12174 18920 12180
rect 18776 12164 18828 12170
rect 18776 12106 18828 12112
rect 18684 11892 18736 11898
rect 18684 11834 18736 11840
rect 18500 11824 18552 11830
rect 18500 11766 18552 11772
rect 18222 11656 18278 11665
rect 18512 11642 18540 11766
rect 18222 11591 18278 11600
rect 18420 11614 18540 11642
rect 18592 11620 18644 11626
rect 18132 11212 18184 11218
rect 18132 11154 18184 11160
rect 18040 11144 18092 11150
rect 18040 11086 18092 11092
rect 18052 10606 18080 11086
rect 18236 11082 18264 11591
rect 18420 11558 18448 11614
rect 18592 11562 18644 11568
rect 18408 11552 18460 11558
rect 18604 11506 18632 11562
rect 18408 11494 18460 11500
rect 18224 11076 18276 11082
rect 18224 11018 18276 11024
rect 18040 10600 18092 10606
rect 18040 10542 18092 10548
rect 18314 10568 18370 10577
rect 18314 10503 18316 10512
rect 18368 10503 18370 10512
rect 18316 10474 18368 10480
rect 18420 9926 18448 11494
rect 18512 11478 18632 11506
rect 18512 11286 18540 11478
rect 18500 11280 18552 11286
rect 18500 11222 18552 11228
rect 18512 11014 18540 11222
rect 18696 11014 18724 11834
rect 18880 11762 18908 12174
rect 19604 12164 19656 12170
rect 19604 12106 19656 12112
rect 19616 11830 19644 12106
rect 19800 11898 19828 12378
rect 20260 12238 20288 12786
rect 20248 12232 20300 12238
rect 20248 12174 20300 12180
rect 20352 12102 20380 13262
rect 20430 12744 20486 12753
rect 20430 12679 20432 12688
rect 20484 12679 20486 12688
rect 20432 12650 20484 12656
rect 20430 12336 20486 12345
rect 20430 12271 20486 12280
rect 20340 12096 20392 12102
rect 20340 12038 20392 12044
rect 19788 11892 19840 11898
rect 19788 11834 19840 11840
rect 19604 11824 19656 11830
rect 19604 11766 19656 11772
rect 18868 11756 18920 11762
rect 18868 11698 18920 11704
rect 18776 11688 18828 11694
rect 18774 11656 18776 11665
rect 18828 11656 18830 11665
rect 18774 11591 18830 11600
rect 19150 11452 19446 11472
rect 19206 11450 19230 11452
rect 19286 11450 19310 11452
rect 19366 11450 19390 11452
rect 19228 11398 19230 11450
rect 19292 11398 19304 11450
rect 19366 11398 19368 11450
rect 19206 11396 19230 11398
rect 19286 11396 19310 11398
rect 19366 11396 19390 11398
rect 19150 11376 19446 11396
rect 20352 11257 20380 12038
rect 20338 11248 20394 11257
rect 18776 11212 18828 11218
rect 20444 11218 20472 12271
rect 20338 11183 20394 11192
rect 20432 11212 20484 11218
rect 18776 11154 18828 11160
rect 20432 11154 20484 11160
rect 18500 11008 18552 11014
rect 18500 10950 18552 10956
rect 18684 11008 18736 11014
rect 18684 10950 18736 10956
rect 18512 10538 18540 10950
rect 18696 10810 18724 10950
rect 18684 10804 18736 10810
rect 18684 10746 18736 10752
rect 18500 10532 18552 10538
rect 18500 10474 18552 10480
rect 18512 10198 18540 10474
rect 18500 10192 18552 10198
rect 18500 10134 18552 10140
rect 18696 10130 18724 10746
rect 18684 10124 18736 10130
rect 18684 10066 18736 10072
rect 17856 9920 17908 9926
rect 17854 9888 17856 9897
rect 18408 9920 18460 9926
rect 17908 9888 17910 9897
rect 18408 9862 18460 9868
rect 18592 9920 18644 9926
rect 18592 9862 18644 9868
rect 17854 9823 17910 9832
rect 18420 9722 18448 9862
rect 18408 9716 18460 9722
rect 18408 9658 18460 9664
rect 17856 9444 17908 9450
rect 17856 9386 17908 9392
rect 17868 8974 17896 9386
rect 18408 9376 18460 9382
rect 18408 9318 18460 9324
rect 17856 8968 17908 8974
rect 17854 8936 17856 8945
rect 17908 8936 17910 8945
rect 17854 8871 17910 8880
rect 18420 8430 18448 9318
rect 18408 8424 18460 8430
rect 18408 8366 18460 8372
rect 16752 8298 16804 8304
rect 17684 8316 17804 8344
rect 16764 8004 16792 8298
rect 16936 8016 16988 8022
rect 16566 7984 16622 7993
rect 16764 7976 16936 8004
rect 16936 7958 16988 7964
rect 16566 7919 16622 7928
rect 16580 7721 16608 7919
rect 16566 7712 16622 7721
rect 16566 7647 16622 7656
rect 16948 7274 16976 7958
rect 17028 7948 17080 7954
rect 17028 7890 17080 7896
rect 17040 7546 17068 7890
rect 17028 7540 17080 7546
rect 17028 7482 17080 7488
rect 16936 7268 16988 7274
rect 16936 7210 16988 7216
rect 16658 7032 16714 7041
rect 16658 6967 16714 6976
rect 16106 6831 16162 6840
rect 16384 6860 16436 6866
rect 16384 6802 16436 6808
rect 16016 6792 16068 6798
rect 16016 6734 16068 6740
rect 15740 6656 15792 6662
rect 15740 6598 15792 6604
rect 15462 5672 15518 5681
rect 15462 5607 15518 5616
rect 15556 5568 15608 5574
rect 15556 5510 15608 5516
rect 15280 5160 15332 5166
rect 15280 5102 15332 5108
rect 15096 4684 15148 4690
rect 15096 4626 15148 4632
rect 14484 4380 14780 4400
rect 14540 4378 14564 4380
rect 14620 4378 14644 4380
rect 14700 4378 14724 4380
rect 14562 4326 14564 4378
rect 14626 4326 14638 4378
rect 14700 4326 14702 4378
rect 14540 4324 14564 4326
rect 14620 4324 14644 4326
rect 14700 4324 14724 4326
rect 14484 4304 14780 4324
rect 14176 4140 14228 4146
rect 14176 4082 14228 4088
rect 14268 4140 14320 4146
rect 14268 4082 14320 4088
rect 14188 3738 14216 4082
rect 14176 3732 14228 3738
rect 14176 3674 14228 3680
rect 13900 3528 13952 3534
rect 13900 3470 13952 3476
rect 13624 3392 13676 3398
rect 13624 3334 13676 3340
rect 13806 3360 13862 3369
rect 13636 3194 13664 3334
rect 13806 3295 13862 3304
rect 13624 3188 13676 3194
rect 13624 3130 13676 3136
rect 13820 3058 13848 3295
rect 14280 3058 14308 4082
rect 14820 3936 14872 3942
rect 14820 3878 14872 3884
rect 14832 3505 14860 3878
rect 15108 3738 15136 4626
rect 15280 4480 15332 4486
rect 15280 4422 15332 4428
rect 15096 3732 15148 3738
rect 15096 3674 15148 3680
rect 14912 3596 14964 3602
rect 14912 3538 14964 3544
rect 14818 3496 14874 3505
rect 14818 3431 14874 3440
rect 14484 3292 14780 3312
rect 14540 3290 14564 3292
rect 14620 3290 14644 3292
rect 14700 3290 14724 3292
rect 14562 3238 14564 3290
rect 14626 3238 14638 3290
rect 14700 3238 14702 3290
rect 14540 3236 14564 3238
rect 14620 3236 14644 3238
rect 14700 3236 14724 3238
rect 14484 3216 14780 3236
rect 13808 3052 13860 3058
rect 13808 2994 13860 3000
rect 14268 3052 14320 3058
rect 14268 2994 14320 3000
rect 14358 2952 14414 2961
rect 14924 2922 14952 3538
rect 15292 3233 15320 4422
rect 15568 4146 15596 5510
rect 15556 4140 15608 4146
rect 15556 4082 15608 4088
rect 15568 3670 15596 4082
rect 15752 3913 15780 6598
rect 16028 6322 16056 6734
rect 16290 6352 16346 6361
rect 16016 6316 16068 6322
rect 16290 6287 16292 6296
rect 16016 6258 16068 6264
rect 16344 6287 16346 6296
rect 16292 6258 16344 6264
rect 16028 5914 16056 6258
rect 16016 5908 16068 5914
rect 16016 5850 16068 5856
rect 16198 5672 16254 5681
rect 16304 5642 16332 6258
rect 16396 6186 16424 6802
rect 16384 6180 16436 6186
rect 16384 6122 16436 6128
rect 16672 5710 16700 6967
rect 16752 6792 16804 6798
rect 16752 6734 16804 6740
rect 16764 5846 16792 6734
rect 16752 5840 16804 5846
rect 16752 5782 16804 5788
rect 16660 5704 16712 5710
rect 16660 5646 16712 5652
rect 16198 5607 16254 5616
rect 16292 5636 16344 5642
rect 16108 5024 16160 5030
rect 16108 4966 16160 4972
rect 16120 4185 16148 4966
rect 16212 4690 16240 5607
rect 16292 5578 16344 5584
rect 16672 5234 16700 5646
rect 16764 5370 16792 5782
rect 16752 5364 16804 5370
rect 16752 5306 16804 5312
rect 16660 5228 16712 5234
rect 16660 5170 16712 5176
rect 16948 5098 16976 7210
rect 17684 6322 17712 8316
rect 17762 8256 17818 8265
rect 17762 8191 17818 8200
rect 17776 8090 17804 8191
rect 18420 8090 18448 8366
rect 17764 8084 17816 8090
rect 17764 8026 17816 8032
rect 18408 8084 18460 8090
rect 18408 8026 18460 8032
rect 17776 6934 17804 8026
rect 18132 7744 18184 7750
rect 18132 7686 18184 7692
rect 17854 7440 17910 7449
rect 17854 7375 17856 7384
rect 17908 7375 17910 7384
rect 17856 7346 17908 7352
rect 17868 7206 17896 7346
rect 18144 7313 18172 7686
rect 18408 7404 18460 7410
rect 18408 7346 18460 7352
rect 18130 7304 18186 7313
rect 18130 7239 18132 7248
rect 18184 7239 18186 7248
rect 18132 7210 18184 7216
rect 17856 7200 17908 7206
rect 18420 7177 18448 7346
rect 17856 7142 17908 7148
rect 18406 7168 18462 7177
rect 18406 7103 18462 7112
rect 17764 6928 17816 6934
rect 17764 6870 17816 6876
rect 17776 6458 17804 6870
rect 18420 6798 18448 7103
rect 18040 6792 18092 6798
rect 18040 6734 18092 6740
rect 18408 6792 18460 6798
rect 18408 6734 18460 6740
rect 17764 6452 17816 6458
rect 17764 6394 17816 6400
rect 17672 6316 17724 6322
rect 17672 6258 17724 6264
rect 17684 5914 17712 6258
rect 18052 5914 18080 6734
rect 18132 6316 18184 6322
rect 18132 6258 18184 6264
rect 17672 5908 17724 5914
rect 17672 5850 17724 5856
rect 18040 5908 18092 5914
rect 18040 5850 18092 5856
rect 17856 5772 17908 5778
rect 17856 5714 17908 5720
rect 17026 5400 17082 5409
rect 17868 5370 17896 5714
rect 17026 5335 17082 5344
rect 17856 5364 17908 5370
rect 17040 5302 17068 5335
rect 17856 5306 17908 5312
rect 17028 5296 17080 5302
rect 17028 5238 17080 5244
rect 16936 5092 16988 5098
rect 16936 5034 16988 5040
rect 16842 4992 16898 5001
rect 16842 4927 16898 4936
rect 16856 4729 16884 4927
rect 16948 4758 16976 5034
rect 16936 4752 16988 4758
rect 16842 4720 16898 4729
rect 16200 4684 16252 4690
rect 16936 4694 16988 4700
rect 16842 4655 16898 4664
rect 16200 4626 16252 4632
rect 16212 4298 16240 4626
rect 16212 4270 16332 4298
rect 16948 4282 16976 4694
rect 17120 4480 17172 4486
rect 17120 4422 17172 4428
rect 17488 4480 17540 4486
rect 17488 4422 17540 4428
rect 16106 4176 16162 4185
rect 16106 4111 16162 4120
rect 16200 4140 16252 4146
rect 16200 4082 16252 4088
rect 15738 3904 15794 3913
rect 15738 3839 15794 3848
rect 15556 3664 15608 3670
rect 16212 3641 16240 4082
rect 16304 3738 16332 4270
rect 16936 4276 16988 4282
rect 16936 4218 16988 4224
rect 16292 3732 16344 3738
rect 16292 3674 16344 3680
rect 17132 3670 17160 4422
rect 17500 4010 17528 4422
rect 17578 4040 17634 4049
rect 17488 4004 17540 4010
rect 17578 3975 17634 3984
rect 17488 3946 17540 3952
rect 17120 3664 17172 3670
rect 15556 3606 15608 3612
rect 16198 3632 16254 3641
rect 15278 3224 15334 3233
rect 15568 3194 15596 3606
rect 17120 3606 17172 3612
rect 16198 3567 16254 3576
rect 16212 3534 16240 3567
rect 16200 3528 16252 3534
rect 16200 3470 16252 3476
rect 16292 3460 16344 3466
rect 16292 3402 16344 3408
rect 16016 3392 16068 3398
rect 16016 3334 16068 3340
rect 15278 3159 15334 3168
rect 15556 3188 15608 3194
rect 15556 3130 15608 3136
rect 16028 3097 16056 3334
rect 16014 3088 16070 3097
rect 16014 3023 16070 3032
rect 14358 2887 14414 2896
rect 14912 2916 14964 2922
rect 13532 2644 13584 2650
rect 13532 2586 13584 2592
rect 13808 2508 13860 2514
rect 13808 2450 13860 2456
rect 13820 1873 13848 2450
rect 13992 2304 14044 2310
rect 13992 2246 14044 2252
rect 14004 1873 14032 2246
rect 14372 1986 14400 2887
rect 14912 2858 14964 2864
rect 14818 2816 14874 2825
rect 14818 2751 14874 2760
rect 14832 2650 14860 2751
rect 16304 2650 16332 3402
rect 17132 3194 17160 3606
rect 17120 3188 17172 3194
rect 17120 3130 17172 3136
rect 16568 2916 16620 2922
rect 16568 2858 16620 2864
rect 14820 2644 14872 2650
rect 14820 2586 14872 2592
rect 16292 2644 16344 2650
rect 16292 2586 16344 2592
rect 14484 2204 14780 2224
rect 14540 2202 14564 2204
rect 14620 2202 14644 2204
rect 14700 2202 14724 2204
rect 14562 2150 14564 2202
rect 14626 2150 14638 2202
rect 14700 2150 14702 2202
rect 14540 2148 14564 2150
rect 14620 2148 14644 2150
rect 14700 2148 14724 2150
rect 14484 2128 14780 2148
rect 15462 2000 15518 2009
rect 14372 1958 14492 1986
rect 13806 1864 13862 1873
rect 13806 1799 13862 1808
rect 13990 1864 14046 1873
rect 13990 1799 14046 1808
rect 14464 480 14492 1958
rect 15462 1935 15518 1944
rect 15476 480 15504 1935
rect 16580 480 16608 2858
rect 17500 2553 17528 3946
rect 17592 3534 17620 3975
rect 17580 3528 17632 3534
rect 17580 3470 17632 3476
rect 18052 3466 18080 5850
rect 18144 3534 18172 6258
rect 18604 5778 18632 9862
rect 18696 9178 18724 10066
rect 18788 9738 18816 11154
rect 18960 11144 19012 11150
rect 20444 11121 20472 11154
rect 18960 11086 19012 11092
rect 20430 11112 20486 11121
rect 18972 10674 19000 11086
rect 19144 11076 19196 11082
rect 19064 11036 19144 11064
rect 18960 10668 19012 10674
rect 18960 10610 19012 10616
rect 18972 10266 19000 10610
rect 18960 10260 19012 10266
rect 18960 10202 19012 10208
rect 18972 10062 19000 10202
rect 18960 10056 19012 10062
rect 18960 9998 19012 10004
rect 18788 9710 18908 9738
rect 18972 9722 19000 9998
rect 18880 9450 18908 9710
rect 18960 9716 19012 9722
rect 18960 9658 19012 9664
rect 18960 9512 19012 9518
rect 18960 9454 19012 9460
rect 18868 9444 18920 9450
rect 18868 9386 18920 9392
rect 18684 9172 18736 9178
rect 18684 9114 18736 9120
rect 18880 9110 18908 9386
rect 18972 9178 19000 9454
rect 18960 9172 19012 9178
rect 18960 9114 19012 9120
rect 18868 9104 18920 9110
rect 18868 9046 18920 9052
rect 19064 8809 19092 11036
rect 20430 11047 20486 11056
rect 19144 11018 19196 11024
rect 19420 11008 19472 11014
rect 19420 10950 19472 10956
rect 19432 10742 19460 10950
rect 19512 10804 19564 10810
rect 19512 10746 19564 10752
rect 19420 10736 19472 10742
rect 19420 10678 19472 10684
rect 19150 10364 19446 10384
rect 19206 10362 19230 10364
rect 19286 10362 19310 10364
rect 19366 10362 19390 10364
rect 19228 10310 19230 10362
rect 19292 10310 19304 10362
rect 19366 10310 19368 10362
rect 19206 10308 19230 10310
rect 19286 10308 19310 10310
rect 19366 10308 19390 10310
rect 19150 10288 19446 10308
rect 19524 10266 19552 10746
rect 19696 10736 19748 10742
rect 19696 10678 19748 10684
rect 19602 10432 19658 10441
rect 19602 10367 19658 10376
rect 19512 10260 19564 10266
rect 19512 10202 19564 10208
rect 19524 9722 19552 10202
rect 19512 9716 19564 9722
rect 19512 9658 19564 9664
rect 19150 9276 19446 9296
rect 19206 9274 19230 9276
rect 19286 9274 19310 9276
rect 19366 9274 19390 9276
rect 19228 9222 19230 9274
rect 19292 9222 19304 9274
rect 19366 9222 19368 9274
rect 19206 9220 19230 9222
rect 19286 9220 19310 9222
rect 19366 9220 19390 9222
rect 19150 9200 19446 9220
rect 19616 9178 19644 10367
rect 19708 10266 19736 10678
rect 19880 10532 19932 10538
rect 19880 10474 19932 10480
rect 19696 10260 19748 10266
rect 19696 10202 19748 10208
rect 19788 9376 19840 9382
rect 19788 9318 19840 9324
rect 19604 9172 19656 9178
rect 19604 9114 19656 9120
rect 19696 9036 19748 9042
rect 19696 8978 19748 8984
rect 19050 8800 19106 8809
rect 19050 8735 19106 8744
rect 18960 8424 19012 8430
rect 18960 8366 19012 8372
rect 18972 7954 19000 8366
rect 19064 7954 19092 8735
rect 19150 8188 19446 8208
rect 19206 8186 19230 8188
rect 19286 8186 19310 8188
rect 19366 8186 19390 8188
rect 19228 8134 19230 8186
rect 19292 8134 19304 8186
rect 19366 8134 19368 8186
rect 19206 8132 19230 8134
rect 19286 8132 19310 8134
rect 19366 8132 19390 8134
rect 19150 8112 19446 8132
rect 19708 8090 19736 8978
rect 19800 8430 19828 9318
rect 19788 8424 19840 8430
rect 19788 8366 19840 8372
rect 19696 8084 19748 8090
rect 19696 8026 19748 8032
rect 18960 7948 19012 7954
rect 18960 7890 19012 7896
rect 19052 7948 19104 7954
rect 19052 7890 19104 7896
rect 18972 7546 19000 7890
rect 18960 7540 19012 7546
rect 18960 7482 19012 7488
rect 19064 7002 19092 7890
rect 19604 7336 19656 7342
rect 19604 7278 19656 7284
rect 19150 7100 19446 7120
rect 19206 7098 19230 7100
rect 19286 7098 19310 7100
rect 19366 7098 19390 7100
rect 19228 7046 19230 7098
rect 19292 7046 19304 7098
rect 19366 7046 19368 7098
rect 19206 7044 19230 7046
rect 19286 7044 19310 7046
rect 19366 7044 19390 7046
rect 19150 7024 19446 7044
rect 19052 6996 19104 7002
rect 19052 6938 19104 6944
rect 19616 6458 19644 7278
rect 19604 6452 19656 6458
rect 19604 6394 19656 6400
rect 19616 6254 19644 6394
rect 19604 6248 19656 6254
rect 19604 6190 19656 6196
rect 18958 6080 19014 6089
rect 18958 6015 19014 6024
rect 18776 5908 18828 5914
rect 18776 5850 18828 5856
rect 18592 5772 18644 5778
rect 18592 5714 18644 5720
rect 18604 5370 18632 5714
rect 18684 5704 18736 5710
rect 18684 5646 18736 5652
rect 18592 5364 18644 5370
rect 18592 5306 18644 5312
rect 18604 4826 18632 5306
rect 18592 4820 18644 4826
rect 18592 4762 18644 4768
rect 18696 4690 18724 5646
rect 18788 5234 18816 5850
rect 18972 5681 19000 6015
rect 19150 6012 19446 6032
rect 19206 6010 19230 6012
rect 19286 6010 19310 6012
rect 19366 6010 19390 6012
rect 19228 5958 19230 6010
rect 19292 5958 19304 6010
rect 19366 5958 19368 6010
rect 19206 5956 19230 5958
rect 19286 5956 19310 5958
rect 19366 5956 19390 5958
rect 19150 5936 19446 5956
rect 19616 5846 19644 6190
rect 19604 5840 19656 5846
rect 19604 5782 19656 5788
rect 18958 5672 19014 5681
rect 18958 5607 19014 5616
rect 18776 5228 18828 5234
rect 18776 5170 18828 5176
rect 18776 5092 18828 5098
rect 18776 5034 18828 5040
rect 18788 4758 18816 5034
rect 19150 4924 19446 4944
rect 19206 4922 19230 4924
rect 19286 4922 19310 4924
rect 19366 4922 19390 4924
rect 19228 4870 19230 4922
rect 19292 4870 19304 4922
rect 19366 4870 19368 4922
rect 19206 4868 19230 4870
rect 19286 4868 19310 4870
rect 19366 4868 19390 4870
rect 19150 4848 19446 4868
rect 18776 4752 18828 4758
rect 18776 4694 18828 4700
rect 18684 4684 18736 4690
rect 18684 4626 18736 4632
rect 18696 4214 18724 4626
rect 18788 4282 18816 4694
rect 19512 4480 19564 4486
rect 19512 4422 19564 4428
rect 18776 4276 18828 4282
rect 18776 4218 18828 4224
rect 18684 4208 18736 4214
rect 18684 4150 18736 4156
rect 19052 4004 19104 4010
rect 19052 3946 19104 3952
rect 18960 3596 19012 3602
rect 18960 3538 19012 3544
rect 18132 3528 18184 3534
rect 18132 3470 18184 3476
rect 18040 3460 18092 3466
rect 18040 3402 18092 3408
rect 17672 3392 17724 3398
rect 17672 3334 17724 3340
rect 17684 3097 17712 3334
rect 17670 3088 17726 3097
rect 18052 3058 18080 3402
rect 18592 3392 18644 3398
rect 18592 3334 18644 3340
rect 17670 3023 17672 3032
rect 17724 3023 17726 3032
rect 18040 3052 18092 3058
rect 17672 2994 17724 3000
rect 18040 2994 18092 3000
rect 18500 2916 18552 2922
rect 18500 2858 18552 2864
rect 17486 2544 17542 2553
rect 16660 2508 16712 2514
rect 17486 2479 17542 2488
rect 16660 2450 16712 2456
rect 16672 1737 16700 2450
rect 17488 2372 17540 2378
rect 17488 2314 17540 2320
rect 16658 1728 16714 1737
rect 16658 1663 16714 1672
rect 17500 1170 17528 2314
rect 17580 2304 17632 2310
rect 17580 2246 17632 2252
rect 17592 1465 17620 2246
rect 18512 1601 18540 2858
rect 18498 1592 18554 1601
rect 18498 1527 18554 1536
rect 17578 1456 17634 1465
rect 17578 1391 17634 1400
rect 17500 1142 17620 1170
rect 17592 480 17620 1142
rect 18604 480 18632 3334
rect 18682 2952 18738 2961
rect 18682 2887 18738 2896
rect 18696 2582 18724 2887
rect 18684 2576 18736 2582
rect 18684 2518 18736 2524
rect 18972 2310 19000 3538
rect 19064 3466 19092 3946
rect 19524 3942 19552 4422
rect 19708 4146 19736 8026
rect 19800 7342 19828 8366
rect 19788 7336 19840 7342
rect 19788 7278 19840 7284
rect 19800 7002 19828 7278
rect 19788 6996 19840 7002
rect 19788 6938 19840 6944
rect 19892 6254 19920 10474
rect 20444 10266 20472 11047
rect 20156 10260 20208 10266
rect 20156 10202 20208 10208
rect 20432 10260 20484 10266
rect 20432 10202 20484 10208
rect 20168 8634 20196 10202
rect 20430 8664 20486 8673
rect 19972 8628 20024 8634
rect 19972 8570 20024 8576
rect 20156 8628 20208 8634
rect 20430 8599 20486 8608
rect 20156 8570 20208 8576
rect 19880 6248 19932 6254
rect 19880 6190 19932 6196
rect 19892 5846 19920 6190
rect 19880 5840 19932 5846
rect 19880 5782 19932 5788
rect 19984 5778 20012 8570
rect 20248 8424 20300 8430
rect 20248 8366 20300 8372
rect 20064 8356 20116 8362
rect 20064 8298 20116 8304
rect 19972 5772 20024 5778
rect 19972 5714 20024 5720
rect 19984 5302 20012 5714
rect 19972 5296 20024 5302
rect 19972 5238 20024 5244
rect 19972 5160 20024 5166
rect 19972 5102 20024 5108
rect 19696 4140 19748 4146
rect 19696 4082 19748 4088
rect 19512 3936 19564 3942
rect 19512 3878 19564 3884
rect 19150 3836 19446 3856
rect 19206 3834 19230 3836
rect 19286 3834 19310 3836
rect 19366 3834 19390 3836
rect 19228 3782 19230 3834
rect 19292 3782 19304 3834
rect 19366 3782 19368 3834
rect 19206 3780 19230 3782
rect 19286 3780 19310 3782
rect 19366 3780 19390 3782
rect 19150 3760 19446 3780
rect 19052 3460 19104 3466
rect 19052 3402 19104 3408
rect 19064 2378 19092 3402
rect 19708 3058 19736 4082
rect 19984 3738 20012 5102
rect 20076 4706 20104 8298
rect 20156 7540 20208 7546
rect 20260 7528 20288 8366
rect 20208 7500 20288 7528
rect 20156 7482 20208 7488
rect 20156 7404 20208 7410
rect 20156 7346 20208 7352
rect 20168 5250 20196 7346
rect 20444 6866 20472 8599
rect 20432 6860 20484 6866
rect 20432 6802 20484 6808
rect 20340 5840 20392 5846
rect 20444 5828 20472 6802
rect 20392 5800 20472 5828
rect 20340 5782 20392 5788
rect 20248 5704 20300 5710
rect 20248 5646 20300 5652
rect 20260 5370 20288 5646
rect 20248 5364 20300 5370
rect 20248 5306 20300 5312
rect 20168 5234 20288 5250
rect 20168 5228 20300 5234
rect 20168 5222 20248 5228
rect 20248 5170 20300 5176
rect 20076 4690 20288 4706
rect 20076 4684 20300 4690
rect 20076 4678 20248 4684
rect 20248 4626 20300 4632
rect 20260 4282 20288 4626
rect 20248 4276 20300 4282
rect 20248 4218 20300 4224
rect 20156 3936 20208 3942
rect 20208 3884 20380 3890
rect 20156 3878 20380 3884
rect 20168 3862 20380 3878
rect 19972 3732 20024 3738
rect 19972 3674 20024 3680
rect 19696 3052 19748 3058
rect 19696 2994 19748 3000
rect 19696 2916 19748 2922
rect 19696 2858 19748 2864
rect 20064 2916 20116 2922
rect 20064 2858 20116 2864
rect 19150 2748 19446 2768
rect 19206 2746 19230 2748
rect 19286 2746 19310 2748
rect 19366 2746 19390 2748
rect 19228 2694 19230 2746
rect 19292 2694 19304 2746
rect 19366 2694 19368 2746
rect 19206 2692 19230 2694
rect 19286 2692 19310 2694
rect 19366 2692 19390 2694
rect 19150 2672 19446 2692
rect 19708 2582 19736 2858
rect 19696 2576 19748 2582
rect 19696 2518 19748 2524
rect 19052 2372 19104 2378
rect 19052 2314 19104 2320
rect 20076 2310 20104 2858
rect 20352 2514 20380 3862
rect 20432 3732 20484 3738
rect 20432 3674 20484 3680
rect 20444 3194 20472 3674
rect 20536 3670 20564 18566
rect 20708 17536 20760 17542
rect 20708 17478 20760 17484
rect 20720 16726 20748 17478
rect 20708 16720 20760 16726
rect 20708 16662 20760 16668
rect 20720 16250 20748 16662
rect 20708 16244 20760 16250
rect 20708 16186 20760 16192
rect 20616 14544 20668 14550
rect 20616 14486 20668 14492
rect 20628 14074 20656 14486
rect 20616 14068 20668 14074
rect 20616 14010 20668 14016
rect 20628 12374 20656 14010
rect 20708 12912 20760 12918
rect 20708 12854 20760 12860
rect 20616 12368 20668 12374
rect 20616 12310 20668 12316
rect 20628 11762 20656 12310
rect 20720 12170 20748 12854
rect 20708 12164 20760 12170
rect 20708 12106 20760 12112
rect 20812 11898 20840 20703
rect 20904 15978 20932 23559
rect 21534 23488 21590 23497
rect 21534 23423 21590 23432
rect 20982 19408 21038 19417
rect 20982 19343 21038 19352
rect 20892 15972 20944 15978
rect 20892 15914 20944 15920
rect 20904 15638 20932 15914
rect 20892 15632 20944 15638
rect 20892 15574 20944 15580
rect 20904 15162 20932 15574
rect 20892 15156 20944 15162
rect 20892 15098 20944 15104
rect 20904 14550 20932 15098
rect 20892 14544 20944 14550
rect 20892 14486 20944 14492
rect 20892 14408 20944 14414
rect 20892 14350 20944 14356
rect 20904 14074 20932 14350
rect 20892 14068 20944 14074
rect 20892 14010 20944 14016
rect 20892 12776 20944 12782
rect 20892 12718 20944 12724
rect 20996 12730 21024 19343
rect 21548 17882 21576 23423
rect 22284 18170 22312 27520
rect 22914 27432 22970 27441
rect 22914 27367 22970 27376
rect 22928 23798 22956 27367
rect 24294 26344 24350 26353
rect 24294 26279 24350 26288
rect 23817 25052 24113 25072
rect 23873 25050 23897 25052
rect 23953 25050 23977 25052
rect 24033 25050 24057 25052
rect 23895 24998 23897 25050
rect 23959 24998 23971 25050
rect 24033 24998 24035 25050
rect 23873 24996 23897 24998
rect 23953 24996 23977 24998
rect 24033 24996 24057 24998
rect 23817 24976 24113 24996
rect 23190 24304 23246 24313
rect 23190 24239 23246 24248
rect 22916 23792 22968 23798
rect 22916 23734 22968 23740
rect 23008 23520 23060 23526
rect 23006 23488 23008 23497
rect 23060 23488 23062 23497
rect 23006 23423 23062 23432
rect 22364 21344 22416 21350
rect 22364 21286 22416 21292
rect 22008 18142 22312 18170
rect 21536 17876 21588 17882
rect 21536 17818 21588 17824
rect 21548 17270 21576 17818
rect 21536 17264 21588 17270
rect 21536 17206 21588 17212
rect 21628 17196 21680 17202
rect 21628 17138 21680 17144
rect 21640 16590 21668 17138
rect 21444 16584 21496 16590
rect 21444 16526 21496 16532
rect 21628 16584 21680 16590
rect 21628 16526 21680 16532
rect 21456 16114 21484 16526
rect 21720 16244 21772 16250
rect 21720 16186 21772 16192
rect 21444 16108 21496 16114
rect 21444 16050 21496 16056
rect 21456 15706 21484 16050
rect 21732 15978 21760 16186
rect 21720 15972 21772 15978
rect 21720 15914 21772 15920
rect 21444 15700 21496 15706
rect 21444 15642 21496 15648
rect 21732 15570 21760 15914
rect 21720 15564 21772 15570
rect 21720 15506 21772 15512
rect 21628 14884 21680 14890
rect 21628 14826 21680 14832
rect 21444 14612 21496 14618
rect 21444 14554 21496 14560
rect 21456 14074 21484 14554
rect 21640 14550 21668 14826
rect 21628 14544 21680 14550
rect 21628 14486 21680 14492
rect 21444 14068 21496 14074
rect 21444 14010 21496 14016
rect 21168 13932 21220 13938
rect 21168 13874 21220 13880
rect 21180 13462 21208 13874
rect 21456 13870 21484 14010
rect 21640 13938 21668 14486
rect 21628 13932 21680 13938
rect 21628 13874 21680 13880
rect 21444 13864 21496 13870
rect 21444 13806 21496 13812
rect 22008 13569 22036 18142
rect 22088 18080 22140 18086
rect 22088 18022 22140 18028
rect 21994 13560 22050 13569
rect 21994 13495 22050 13504
rect 21168 13456 21220 13462
rect 21168 13398 21220 13404
rect 21076 13184 21128 13190
rect 21076 13126 21128 13132
rect 21088 12850 21116 13126
rect 21076 12844 21128 12850
rect 21076 12786 21128 12792
rect 21444 12776 21496 12782
rect 21442 12744 21444 12753
rect 21496 12744 21498 12753
rect 20904 12442 20932 12718
rect 20996 12702 21208 12730
rect 20892 12436 20944 12442
rect 20892 12378 20944 12384
rect 20800 11892 20852 11898
rect 20800 11834 20852 11840
rect 20616 11756 20668 11762
rect 20616 11698 20668 11704
rect 20892 11620 20944 11626
rect 20892 11562 20944 11568
rect 20708 11552 20760 11558
rect 20708 11494 20760 11500
rect 20720 11286 20748 11494
rect 20708 11280 20760 11286
rect 20708 11222 20760 11228
rect 20904 11218 20932 11562
rect 20892 11212 20944 11218
rect 20892 11154 20944 11160
rect 20614 10704 20670 10713
rect 20614 10639 20616 10648
rect 20668 10639 20670 10648
rect 20616 10610 20668 10616
rect 20628 8634 20656 10610
rect 20904 10606 20932 11154
rect 20984 11144 21036 11150
rect 20984 11086 21036 11092
rect 20892 10600 20944 10606
rect 20892 10542 20944 10548
rect 20996 10130 21024 11086
rect 20984 10124 21036 10130
rect 20984 10066 21036 10072
rect 21180 10010 21208 12702
rect 21442 12679 21498 12688
rect 21904 12300 21956 12306
rect 21904 12242 21956 12248
rect 21536 11756 21588 11762
rect 21536 11698 21588 11704
rect 21352 11688 21404 11694
rect 21352 11630 21404 11636
rect 21364 11354 21392 11630
rect 21352 11348 21404 11354
rect 21352 11290 21404 11296
rect 21548 10742 21576 11698
rect 21916 11286 21944 12242
rect 21904 11280 21956 11286
rect 21904 11222 21956 11228
rect 21904 10804 21956 10810
rect 21904 10746 21956 10752
rect 21536 10736 21588 10742
rect 21536 10678 21588 10684
rect 21260 10668 21312 10674
rect 21260 10610 21312 10616
rect 20996 9982 21208 10010
rect 20800 9648 20852 9654
rect 20800 9590 20852 9596
rect 20616 8628 20668 8634
rect 20616 8570 20668 8576
rect 20812 8022 20840 9590
rect 20996 9178 21024 9982
rect 21272 9586 21300 10610
rect 21548 10198 21576 10678
rect 21916 10266 21944 10746
rect 21904 10260 21956 10266
rect 21904 10202 21956 10208
rect 21536 10192 21588 10198
rect 21536 10134 21588 10140
rect 21548 9654 21576 10134
rect 21628 10124 21680 10130
rect 21628 10066 21680 10072
rect 21640 9722 21668 10066
rect 22100 10062 22128 18022
rect 22180 17536 22232 17542
rect 22180 17478 22232 17484
rect 22088 10056 22140 10062
rect 22088 9998 22140 10004
rect 22192 9722 22220 17478
rect 22270 15736 22326 15745
rect 22270 15671 22326 15680
rect 22284 15638 22312 15671
rect 22272 15632 22324 15638
rect 22272 15574 22324 15580
rect 22284 15026 22312 15574
rect 22272 15020 22324 15026
rect 22272 14962 22324 14968
rect 22272 14408 22324 14414
rect 22272 14350 22324 14356
rect 22284 13530 22312 14350
rect 22272 13524 22324 13530
rect 22272 13466 22324 13472
rect 22284 13433 22312 13466
rect 22270 13424 22326 13433
rect 22270 13359 22326 13368
rect 21628 9716 21680 9722
rect 21628 9658 21680 9664
rect 21812 9716 21864 9722
rect 21812 9658 21864 9664
rect 22180 9716 22232 9722
rect 22180 9658 22232 9664
rect 21536 9648 21588 9654
rect 21536 9590 21588 9596
rect 21824 9602 21852 9658
rect 21260 9580 21312 9586
rect 21260 9522 21312 9528
rect 21548 9450 21576 9590
rect 21824 9574 21944 9602
rect 21536 9444 21588 9450
rect 21536 9386 21588 9392
rect 20984 9172 21036 9178
rect 20984 9114 21036 9120
rect 21352 9172 21404 9178
rect 21352 9114 21404 9120
rect 20892 8832 20944 8838
rect 20890 8800 20892 8809
rect 20944 8800 20946 8809
rect 20946 8758 21024 8786
rect 20890 8735 20946 8744
rect 20996 8430 21024 8758
rect 20984 8424 21036 8430
rect 20984 8366 21036 8372
rect 21168 8288 21220 8294
rect 21168 8230 21220 8236
rect 20800 8016 20852 8022
rect 20800 7958 20852 7964
rect 20812 7546 20840 7958
rect 20892 7880 20944 7886
rect 20892 7822 20944 7828
rect 20800 7540 20852 7546
rect 20800 7482 20852 7488
rect 20614 7304 20670 7313
rect 20614 7239 20670 7248
rect 20628 6866 20656 7239
rect 20904 7002 20932 7822
rect 21180 7410 21208 8230
rect 21364 7834 21392 9114
rect 21444 9104 21496 9110
rect 21444 9046 21496 9052
rect 21456 8634 21484 9046
rect 21536 8968 21588 8974
rect 21536 8910 21588 8916
rect 21444 8628 21496 8634
rect 21444 8570 21496 8576
rect 21548 8242 21576 8910
rect 21916 8634 21944 9574
rect 21904 8628 21956 8634
rect 21904 8570 21956 8576
rect 21548 8214 21668 8242
rect 21640 8090 21668 8214
rect 21628 8084 21680 8090
rect 21628 8026 21680 8032
rect 21640 7993 21668 8026
rect 21626 7984 21682 7993
rect 21626 7919 21682 7928
rect 22376 7886 22404 21286
rect 23204 20777 23232 24239
rect 23817 23964 24113 23984
rect 23873 23962 23897 23964
rect 23953 23962 23977 23964
rect 24033 23962 24057 23964
rect 23895 23910 23897 23962
rect 23959 23910 23971 23962
rect 24033 23910 24035 23962
rect 23873 23908 23897 23910
rect 23953 23908 23977 23910
rect 24033 23908 24057 23910
rect 23817 23888 24113 23908
rect 24308 23866 24336 26279
rect 24938 25392 24994 25401
rect 24938 25327 24994 25336
rect 24296 23860 24348 23866
rect 24296 23802 24348 23808
rect 24308 23662 24336 23802
rect 24296 23656 24348 23662
rect 24296 23598 24348 23604
rect 24294 23216 24350 23225
rect 24294 23151 24350 23160
rect 23817 22876 24113 22896
rect 23873 22874 23897 22876
rect 23953 22874 23977 22876
rect 24033 22874 24057 22876
rect 23895 22822 23897 22874
rect 23959 22822 23971 22874
rect 24033 22822 24035 22874
rect 23873 22820 23897 22822
rect 23953 22820 23977 22822
rect 24033 22820 24057 22822
rect 23817 22800 24113 22820
rect 24202 22264 24258 22273
rect 24202 22199 24258 22208
rect 23817 21788 24113 21808
rect 23873 21786 23897 21788
rect 23953 21786 23977 21788
rect 24033 21786 24057 21788
rect 23895 21734 23897 21786
rect 23959 21734 23971 21786
rect 24033 21734 24035 21786
rect 23873 21732 23897 21734
rect 23953 21732 23977 21734
rect 24033 21732 24057 21734
rect 23817 21712 24113 21732
rect 24216 21010 24244 22199
rect 24308 21690 24336 23151
rect 24296 21684 24348 21690
rect 24296 21626 24348 21632
rect 24308 21486 24336 21626
rect 24296 21480 24348 21486
rect 24296 21422 24348 21428
rect 24204 21004 24256 21010
rect 24204 20946 24256 20952
rect 23284 20800 23336 20806
rect 23190 20768 23246 20777
rect 23284 20742 23336 20748
rect 23190 20703 23246 20712
rect 23008 19712 23060 19718
rect 23008 19654 23060 19660
rect 23020 19417 23048 19654
rect 23006 19408 23062 19417
rect 23006 19343 23062 19352
rect 23006 19272 23062 19281
rect 23006 19207 23008 19216
rect 23060 19207 23062 19216
rect 23008 19178 23060 19184
rect 23006 18728 23062 18737
rect 23006 18663 23008 18672
rect 23060 18663 23062 18672
rect 23008 18634 23060 18640
rect 23100 18624 23152 18630
rect 23100 18566 23152 18572
rect 23112 18329 23140 18566
rect 23098 18320 23154 18329
rect 23098 18255 23154 18264
rect 22640 18080 22692 18086
rect 22638 18048 22640 18057
rect 22692 18048 22694 18057
rect 22638 17983 22694 17992
rect 22732 17740 22784 17746
rect 22732 17682 22784 17688
rect 22744 16998 22772 17682
rect 23008 17536 23060 17542
rect 23008 17478 23060 17484
rect 22732 16992 22784 16998
rect 22732 16934 22784 16940
rect 22548 16652 22600 16658
rect 22548 16594 22600 16600
rect 22456 16448 22508 16454
rect 22456 16390 22508 16396
rect 22468 15638 22496 16390
rect 22560 16250 22588 16594
rect 22548 16244 22600 16250
rect 22548 16186 22600 16192
rect 22548 15972 22600 15978
rect 22548 15914 22600 15920
rect 22456 15632 22508 15638
rect 22456 15574 22508 15580
rect 22468 15162 22496 15574
rect 22560 15502 22588 15914
rect 22548 15496 22600 15502
rect 22548 15438 22600 15444
rect 22456 15156 22508 15162
rect 22456 15098 22508 15104
rect 22640 14544 22692 14550
rect 22640 14486 22692 14492
rect 22652 14074 22680 14486
rect 22640 14068 22692 14074
rect 22640 14010 22692 14016
rect 22456 13456 22508 13462
rect 22456 13398 22508 13404
rect 22468 12986 22496 13398
rect 22548 13320 22600 13326
rect 22548 13262 22600 13268
rect 22456 12980 22508 12986
rect 22456 12922 22508 12928
rect 22560 12102 22588 13262
rect 22640 12776 22692 12782
rect 22640 12718 22692 12724
rect 22652 12345 22680 12718
rect 22638 12336 22694 12345
rect 22638 12271 22694 12280
rect 22548 12096 22600 12102
rect 22548 12038 22600 12044
rect 22560 11506 22588 12038
rect 22468 11478 22588 11506
rect 22468 10033 22496 11478
rect 22744 11286 22772 16934
rect 23020 15337 23048 17478
rect 23296 16130 23324 20742
rect 23817 20700 24113 20720
rect 23873 20698 23897 20700
rect 23953 20698 23977 20700
rect 24033 20698 24057 20700
rect 23895 20646 23897 20698
rect 23959 20646 23971 20698
rect 24033 20646 24035 20698
rect 23873 20644 23897 20646
rect 23953 20644 23977 20646
rect 24033 20644 24057 20646
rect 23817 20624 24113 20644
rect 24216 20602 24244 20946
rect 24204 20596 24256 20602
rect 24204 20538 24256 20544
rect 23817 19612 24113 19632
rect 23873 19610 23897 19612
rect 23953 19610 23977 19612
rect 24033 19610 24057 19612
rect 23895 19558 23897 19610
rect 23959 19558 23971 19610
rect 24033 19558 24035 19610
rect 23873 19556 23897 19558
rect 23953 19556 23977 19558
rect 24033 19556 24057 19558
rect 23817 19536 24113 19556
rect 24202 19136 24258 19145
rect 24202 19071 24258 19080
rect 23468 18828 23520 18834
rect 23468 18770 23520 18776
rect 23480 18290 23508 18770
rect 23817 18524 24113 18544
rect 23873 18522 23897 18524
rect 23953 18522 23977 18524
rect 24033 18522 24057 18524
rect 23895 18470 23897 18522
rect 23959 18470 23971 18522
rect 24033 18470 24035 18522
rect 23873 18468 23897 18470
rect 23953 18468 23977 18470
rect 24033 18468 24057 18470
rect 23817 18448 24113 18468
rect 23468 18284 23520 18290
rect 23468 18226 23520 18232
rect 23558 18184 23614 18193
rect 23558 18119 23614 18128
rect 23652 18148 23704 18154
rect 23468 18080 23520 18086
rect 23468 18022 23520 18028
rect 23480 17377 23508 18022
rect 23466 17368 23522 17377
rect 23466 17303 23522 17312
rect 23572 17252 23600 18119
rect 23652 18090 23704 18096
rect 23480 17224 23600 17252
rect 23376 16992 23428 16998
rect 23376 16934 23428 16940
rect 23112 16102 23324 16130
rect 23006 15328 23062 15337
rect 23006 15263 23062 15272
rect 23008 14952 23060 14958
rect 23008 14894 23060 14900
rect 23020 14618 23048 14894
rect 23008 14612 23060 14618
rect 23008 14554 23060 14560
rect 23112 14498 23140 16102
rect 23284 16040 23336 16046
rect 23282 16008 23284 16017
rect 23336 16008 23338 16017
rect 23282 15943 23338 15952
rect 23192 14884 23244 14890
rect 23192 14826 23244 14832
rect 23204 14550 23232 14826
rect 22836 14470 23140 14498
rect 23192 14544 23244 14550
rect 23192 14486 23244 14492
rect 22836 12617 22864 14470
rect 22916 14408 22968 14414
rect 22914 14376 22916 14385
rect 23008 14408 23060 14414
rect 22968 14376 22970 14385
rect 23008 14350 23060 14356
rect 22914 14311 22970 14320
rect 22928 14074 22956 14311
rect 22916 14068 22968 14074
rect 22916 14010 22968 14016
rect 23020 13954 23048 14350
rect 23192 14272 23244 14278
rect 23192 14214 23244 14220
rect 22928 13926 23048 13954
rect 22928 13462 22956 13926
rect 23008 13864 23060 13870
rect 23204 13852 23232 14214
rect 23284 13864 23336 13870
rect 23204 13824 23284 13852
rect 23008 13806 23060 13812
rect 23284 13806 23336 13812
rect 22916 13456 22968 13462
rect 22916 13398 22968 13404
rect 23020 12782 23048 13806
rect 23192 13728 23244 13734
rect 23192 13670 23244 13676
rect 23100 13320 23152 13326
rect 23100 13262 23152 13268
rect 23112 12850 23140 13262
rect 23100 12844 23152 12850
rect 23100 12786 23152 12792
rect 23008 12776 23060 12782
rect 23008 12718 23060 12724
rect 22916 12708 22968 12714
rect 22916 12650 22968 12656
rect 22822 12608 22878 12617
rect 22822 12543 22878 12552
rect 22822 12472 22878 12481
rect 22928 12442 22956 12650
rect 22822 12407 22878 12416
rect 22916 12436 22968 12442
rect 22836 11778 22864 12407
rect 22916 12378 22968 12384
rect 23008 12368 23060 12374
rect 23008 12310 23060 12316
rect 23020 11898 23048 12310
rect 23008 11892 23060 11898
rect 23008 11834 23060 11840
rect 22836 11750 23048 11778
rect 23112 11762 23140 12786
rect 23204 12306 23232 13670
rect 23284 13524 23336 13530
rect 23284 13466 23336 13472
rect 23296 12714 23324 13466
rect 23284 12708 23336 12714
rect 23284 12650 23336 12656
rect 23282 12608 23338 12617
rect 23282 12543 23338 12552
rect 23192 12300 23244 12306
rect 23192 12242 23244 12248
rect 22732 11280 22784 11286
rect 22732 11222 22784 11228
rect 22640 11144 22692 11150
rect 22640 11086 22692 11092
rect 22546 10568 22602 10577
rect 22546 10503 22548 10512
rect 22600 10503 22602 10512
rect 22548 10474 22600 10480
rect 22652 10266 22680 11086
rect 22744 10810 22772 11222
rect 22916 11144 22968 11150
rect 22916 11086 22968 11092
rect 22732 10804 22784 10810
rect 22732 10746 22784 10752
rect 22640 10260 22692 10266
rect 22640 10202 22692 10208
rect 22454 10024 22510 10033
rect 22454 9959 22510 9968
rect 22640 9512 22692 9518
rect 22640 9454 22692 9460
rect 22652 8634 22680 9454
rect 22928 9110 22956 11086
rect 22916 9104 22968 9110
rect 22916 9046 22968 9052
rect 23020 8634 23048 11750
rect 23100 11756 23152 11762
rect 23100 11698 23152 11704
rect 23296 9058 23324 12543
rect 23388 12356 23416 16934
rect 23480 13433 23508 17224
rect 23664 16017 23692 18090
rect 24216 17746 24244 19071
rect 24296 18284 24348 18290
rect 24296 18226 24348 18232
rect 24204 17740 24256 17746
rect 24204 17682 24256 17688
rect 23817 17436 24113 17456
rect 23873 17434 23897 17436
rect 23953 17434 23977 17436
rect 24033 17434 24057 17436
rect 23895 17382 23897 17434
rect 23959 17382 23971 17434
rect 24033 17382 24035 17434
rect 23873 17380 23897 17382
rect 23953 17380 23977 17382
rect 24033 17380 24057 17382
rect 23817 17360 24113 17380
rect 24216 17338 24244 17682
rect 24204 17332 24256 17338
rect 24204 17274 24256 17280
rect 24308 17218 24336 18226
rect 24308 17190 24520 17218
rect 24386 17096 24442 17105
rect 24386 17031 24388 17040
rect 24440 17031 24442 17040
rect 24388 17002 24440 17008
rect 24296 16992 24348 16998
rect 24296 16934 24348 16940
rect 23744 16652 23796 16658
rect 23744 16594 23796 16600
rect 24204 16652 24256 16658
rect 24204 16594 24256 16600
rect 23650 16008 23706 16017
rect 23756 15978 23784 16594
rect 23817 16348 24113 16368
rect 23873 16346 23897 16348
rect 23953 16346 23977 16348
rect 24033 16346 24057 16348
rect 23895 16294 23897 16346
rect 23959 16294 23971 16346
rect 24033 16294 24035 16346
rect 23873 16292 23897 16294
rect 23953 16292 23977 16294
rect 24033 16292 24057 16294
rect 23817 16272 24113 16292
rect 23650 15943 23706 15952
rect 23744 15972 23796 15978
rect 23744 15914 23796 15920
rect 23560 15904 23612 15910
rect 23560 15846 23612 15852
rect 23466 13424 23522 13433
rect 23466 13359 23522 13368
rect 23572 12617 23600 15846
rect 23817 15260 24113 15280
rect 23873 15258 23897 15260
rect 23953 15258 23977 15260
rect 24033 15258 24057 15260
rect 23895 15206 23897 15258
rect 23959 15206 23971 15258
rect 24033 15206 24035 15258
rect 23873 15204 23897 15206
rect 23953 15204 23977 15206
rect 24033 15204 24057 15206
rect 23817 15184 24113 15204
rect 23652 14476 23704 14482
rect 23652 14418 23704 14424
rect 23664 14074 23692 14418
rect 23817 14172 24113 14192
rect 23873 14170 23897 14172
rect 23953 14170 23977 14172
rect 24033 14170 24057 14172
rect 23895 14118 23897 14170
rect 23959 14118 23971 14170
rect 24033 14118 24035 14170
rect 23873 14116 23897 14118
rect 23953 14116 23977 14118
rect 24033 14116 24057 14118
rect 23817 14096 24113 14116
rect 23652 14068 23704 14074
rect 23652 14010 23704 14016
rect 23664 12714 23692 14010
rect 24020 13864 24072 13870
rect 24216 13852 24244 16594
rect 24308 14929 24336 16934
rect 24388 16720 24440 16726
rect 24386 16688 24388 16697
rect 24440 16688 24442 16697
rect 24386 16623 24442 16632
rect 24492 16572 24520 17190
rect 24492 16544 24704 16572
rect 24572 15564 24624 15570
rect 24572 15506 24624 15512
rect 24294 14920 24350 14929
rect 24584 14890 24612 15506
rect 24294 14855 24350 14864
rect 24572 14884 24624 14890
rect 24572 14826 24624 14832
rect 24480 14816 24532 14822
rect 24480 14758 24532 14764
rect 24388 13864 24440 13870
rect 24216 13824 24388 13852
rect 24020 13806 24072 13812
rect 24388 13806 24440 13812
rect 24032 13569 24060 13806
rect 24492 13682 24520 14758
rect 24308 13654 24520 13682
rect 24018 13560 24074 13569
rect 24308 13530 24336 13654
rect 24478 13560 24534 13569
rect 24018 13495 24074 13504
rect 24296 13524 24348 13530
rect 24478 13495 24534 13504
rect 24296 13466 24348 13472
rect 24294 13424 24350 13433
rect 24204 13388 24256 13394
rect 24294 13359 24350 13368
rect 24204 13330 24256 13336
rect 23744 13320 23796 13326
rect 23744 13262 23796 13268
rect 23652 12708 23704 12714
rect 23652 12650 23704 12656
rect 23558 12608 23614 12617
rect 23756 12594 23784 13262
rect 23817 13084 24113 13104
rect 23873 13082 23897 13084
rect 23953 13082 23977 13084
rect 24033 13082 24057 13084
rect 23895 13030 23897 13082
rect 23959 13030 23971 13082
rect 24033 13030 24035 13082
rect 23873 13028 23897 13030
rect 23953 13028 23977 13030
rect 24033 13028 24057 13030
rect 23817 13008 24113 13028
rect 24216 12986 24244 13330
rect 24204 12980 24256 12986
rect 24204 12922 24256 12928
rect 23756 12566 23876 12594
rect 23558 12543 23614 12552
rect 23848 12374 23876 12566
rect 23836 12368 23888 12374
rect 23388 12328 23508 12356
rect 23480 12238 23508 12328
rect 24216 12356 24244 12922
rect 24308 12730 24336 13359
rect 24492 12753 24520 13495
rect 24584 12764 24612 14826
rect 24676 12889 24704 16544
rect 24756 15904 24808 15910
rect 24756 15846 24808 15852
rect 24768 15745 24796 15846
rect 24754 15736 24810 15745
rect 24754 15671 24810 15680
rect 24848 15496 24900 15502
rect 24848 15438 24900 15444
rect 24860 14464 24888 15438
rect 24952 15162 24980 25327
rect 25780 23633 25808 27520
rect 25766 23624 25822 23633
rect 25766 23559 25822 23568
rect 25030 21176 25086 21185
rect 25030 21111 25086 21120
rect 25044 19922 25072 21111
rect 25032 19916 25084 19922
rect 25032 19858 25084 19864
rect 25044 19310 25072 19858
rect 25032 19304 25084 19310
rect 25032 19246 25084 19252
rect 25492 19168 25544 19174
rect 25492 19110 25544 19116
rect 25032 18828 25084 18834
rect 25032 18770 25084 18776
rect 25044 18086 25072 18770
rect 25124 18216 25176 18222
rect 25122 18184 25124 18193
rect 25176 18184 25178 18193
rect 25122 18119 25178 18128
rect 25032 18080 25084 18086
rect 25032 18022 25084 18028
rect 25216 18080 25268 18086
rect 25216 18022 25268 18028
rect 25044 17105 25072 18022
rect 25030 17096 25086 17105
rect 25030 17031 25086 17040
rect 24940 15156 24992 15162
rect 24940 15098 24992 15104
rect 24952 14958 24980 15098
rect 24940 14952 24992 14958
rect 24940 14894 24992 14900
rect 24860 14436 24980 14464
rect 24846 14376 24902 14385
rect 24846 14311 24902 14320
rect 24662 12880 24718 12889
rect 24662 12815 24718 12824
rect 24478 12744 24534 12753
rect 24308 12702 24428 12730
rect 24296 12640 24348 12646
rect 24296 12582 24348 12588
rect 24308 12374 24336 12582
rect 23836 12310 23888 12316
rect 24124 12328 24244 12356
rect 24296 12368 24348 12374
rect 23468 12232 23520 12238
rect 23374 12200 23430 12209
rect 23468 12174 23520 12180
rect 23652 12232 23704 12238
rect 23652 12174 23704 12180
rect 23374 12135 23430 12144
rect 23388 9518 23416 12135
rect 23480 11354 23508 12174
rect 23560 12164 23612 12170
rect 23560 12106 23612 12112
rect 23572 11626 23600 12106
rect 23664 11801 23692 12174
rect 24124 12170 24152 12328
rect 24296 12310 24348 12316
rect 24400 12186 24428 12702
rect 24584 12736 24704 12764
rect 24478 12679 24534 12688
rect 24112 12164 24164 12170
rect 24112 12106 24164 12112
rect 24216 12158 24428 12186
rect 23817 11996 24113 12016
rect 23873 11994 23897 11996
rect 23953 11994 23977 11996
rect 24033 11994 24057 11996
rect 23895 11942 23897 11994
rect 23959 11942 23971 11994
rect 24033 11942 24035 11994
rect 23873 11940 23897 11942
rect 23953 11940 23977 11942
rect 24033 11940 24057 11942
rect 23817 11920 24113 11940
rect 23650 11792 23706 11801
rect 23650 11727 23652 11736
rect 23704 11727 23706 11736
rect 23652 11698 23704 11704
rect 23560 11620 23612 11626
rect 23560 11562 23612 11568
rect 23652 11620 23704 11626
rect 23652 11562 23704 11568
rect 23468 11348 23520 11354
rect 23468 11290 23520 11296
rect 23468 10124 23520 10130
rect 23468 10066 23520 10072
rect 23376 9512 23428 9518
rect 23376 9454 23428 9460
rect 23388 9110 23416 9454
rect 23480 9382 23508 10066
rect 23560 9920 23612 9926
rect 23560 9862 23612 9868
rect 23468 9376 23520 9382
rect 23468 9318 23520 9324
rect 23112 9030 23324 9058
rect 23376 9104 23428 9110
rect 23376 9046 23428 9052
rect 22640 8628 22692 8634
rect 22640 8570 22692 8576
rect 23008 8628 23060 8634
rect 23008 8570 23060 8576
rect 22456 8016 22508 8022
rect 22456 7958 22508 7964
rect 22364 7880 22416 7886
rect 21626 7848 21682 7857
rect 21364 7806 21484 7834
rect 21352 7744 21404 7750
rect 21350 7712 21352 7721
rect 21404 7712 21406 7721
rect 21350 7647 21406 7656
rect 21364 7546 21392 7647
rect 21352 7540 21404 7546
rect 21352 7482 21404 7488
rect 21258 7440 21314 7449
rect 21168 7404 21220 7410
rect 21258 7375 21314 7384
rect 21168 7346 21220 7352
rect 20984 7268 21036 7274
rect 20984 7210 21036 7216
rect 20892 6996 20944 7002
rect 20892 6938 20944 6944
rect 20616 6860 20668 6866
rect 20616 6802 20668 6808
rect 20996 6458 21024 7210
rect 21180 7002 21208 7346
rect 21168 6996 21220 7002
rect 21168 6938 21220 6944
rect 20984 6452 21036 6458
rect 20984 6394 21036 6400
rect 20984 6180 21036 6186
rect 20984 6122 21036 6128
rect 20800 6112 20852 6118
rect 20800 6054 20852 6060
rect 20616 5840 20668 5846
rect 20616 5782 20668 5788
rect 20706 5808 20762 5817
rect 20628 5681 20656 5782
rect 20706 5743 20708 5752
rect 20760 5743 20762 5752
rect 20708 5714 20760 5720
rect 20614 5672 20670 5681
rect 20614 5607 20670 5616
rect 20812 5370 20840 6054
rect 20996 5778 21024 6122
rect 20984 5772 21036 5778
rect 20984 5714 21036 5720
rect 20800 5364 20852 5370
rect 20800 5306 20852 5312
rect 20812 5098 20840 5306
rect 20800 5092 20852 5098
rect 20800 5034 20852 5040
rect 20812 4758 20840 5034
rect 20800 4752 20852 4758
rect 20800 4694 20852 4700
rect 20812 4214 20840 4694
rect 20800 4208 20852 4214
rect 20800 4150 20852 4156
rect 20524 3664 20576 3670
rect 20524 3606 20576 3612
rect 20432 3188 20484 3194
rect 20432 3130 20484 3136
rect 21272 2922 21300 7375
rect 21352 6792 21404 6798
rect 21352 6734 21404 6740
rect 21364 5846 21392 6734
rect 21352 5840 21404 5846
rect 21352 5782 21404 5788
rect 21350 4856 21406 4865
rect 21350 4791 21352 4800
rect 21404 4791 21406 4800
rect 21352 4762 21404 4768
rect 21364 4282 21392 4762
rect 21352 4276 21404 4282
rect 21352 4218 21404 4224
rect 21364 4010 21392 4218
rect 21456 4214 21484 7806
rect 22364 7822 22416 7828
rect 21626 7783 21682 7792
rect 21640 6934 21668 7783
rect 22376 7002 22404 7822
rect 22468 7546 22496 7958
rect 22548 7880 22600 7886
rect 22548 7822 22600 7828
rect 22456 7540 22508 7546
rect 22456 7482 22508 7488
rect 22560 7410 22588 7822
rect 22548 7404 22600 7410
rect 22548 7346 22600 7352
rect 22364 6996 22416 7002
rect 22364 6938 22416 6944
rect 22560 6934 22588 7346
rect 23112 6984 23140 9030
rect 23192 8968 23244 8974
rect 23192 8910 23244 8916
rect 23204 8673 23232 8910
rect 23480 8838 23508 9318
rect 23468 8832 23520 8838
rect 23468 8774 23520 8780
rect 23190 8664 23246 8673
rect 23190 8599 23246 8608
rect 23376 8628 23428 8634
rect 23204 8566 23232 8599
rect 23376 8570 23428 8576
rect 23192 8560 23244 8566
rect 23192 8502 23244 8508
rect 23282 8392 23338 8401
rect 23388 8362 23416 8570
rect 23282 8327 23284 8336
rect 23336 8327 23338 8336
rect 23376 8356 23428 8362
rect 23284 8298 23336 8304
rect 23376 8298 23428 8304
rect 23296 8090 23324 8298
rect 23284 8084 23336 8090
rect 23284 8026 23336 8032
rect 23192 7948 23244 7954
rect 23192 7890 23244 7896
rect 23204 7206 23232 7890
rect 23572 7528 23600 9862
rect 23296 7500 23600 7528
rect 23192 7200 23244 7206
rect 23192 7142 23244 7148
rect 23020 6956 23140 6984
rect 21628 6928 21680 6934
rect 21628 6870 21680 6876
rect 22548 6928 22600 6934
rect 22548 6870 22600 6876
rect 21640 5914 21668 6870
rect 21904 6112 21956 6118
rect 21904 6054 21956 6060
rect 22272 6112 22324 6118
rect 22272 6054 22324 6060
rect 21628 5908 21680 5914
rect 21628 5850 21680 5856
rect 21916 5846 21944 6054
rect 22284 5953 22312 6054
rect 22270 5944 22326 5953
rect 22326 5914 22496 5930
rect 22326 5908 22508 5914
rect 22326 5902 22456 5908
rect 22270 5879 22326 5888
rect 22456 5850 22508 5856
rect 21904 5840 21956 5846
rect 21904 5782 21956 5788
rect 23020 5710 23048 6956
rect 23098 6896 23154 6905
rect 23098 6831 23154 6840
rect 23112 6798 23140 6831
rect 23100 6792 23152 6798
rect 23100 6734 23152 6740
rect 23112 5778 23140 6734
rect 23192 6248 23244 6254
rect 23192 6190 23244 6196
rect 23204 5846 23232 6190
rect 23192 5840 23244 5846
rect 23190 5808 23192 5817
rect 23244 5808 23246 5817
rect 23100 5772 23152 5778
rect 23190 5743 23246 5752
rect 23100 5714 23152 5720
rect 22088 5704 22140 5710
rect 22088 5646 22140 5652
rect 23008 5704 23060 5710
rect 23008 5646 23060 5652
rect 21902 5128 21958 5137
rect 21902 5063 21958 5072
rect 21536 5024 21588 5030
rect 21536 4966 21588 4972
rect 21548 4321 21576 4966
rect 21720 4548 21772 4554
rect 21720 4490 21772 4496
rect 21534 4312 21590 4321
rect 21534 4247 21590 4256
rect 21444 4208 21496 4214
rect 21444 4150 21496 4156
rect 21352 4004 21404 4010
rect 21352 3946 21404 3952
rect 21456 3738 21484 4150
rect 21444 3732 21496 3738
rect 21444 3674 21496 3680
rect 21260 2916 21312 2922
rect 21260 2858 21312 2864
rect 20340 2508 20392 2514
rect 20340 2450 20392 2456
rect 18960 2304 19012 2310
rect 18960 2246 19012 2252
rect 19420 2304 19472 2310
rect 19420 2246 19472 2252
rect 20064 2304 20116 2310
rect 20064 2246 20116 2252
rect 19432 1057 19460 2246
rect 19602 1456 19658 1465
rect 19602 1391 19658 1400
rect 19418 1048 19474 1057
rect 19418 983 19474 992
rect 19616 480 19644 1391
rect 20076 921 20104 2246
rect 20706 1864 20762 1873
rect 20706 1799 20762 1808
rect 20062 912 20118 921
rect 20062 847 20118 856
rect 20720 480 20748 1799
rect 21732 480 21760 4490
rect 21916 4146 21944 5063
rect 22100 4826 22128 5646
rect 22916 5568 22968 5574
rect 22916 5510 22968 5516
rect 22178 5128 22234 5137
rect 22178 5063 22234 5072
rect 22088 4820 22140 4826
rect 22088 4762 22140 4768
rect 22192 4690 22220 5063
rect 22928 5012 22956 5510
rect 23190 5400 23246 5409
rect 23190 5335 23246 5344
rect 23204 5137 23232 5335
rect 23190 5128 23246 5137
rect 23190 5063 23246 5072
rect 23008 5024 23060 5030
rect 22928 4984 23008 5012
rect 23008 4966 23060 4972
rect 22180 4684 22232 4690
rect 22180 4626 22232 4632
rect 22086 4584 22142 4593
rect 22086 4519 22142 4528
rect 21904 4140 21956 4146
rect 21904 4082 21956 4088
rect 22100 3534 22128 4519
rect 23020 4457 23048 4966
rect 23192 4616 23244 4622
rect 23192 4558 23244 4564
rect 23006 4448 23062 4457
rect 23006 4383 23062 4392
rect 23204 4214 23232 4558
rect 23192 4208 23244 4214
rect 22730 4176 22786 4185
rect 23192 4150 23244 4156
rect 22730 4111 22786 4120
rect 22456 4004 22508 4010
rect 22456 3946 22508 3952
rect 22180 3664 22232 3670
rect 22180 3606 22232 3612
rect 22362 3632 22418 3641
rect 22088 3528 22140 3534
rect 22088 3470 22140 3476
rect 22100 3126 22128 3470
rect 22088 3120 22140 3126
rect 22088 3062 22140 3068
rect 22192 2854 22220 3606
rect 22362 3567 22418 3576
rect 22376 3534 22404 3567
rect 22468 3534 22496 3946
rect 22364 3528 22416 3534
rect 22364 3470 22416 3476
rect 22456 3528 22508 3534
rect 22456 3470 22508 3476
rect 22468 3058 22496 3470
rect 22456 3052 22508 3058
rect 22456 2994 22508 3000
rect 22180 2848 22232 2854
rect 22180 2790 22232 2796
rect 22272 2508 22324 2514
rect 22272 2450 22324 2456
rect 22284 2417 22312 2450
rect 22270 2408 22326 2417
rect 22270 2343 22326 2352
rect 22456 2304 22508 2310
rect 22456 2246 22508 2252
rect 22468 1465 22496 2246
rect 22454 1456 22510 1465
rect 22454 1391 22510 1400
rect 22744 480 22772 4111
rect 23296 4049 23324 7500
rect 23560 7404 23612 7410
rect 23560 7346 23612 7352
rect 23572 6798 23600 7346
rect 23664 6934 23692 11562
rect 23744 11552 23796 11558
rect 23744 11494 23796 11500
rect 23756 8945 23784 11494
rect 23817 10908 24113 10928
rect 23873 10906 23897 10908
rect 23953 10906 23977 10908
rect 24033 10906 24057 10908
rect 23895 10854 23897 10906
rect 23959 10854 23971 10906
rect 24033 10854 24035 10906
rect 23873 10852 23897 10854
rect 23953 10852 23977 10854
rect 24033 10852 24057 10854
rect 23817 10832 24113 10852
rect 24216 10849 24244 12158
rect 24296 12096 24348 12102
rect 24296 12038 24348 12044
rect 24308 11558 24336 12038
rect 24296 11552 24348 11558
rect 24296 11494 24348 11500
rect 24388 11552 24440 11558
rect 24388 11494 24440 11500
rect 24400 11098 24428 11494
rect 24492 11218 24520 12679
rect 24480 11212 24532 11218
rect 24480 11154 24532 11160
rect 24308 11070 24428 11098
rect 24202 10840 24258 10849
rect 24202 10775 24258 10784
rect 24112 10464 24164 10470
rect 24112 10406 24164 10412
rect 24124 10198 24152 10406
rect 24112 10192 24164 10198
rect 24164 10152 24244 10180
rect 24112 10134 24164 10140
rect 23817 9820 24113 9840
rect 23873 9818 23897 9820
rect 23953 9818 23977 9820
rect 24033 9818 24057 9820
rect 23895 9766 23897 9818
rect 23959 9766 23971 9818
rect 24033 9766 24035 9818
rect 23873 9764 23897 9766
rect 23953 9764 23977 9766
rect 24033 9764 24057 9766
rect 23817 9744 24113 9764
rect 23926 9480 23982 9489
rect 23926 9415 23928 9424
rect 23980 9415 23982 9424
rect 23928 9386 23980 9392
rect 24216 9178 24244 10152
rect 24308 9568 24336 11070
rect 24388 11008 24440 11014
rect 24388 10950 24440 10956
rect 24400 10742 24428 10950
rect 24492 10810 24520 11154
rect 24480 10804 24532 10810
rect 24480 10746 24532 10752
rect 24388 10736 24440 10742
rect 24386 10704 24388 10713
rect 24440 10704 24442 10713
rect 24386 10639 24442 10648
rect 24480 10464 24532 10470
rect 24480 10406 24532 10412
rect 24308 9540 24428 9568
rect 24296 9444 24348 9450
rect 24296 9386 24348 9392
rect 24204 9172 24256 9178
rect 24204 9114 24256 9120
rect 23742 8936 23798 8945
rect 23742 8871 23798 8880
rect 23817 8732 24113 8752
rect 23873 8730 23897 8732
rect 23953 8730 23977 8732
rect 24033 8730 24057 8732
rect 23895 8678 23897 8730
rect 23959 8678 23971 8730
rect 24033 8678 24035 8730
rect 23873 8676 23897 8678
rect 23953 8676 23977 8678
rect 24033 8676 24057 8678
rect 23817 8656 24113 8676
rect 24216 8634 24244 9114
rect 24308 9110 24336 9386
rect 24296 9104 24348 9110
rect 24296 9046 24348 9052
rect 24400 8956 24428 9540
rect 24308 8928 24428 8956
rect 24204 8628 24256 8634
rect 24204 8570 24256 8576
rect 24204 8492 24256 8498
rect 24204 8434 24256 8440
rect 23744 7880 23796 7886
rect 23744 7822 23796 7828
rect 23756 7449 23784 7822
rect 23817 7644 24113 7664
rect 23873 7642 23897 7644
rect 23953 7642 23977 7644
rect 24033 7642 24057 7644
rect 23895 7590 23897 7642
rect 23959 7590 23971 7642
rect 24033 7590 24035 7642
rect 23873 7588 23897 7590
rect 23953 7588 23977 7590
rect 24033 7588 24057 7590
rect 23817 7568 24113 7588
rect 23742 7440 23798 7449
rect 23742 7375 23798 7384
rect 23744 7200 23796 7206
rect 23744 7142 23796 7148
rect 23652 6928 23704 6934
rect 23652 6870 23704 6876
rect 23560 6792 23612 6798
rect 23558 6760 23560 6769
rect 23612 6760 23614 6769
rect 23558 6695 23614 6704
rect 23664 6458 23692 6870
rect 23652 6452 23704 6458
rect 23652 6394 23704 6400
rect 23756 6338 23784 7142
rect 23817 6556 24113 6576
rect 23873 6554 23897 6556
rect 23953 6554 23977 6556
rect 24033 6554 24057 6556
rect 23895 6502 23897 6554
rect 23959 6502 23971 6554
rect 24033 6502 24035 6554
rect 23873 6500 23897 6502
rect 23953 6500 23977 6502
rect 24033 6500 24057 6502
rect 23817 6480 24113 6500
rect 23664 6310 23784 6338
rect 23376 5228 23428 5234
rect 23376 5170 23428 5176
rect 23388 4826 23416 5170
rect 23664 4865 23692 6310
rect 23744 6112 23796 6118
rect 23744 6054 23796 6060
rect 23650 4856 23706 4865
rect 23376 4820 23428 4826
rect 23428 4780 23508 4808
rect 23650 4791 23706 4800
rect 23376 4762 23428 4768
rect 23480 4146 23508 4780
rect 23652 4752 23704 4758
rect 23650 4720 23652 4729
rect 23704 4720 23706 4729
rect 23650 4655 23706 4664
rect 23558 4312 23614 4321
rect 23664 4282 23692 4655
rect 23558 4247 23614 4256
rect 23652 4276 23704 4282
rect 23376 4140 23428 4146
rect 23376 4082 23428 4088
rect 23468 4140 23520 4146
rect 23468 4082 23520 4088
rect 23282 4040 23338 4049
rect 23388 4010 23416 4082
rect 23282 3975 23338 3984
rect 23376 4004 23428 4010
rect 23376 3946 23428 3952
rect 23192 3936 23244 3942
rect 23192 3878 23244 3884
rect 23204 3398 23232 3878
rect 23192 3392 23244 3398
rect 23192 3334 23244 3340
rect 23098 3224 23154 3233
rect 23098 3159 23154 3168
rect 23006 2952 23062 2961
rect 23006 2887 23008 2896
rect 23060 2887 23062 2896
rect 23008 2858 23060 2864
rect 22916 2848 22968 2854
rect 22968 2796 23048 2802
rect 22916 2790 23048 2796
rect 22928 2774 23048 2790
rect 23020 2582 23048 2774
rect 23008 2576 23060 2582
rect 23112 2553 23140 3159
rect 23008 2518 23060 2524
rect 23098 2544 23154 2553
rect 23098 2479 23154 2488
rect 23204 1193 23232 3334
rect 23388 1329 23416 3946
rect 23572 3738 23600 4247
rect 23652 4218 23704 4224
rect 23560 3732 23612 3738
rect 23560 3674 23612 3680
rect 23572 3346 23600 3674
rect 23652 3528 23704 3534
rect 23652 3470 23704 3476
rect 23480 3318 23600 3346
rect 23480 3126 23508 3318
rect 23664 3194 23692 3470
rect 23652 3188 23704 3194
rect 23652 3130 23704 3136
rect 23468 3120 23520 3126
rect 23468 3062 23520 3068
rect 23480 2650 23508 3062
rect 23560 2984 23612 2990
rect 23560 2926 23612 2932
rect 23468 2644 23520 2650
rect 23468 2586 23520 2592
rect 23572 1465 23600 2926
rect 23558 1456 23614 1465
rect 23558 1391 23614 1400
rect 23374 1320 23430 1329
rect 23374 1255 23430 1264
rect 23190 1184 23246 1193
rect 23190 1119 23246 1128
rect 23756 480 23784 6054
rect 23817 5468 24113 5488
rect 23873 5466 23897 5468
rect 23953 5466 23977 5468
rect 24033 5466 24057 5468
rect 23895 5414 23897 5466
rect 23959 5414 23971 5466
rect 24033 5414 24035 5466
rect 23873 5412 23897 5414
rect 23953 5412 23977 5414
rect 24033 5412 24057 5414
rect 23817 5392 24113 5412
rect 23817 4380 24113 4400
rect 23873 4378 23897 4380
rect 23953 4378 23977 4380
rect 24033 4378 24057 4380
rect 23895 4326 23897 4378
rect 23959 4326 23971 4378
rect 24033 4326 24035 4378
rect 23873 4324 23897 4326
rect 23953 4324 23977 4326
rect 24033 4324 24057 4326
rect 23817 4304 24113 4324
rect 23817 3292 24113 3312
rect 23873 3290 23897 3292
rect 23953 3290 23977 3292
rect 24033 3290 24057 3292
rect 23895 3238 23897 3290
rect 23959 3238 23971 3290
rect 24033 3238 24035 3290
rect 23873 3236 23897 3238
rect 23953 3236 23977 3238
rect 24033 3236 24057 3238
rect 23817 3216 24113 3236
rect 24216 2990 24244 8434
rect 24308 6633 24336 8928
rect 24492 8498 24520 10406
rect 24572 10056 24624 10062
rect 24572 9998 24624 10004
rect 24584 9450 24612 9998
rect 24572 9444 24624 9450
rect 24572 9386 24624 9392
rect 24480 8492 24532 8498
rect 24480 8434 24532 8440
rect 24676 7274 24704 12736
rect 24860 12306 24888 14311
rect 24848 12300 24900 12306
rect 24848 12242 24900 12248
rect 24860 11898 24888 12242
rect 24848 11892 24900 11898
rect 24848 11834 24900 11840
rect 24848 11688 24900 11694
rect 24846 11656 24848 11665
rect 24900 11656 24902 11665
rect 24952 11626 24980 14436
rect 25032 12776 25084 12782
rect 25032 12718 25084 12724
rect 25044 12442 25072 12718
rect 25032 12436 25084 12442
rect 25032 12378 25084 12384
rect 24846 11591 24902 11600
rect 24940 11620 24992 11626
rect 24940 11562 24992 11568
rect 24940 10600 24992 10606
rect 24940 10542 24992 10548
rect 24952 10441 24980 10542
rect 24938 10432 24994 10441
rect 24938 10367 24994 10376
rect 24756 10056 24808 10062
rect 24756 9998 24808 10004
rect 24768 9636 24796 9998
rect 24938 9752 24994 9761
rect 24938 9687 24994 9696
rect 24768 9608 24888 9636
rect 24860 9518 24888 9608
rect 24848 9512 24900 9518
rect 24846 9480 24848 9489
rect 24900 9480 24902 9489
rect 24846 9415 24902 9424
rect 24952 8634 24980 9687
rect 25228 9081 25256 18022
rect 25400 16652 25452 16658
rect 25400 16594 25452 16600
rect 25412 15910 25440 16594
rect 25400 15904 25452 15910
rect 25400 15846 25452 15852
rect 25308 14000 25360 14006
rect 25412 13977 25440 15846
rect 25308 13942 25360 13948
rect 25398 13968 25454 13977
rect 25214 9072 25270 9081
rect 25214 9007 25270 9016
rect 25124 8832 25176 8838
rect 25124 8774 25176 8780
rect 24940 8628 24992 8634
rect 24940 8570 24992 8576
rect 24754 8528 24810 8537
rect 24754 8463 24810 8472
rect 24768 8430 24796 8463
rect 24756 8424 24808 8430
rect 24756 8366 24808 8372
rect 24756 7336 24808 7342
rect 24754 7304 24756 7313
rect 24808 7304 24810 7313
rect 24664 7268 24716 7274
rect 24754 7239 24810 7248
rect 24664 7210 24716 7216
rect 24940 7200 24992 7206
rect 24940 7142 24992 7148
rect 24572 6860 24624 6866
rect 24572 6802 24624 6808
rect 24294 6624 24350 6633
rect 24294 6559 24350 6568
rect 24584 6497 24612 6802
rect 24570 6488 24626 6497
rect 24570 6423 24572 6432
rect 24624 6423 24626 6432
rect 24572 6394 24624 6400
rect 24756 6248 24808 6254
rect 24754 6216 24756 6225
rect 24808 6216 24810 6225
rect 24754 6151 24810 6160
rect 24480 5840 24532 5846
rect 24480 5782 24532 5788
rect 24296 5704 24348 5710
rect 24296 5646 24348 5652
rect 24308 5370 24336 5646
rect 24388 5636 24440 5642
rect 24388 5578 24440 5584
rect 24296 5364 24348 5370
rect 24296 5306 24348 5312
rect 24400 5250 24428 5578
rect 24492 5370 24520 5782
rect 24952 5681 24980 7142
rect 24938 5672 24994 5681
rect 24938 5607 24994 5616
rect 24480 5364 24532 5370
rect 24480 5306 24532 5312
rect 24308 5234 24428 5250
rect 24296 5228 24428 5234
rect 24348 5222 24428 5228
rect 25030 5264 25086 5273
rect 25030 5199 25086 5208
rect 24296 5170 24348 5176
rect 25044 5166 25072 5199
rect 25032 5160 25084 5166
rect 24846 5128 24902 5137
rect 24296 5092 24348 5098
rect 25032 5102 25084 5108
rect 24846 5063 24902 5072
rect 24296 5034 24348 5040
rect 24308 4622 24336 5034
rect 24296 4616 24348 4622
rect 24296 4558 24348 4564
rect 24204 2984 24256 2990
rect 24204 2926 24256 2932
rect 24308 2530 24336 4558
rect 24756 4072 24808 4078
rect 24756 4014 24808 4020
rect 24768 3505 24796 4014
rect 24754 3496 24810 3505
rect 24754 3431 24810 3440
rect 24308 2514 24428 2530
rect 24308 2508 24440 2514
rect 24308 2502 24388 2508
rect 24388 2450 24440 2456
rect 23817 2204 24113 2224
rect 23873 2202 23897 2204
rect 23953 2202 23977 2204
rect 24033 2202 24057 2204
rect 23895 2150 23897 2202
rect 23959 2150 23971 2202
rect 24033 2150 24035 2202
rect 23873 2148 23897 2150
rect 23953 2148 23977 2150
rect 24033 2148 24057 2150
rect 23817 2128 24113 2148
rect 24860 480 24888 5063
rect 24938 4584 24994 4593
rect 24938 4519 24994 4528
rect 24952 3942 24980 4519
rect 24940 3936 24992 3942
rect 24940 3878 24992 3884
rect 24938 3496 24994 3505
rect 24938 3431 24994 3440
rect 24952 3194 24980 3431
rect 24940 3188 24992 3194
rect 24940 3130 24992 3136
rect 25136 513 25164 8774
rect 25320 7721 25348 13942
rect 25398 13903 25454 13912
rect 25504 11801 25532 19110
rect 25490 11792 25546 11801
rect 25490 11727 25546 11736
rect 25306 7712 25362 7721
rect 25306 7647 25362 7656
rect 25860 6656 25912 6662
rect 25860 6598 25912 6604
rect 25216 5024 25268 5030
rect 25216 4966 25268 4972
rect 25228 4185 25256 4966
rect 25214 4176 25270 4185
rect 25214 4111 25270 4120
rect 25216 2984 25268 2990
rect 25216 2926 25268 2932
rect 25228 2650 25256 2926
rect 25216 2644 25268 2650
rect 25216 2586 25268 2592
rect 25122 504 25178 513
rect 6 0 62 480
rect 1018 0 1074 480
rect 2030 0 2086 480
rect 3042 0 3098 480
rect 4146 0 4202 480
rect 5158 0 5214 480
rect 6170 0 6226 480
rect 7182 0 7238 480
rect 8286 0 8342 480
rect 9298 0 9354 480
rect 10310 0 10366 480
rect 11322 0 11378 480
rect 12426 0 12482 480
rect 13438 0 13494 480
rect 14450 0 14506 480
rect 15462 0 15518 480
rect 16566 0 16622 480
rect 17578 0 17634 480
rect 18590 0 18646 480
rect 19602 0 19658 480
rect 20706 0 20762 480
rect 21718 0 21774 480
rect 22730 0 22786 480
rect 23742 0 23798 480
rect 24846 0 24902 480
rect 25872 480 25900 6598
rect 26870 1728 26926 1737
rect 26870 1663 26926 1672
rect 26884 480 26912 1663
rect 25122 439 25178 448
rect 25858 0 25914 480
rect 26870 0 26926 480
<< via2 >>
rect 1018 14320 1074 14376
rect 5150 25050 5206 25052
rect 5230 25050 5286 25052
rect 5310 25050 5366 25052
rect 5390 25050 5446 25052
rect 5150 24998 5176 25050
rect 5176 24998 5206 25050
rect 5230 24998 5240 25050
rect 5240 24998 5286 25050
rect 5310 24998 5356 25050
rect 5356 24998 5366 25050
rect 5390 24998 5420 25050
rect 5420 24998 5446 25050
rect 5150 24996 5206 24998
rect 5230 24996 5286 24998
rect 5310 24996 5366 24998
rect 5390 24996 5446 24998
rect 5150 23962 5206 23964
rect 5230 23962 5286 23964
rect 5310 23962 5366 23964
rect 5390 23962 5446 23964
rect 5150 23910 5176 23962
rect 5176 23910 5206 23962
rect 5230 23910 5240 23962
rect 5240 23910 5286 23962
rect 5310 23910 5356 23962
rect 5356 23910 5366 23962
rect 5390 23910 5420 23962
rect 5420 23910 5446 23962
rect 5150 23908 5206 23910
rect 5230 23908 5286 23910
rect 5310 23908 5366 23910
rect 5390 23908 5446 23910
rect 5150 22874 5206 22876
rect 5230 22874 5286 22876
rect 5310 22874 5366 22876
rect 5390 22874 5446 22876
rect 5150 22822 5176 22874
rect 5176 22822 5206 22874
rect 5230 22822 5240 22874
rect 5240 22822 5286 22874
rect 5310 22822 5356 22874
rect 5356 22822 5366 22874
rect 5390 22822 5420 22874
rect 5420 22822 5446 22874
rect 5150 22820 5206 22822
rect 5230 22820 5286 22822
rect 5310 22820 5366 22822
rect 5390 22820 5446 22822
rect 5150 21786 5206 21788
rect 5230 21786 5286 21788
rect 5310 21786 5366 21788
rect 5390 21786 5446 21788
rect 5150 21734 5176 21786
rect 5176 21734 5206 21786
rect 5230 21734 5240 21786
rect 5240 21734 5286 21786
rect 5310 21734 5356 21786
rect 5356 21734 5366 21786
rect 5390 21734 5420 21786
rect 5420 21734 5446 21786
rect 5150 21732 5206 21734
rect 5230 21732 5286 21734
rect 5310 21732 5366 21734
rect 5390 21732 5446 21734
rect 5150 20698 5206 20700
rect 5230 20698 5286 20700
rect 5310 20698 5366 20700
rect 5390 20698 5446 20700
rect 5150 20646 5176 20698
rect 5176 20646 5206 20698
rect 5230 20646 5240 20698
rect 5240 20646 5286 20698
rect 5310 20646 5356 20698
rect 5356 20646 5366 20698
rect 5390 20646 5420 20698
rect 5420 20646 5446 20698
rect 5150 20644 5206 20646
rect 5230 20644 5286 20646
rect 5310 20644 5366 20646
rect 5390 20644 5446 20646
rect 5150 19610 5206 19612
rect 5230 19610 5286 19612
rect 5310 19610 5366 19612
rect 5390 19610 5446 19612
rect 5150 19558 5176 19610
rect 5176 19558 5206 19610
rect 5230 19558 5240 19610
rect 5240 19558 5286 19610
rect 5310 19558 5356 19610
rect 5356 19558 5366 19610
rect 5390 19558 5420 19610
rect 5420 19558 5446 19610
rect 5150 19556 5206 19558
rect 5230 19556 5286 19558
rect 5310 19556 5366 19558
rect 5390 19556 5446 19558
rect 5150 18522 5206 18524
rect 5230 18522 5286 18524
rect 5310 18522 5366 18524
rect 5390 18522 5446 18524
rect 5150 18470 5176 18522
rect 5176 18470 5206 18522
rect 5230 18470 5240 18522
rect 5240 18470 5286 18522
rect 5310 18470 5356 18522
rect 5356 18470 5366 18522
rect 5390 18470 5420 18522
rect 5420 18470 5446 18522
rect 5150 18468 5206 18470
rect 5230 18468 5286 18470
rect 5310 18468 5366 18470
rect 5390 18468 5446 18470
rect 9817 25594 9873 25596
rect 9897 25594 9953 25596
rect 9977 25594 10033 25596
rect 10057 25594 10113 25596
rect 9817 25542 9843 25594
rect 9843 25542 9873 25594
rect 9897 25542 9907 25594
rect 9907 25542 9953 25594
rect 9977 25542 10023 25594
rect 10023 25542 10033 25594
rect 10057 25542 10087 25594
rect 10087 25542 10113 25594
rect 9817 25540 9873 25542
rect 9897 25540 9953 25542
rect 9977 25540 10033 25542
rect 10057 25540 10113 25542
rect 9817 24506 9873 24508
rect 9897 24506 9953 24508
rect 9977 24506 10033 24508
rect 10057 24506 10113 24508
rect 9817 24454 9843 24506
rect 9843 24454 9873 24506
rect 9897 24454 9907 24506
rect 9907 24454 9953 24506
rect 9977 24454 10023 24506
rect 10023 24454 10033 24506
rect 10057 24454 10087 24506
rect 10087 24454 10113 24506
rect 9817 24452 9873 24454
rect 9897 24452 9953 24454
rect 9977 24452 10033 24454
rect 10057 24452 10113 24454
rect 9817 23418 9873 23420
rect 9897 23418 9953 23420
rect 9977 23418 10033 23420
rect 10057 23418 10113 23420
rect 9817 23366 9843 23418
rect 9843 23366 9873 23418
rect 9897 23366 9907 23418
rect 9907 23366 9953 23418
rect 9977 23366 10023 23418
rect 10023 23366 10033 23418
rect 10057 23366 10087 23418
rect 10087 23366 10113 23418
rect 9817 23364 9873 23366
rect 9897 23364 9953 23366
rect 9977 23364 10033 23366
rect 10057 23364 10113 23366
rect 9817 22330 9873 22332
rect 9897 22330 9953 22332
rect 9977 22330 10033 22332
rect 10057 22330 10113 22332
rect 9817 22278 9843 22330
rect 9843 22278 9873 22330
rect 9897 22278 9907 22330
rect 9907 22278 9953 22330
rect 9977 22278 10023 22330
rect 10023 22278 10033 22330
rect 10057 22278 10087 22330
rect 10087 22278 10113 22330
rect 9817 22276 9873 22278
rect 9897 22276 9953 22278
rect 9977 22276 10033 22278
rect 10057 22276 10113 22278
rect 9817 21242 9873 21244
rect 9897 21242 9953 21244
rect 9977 21242 10033 21244
rect 10057 21242 10113 21244
rect 9817 21190 9843 21242
rect 9843 21190 9873 21242
rect 9897 21190 9907 21242
rect 9907 21190 9953 21242
rect 9977 21190 10023 21242
rect 10023 21190 10033 21242
rect 10057 21190 10087 21242
rect 10087 21190 10113 21242
rect 9817 21188 9873 21190
rect 9897 21188 9953 21190
rect 9977 21188 10033 21190
rect 10057 21188 10113 21190
rect 9817 20154 9873 20156
rect 9897 20154 9953 20156
rect 9977 20154 10033 20156
rect 10057 20154 10113 20156
rect 9817 20102 9843 20154
rect 9843 20102 9873 20154
rect 9897 20102 9907 20154
rect 9907 20102 9953 20154
rect 9977 20102 10023 20154
rect 10023 20102 10033 20154
rect 10057 20102 10087 20154
rect 10087 20102 10113 20154
rect 9817 20100 9873 20102
rect 9897 20100 9953 20102
rect 9977 20100 10033 20102
rect 10057 20100 10113 20102
rect 9817 19066 9873 19068
rect 9897 19066 9953 19068
rect 9977 19066 10033 19068
rect 10057 19066 10113 19068
rect 9817 19014 9843 19066
rect 9843 19014 9873 19066
rect 9897 19014 9907 19066
rect 9907 19014 9953 19066
rect 9977 19014 10023 19066
rect 10023 19014 10033 19066
rect 10057 19014 10087 19066
rect 10087 19014 10113 19066
rect 9817 19012 9873 19014
rect 9897 19012 9953 19014
rect 9977 19012 10033 19014
rect 10057 19012 10113 19014
rect 10402 18672 10458 18728
rect 8286 17992 8342 18048
rect 9574 17992 9630 18048
rect 5150 17434 5206 17436
rect 5230 17434 5286 17436
rect 5310 17434 5366 17436
rect 5390 17434 5446 17436
rect 5150 17382 5176 17434
rect 5176 17382 5206 17434
rect 5230 17382 5240 17434
rect 5240 17382 5286 17434
rect 5310 17382 5356 17434
rect 5356 17382 5366 17434
rect 5390 17382 5420 17434
rect 5420 17382 5446 17434
rect 5150 17380 5206 17382
rect 5230 17380 5286 17382
rect 5310 17380 5366 17382
rect 5390 17380 5446 17382
rect 5150 16346 5206 16348
rect 5230 16346 5286 16348
rect 5310 16346 5366 16348
rect 5390 16346 5446 16348
rect 5150 16294 5176 16346
rect 5176 16294 5206 16346
rect 5230 16294 5240 16346
rect 5240 16294 5286 16346
rect 5310 16294 5356 16346
rect 5356 16294 5366 16346
rect 5390 16294 5420 16346
rect 5420 16294 5446 16346
rect 5150 16292 5206 16294
rect 5230 16292 5286 16294
rect 5310 16292 5366 16294
rect 5390 16292 5446 16294
rect 5526 16088 5582 16144
rect 5150 15258 5206 15260
rect 5230 15258 5286 15260
rect 5310 15258 5366 15260
rect 5390 15258 5446 15260
rect 5150 15206 5176 15258
rect 5176 15206 5206 15258
rect 5230 15206 5240 15258
rect 5240 15206 5286 15258
rect 5310 15206 5356 15258
rect 5356 15206 5366 15258
rect 5390 15206 5420 15258
rect 5420 15206 5446 15258
rect 5150 15204 5206 15206
rect 5230 15204 5286 15206
rect 5310 15204 5366 15206
rect 5390 15204 5446 15206
rect 5150 14170 5206 14172
rect 5230 14170 5286 14172
rect 5310 14170 5366 14172
rect 5390 14170 5446 14172
rect 5150 14118 5176 14170
rect 5176 14118 5206 14170
rect 5230 14118 5240 14170
rect 5240 14118 5286 14170
rect 5310 14118 5356 14170
rect 5356 14118 5366 14170
rect 5390 14118 5420 14170
rect 5420 14118 5446 14170
rect 5150 14116 5206 14118
rect 5230 14116 5286 14118
rect 5310 14116 5366 14118
rect 5390 14116 5446 14118
rect 5150 13082 5206 13084
rect 5230 13082 5286 13084
rect 5310 13082 5366 13084
rect 5390 13082 5446 13084
rect 5150 13030 5176 13082
rect 5176 13030 5206 13082
rect 5230 13030 5240 13082
rect 5240 13030 5286 13082
rect 5310 13030 5356 13082
rect 5356 13030 5366 13082
rect 5390 13030 5420 13082
rect 5420 13030 5446 13082
rect 5150 13028 5206 13030
rect 5230 13028 5286 13030
rect 5310 13028 5366 13030
rect 5390 13028 5446 13030
rect 5066 12688 5122 12744
rect 3686 11192 3742 11248
rect 4422 10512 4478 10568
rect 3318 8200 3374 8256
rect 1662 7112 1718 7168
rect 6 3712 62 3768
rect 1018 2896 1074 2952
rect 2766 6976 2822 7032
rect 2030 2760 2086 2816
rect 2122 1672 2178 1728
rect 3042 1944 3098 2000
rect 3226 1672 3282 1728
rect 2858 1400 2914 1456
rect 3778 6704 3834 6760
rect 3410 4800 3466 4856
rect 3594 3984 3650 4040
rect 4054 6432 4110 6488
rect 3962 3596 4018 3632
rect 3962 3576 3964 3596
rect 3964 3576 4016 3596
rect 4016 3576 4018 3596
rect 4974 4548 5030 4584
rect 4974 4528 4976 4548
rect 4976 4528 5028 4548
rect 5028 4528 5030 4548
rect 4606 3440 4662 3496
rect 4238 2932 4240 2952
rect 4240 2932 4292 2952
rect 4292 2932 4294 2952
rect 4238 2896 4294 2932
rect 4330 2760 4386 2816
rect 4514 2644 4570 2680
rect 4514 2624 4516 2644
rect 4516 2624 4568 2644
rect 4568 2624 4570 2644
rect 5150 11994 5206 11996
rect 5230 11994 5286 11996
rect 5310 11994 5366 11996
rect 5390 11994 5446 11996
rect 5150 11942 5176 11994
rect 5176 11942 5206 11994
rect 5230 11942 5240 11994
rect 5240 11942 5286 11994
rect 5310 11942 5356 11994
rect 5356 11942 5366 11994
rect 5390 11942 5420 11994
rect 5420 11942 5446 11994
rect 5150 11940 5206 11942
rect 5230 11940 5286 11942
rect 5310 11940 5366 11942
rect 5390 11940 5446 11942
rect 5150 10906 5206 10908
rect 5230 10906 5286 10908
rect 5310 10906 5366 10908
rect 5390 10906 5446 10908
rect 5150 10854 5176 10906
rect 5176 10854 5206 10906
rect 5230 10854 5240 10906
rect 5240 10854 5286 10906
rect 5310 10854 5356 10906
rect 5356 10854 5366 10906
rect 5390 10854 5420 10906
rect 5420 10854 5446 10906
rect 5150 10852 5206 10854
rect 5230 10852 5286 10854
rect 5310 10852 5366 10854
rect 5390 10852 5446 10854
rect 5150 9818 5206 9820
rect 5230 9818 5286 9820
rect 5310 9818 5366 9820
rect 5390 9818 5446 9820
rect 5150 9766 5176 9818
rect 5176 9766 5206 9818
rect 5230 9766 5240 9818
rect 5240 9766 5286 9818
rect 5310 9766 5356 9818
rect 5356 9766 5366 9818
rect 5390 9766 5420 9818
rect 5420 9766 5446 9818
rect 5150 9764 5206 9766
rect 5230 9764 5286 9766
rect 5310 9764 5366 9766
rect 5390 9764 5446 9766
rect 5150 8730 5206 8732
rect 5230 8730 5286 8732
rect 5310 8730 5366 8732
rect 5390 8730 5446 8732
rect 5150 8678 5176 8730
rect 5176 8678 5206 8730
rect 5230 8678 5240 8730
rect 5240 8678 5286 8730
rect 5310 8678 5356 8730
rect 5356 8678 5366 8730
rect 5390 8678 5420 8730
rect 5420 8678 5446 8730
rect 5150 8676 5206 8678
rect 5230 8676 5286 8678
rect 5310 8676 5366 8678
rect 5390 8676 5446 8678
rect 5150 7642 5206 7644
rect 5230 7642 5286 7644
rect 5310 7642 5366 7644
rect 5390 7642 5446 7644
rect 5150 7590 5176 7642
rect 5176 7590 5206 7642
rect 5230 7590 5240 7642
rect 5240 7590 5286 7642
rect 5310 7590 5356 7642
rect 5356 7590 5366 7642
rect 5390 7590 5420 7642
rect 5420 7590 5446 7642
rect 5150 7588 5206 7590
rect 5230 7588 5286 7590
rect 5310 7588 5366 7590
rect 5390 7588 5446 7590
rect 5150 6554 5206 6556
rect 5230 6554 5286 6556
rect 5310 6554 5366 6556
rect 5390 6554 5446 6556
rect 5150 6502 5176 6554
rect 5176 6502 5206 6554
rect 5230 6502 5240 6554
rect 5240 6502 5286 6554
rect 5310 6502 5356 6554
rect 5356 6502 5366 6554
rect 5390 6502 5420 6554
rect 5420 6502 5446 6554
rect 5150 6500 5206 6502
rect 5230 6500 5286 6502
rect 5310 6500 5366 6502
rect 5390 6500 5446 6502
rect 5150 5466 5206 5468
rect 5230 5466 5286 5468
rect 5310 5466 5366 5468
rect 5390 5466 5446 5468
rect 5150 5414 5176 5466
rect 5176 5414 5206 5466
rect 5230 5414 5240 5466
rect 5240 5414 5286 5466
rect 5310 5414 5356 5466
rect 5356 5414 5366 5466
rect 5390 5414 5420 5466
rect 5420 5414 5446 5466
rect 5150 5412 5206 5414
rect 5230 5412 5286 5414
rect 5310 5412 5366 5414
rect 5390 5412 5446 5414
rect 5150 4378 5206 4380
rect 5230 4378 5286 4380
rect 5310 4378 5366 4380
rect 5390 4378 5446 4380
rect 5150 4326 5176 4378
rect 5176 4326 5206 4378
rect 5230 4326 5240 4378
rect 5240 4326 5286 4378
rect 5310 4326 5356 4378
rect 5356 4326 5366 4378
rect 5390 4326 5420 4378
rect 5420 4326 5446 4378
rect 5150 4324 5206 4326
rect 5230 4324 5286 4326
rect 5310 4324 5366 4326
rect 5390 4324 5446 4326
rect 8194 15408 8250 15464
rect 7734 12008 7790 12064
rect 8102 11212 8158 11248
rect 8102 11192 8104 11212
rect 8104 11192 8156 11212
rect 8156 11192 8158 11212
rect 7366 10784 7422 10840
rect 9817 17978 9873 17980
rect 9897 17978 9953 17980
rect 9977 17978 10033 17980
rect 10057 17978 10113 17980
rect 9817 17926 9843 17978
rect 9843 17926 9873 17978
rect 9897 17926 9907 17978
rect 9907 17926 9953 17978
rect 9977 17926 10023 17978
rect 10023 17926 10033 17978
rect 10057 17926 10087 17978
rect 10087 17926 10113 17978
rect 9817 17924 9873 17926
rect 9897 17924 9953 17926
rect 9977 17924 10033 17926
rect 10057 17924 10113 17926
rect 9817 16890 9873 16892
rect 9897 16890 9953 16892
rect 9977 16890 10033 16892
rect 10057 16890 10113 16892
rect 9817 16838 9843 16890
rect 9843 16838 9873 16890
rect 9897 16838 9907 16890
rect 9907 16838 9953 16890
rect 9977 16838 10023 16890
rect 10023 16838 10033 16890
rect 10057 16838 10087 16890
rect 10087 16838 10113 16890
rect 9817 16836 9873 16838
rect 9897 16836 9953 16838
rect 9977 16836 10033 16838
rect 10057 16836 10113 16838
rect 9817 15802 9873 15804
rect 9897 15802 9953 15804
rect 9977 15802 10033 15804
rect 10057 15802 10113 15804
rect 9817 15750 9843 15802
rect 9843 15750 9873 15802
rect 9897 15750 9907 15802
rect 9907 15750 9953 15802
rect 9977 15750 10023 15802
rect 10023 15750 10033 15802
rect 10057 15750 10087 15802
rect 10087 15750 10113 15802
rect 9817 15748 9873 15750
rect 9897 15748 9953 15750
rect 9977 15748 10033 15750
rect 10057 15748 10113 15750
rect 9817 14714 9873 14716
rect 9897 14714 9953 14716
rect 9977 14714 10033 14716
rect 10057 14714 10113 14716
rect 9817 14662 9843 14714
rect 9843 14662 9873 14714
rect 9897 14662 9907 14714
rect 9907 14662 9953 14714
rect 9977 14662 10023 14714
rect 10023 14662 10033 14714
rect 10057 14662 10087 14714
rect 10087 14662 10113 14714
rect 9817 14660 9873 14662
rect 9897 14660 9953 14662
rect 9977 14660 10033 14662
rect 10057 14660 10113 14662
rect 8930 14320 8986 14376
rect 9817 13626 9873 13628
rect 9897 13626 9953 13628
rect 9977 13626 10033 13628
rect 10057 13626 10113 13628
rect 9817 13574 9843 13626
rect 9843 13574 9873 13626
rect 9897 13574 9907 13626
rect 9907 13574 9953 13626
rect 9977 13574 10023 13626
rect 10023 13574 10033 13626
rect 10057 13574 10087 13626
rect 10087 13574 10113 13626
rect 9817 13572 9873 13574
rect 9897 13572 9953 13574
rect 9977 13572 10033 13574
rect 10057 13572 10113 13574
rect 9482 12960 9538 13016
rect 8654 11892 8710 11928
rect 8654 11872 8656 11892
rect 8656 11872 8708 11892
rect 8708 11872 8710 11892
rect 8286 11736 8342 11792
rect 8286 11076 8342 11112
rect 8286 11056 8288 11076
rect 8288 11056 8340 11076
rect 8340 11056 8342 11076
rect 9817 12538 9873 12540
rect 9897 12538 9953 12540
rect 9977 12538 10033 12540
rect 10057 12538 10113 12540
rect 9817 12486 9843 12538
rect 9843 12486 9873 12538
rect 9897 12486 9907 12538
rect 9907 12486 9953 12538
rect 9977 12486 10023 12538
rect 10023 12486 10033 12538
rect 10057 12486 10087 12538
rect 10087 12486 10113 12538
rect 9817 12484 9873 12486
rect 9897 12484 9953 12486
rect 9977 12484 10033 12486
rect 10057 12484 10113 12486
rect 9390 12280 9446 12336
rect 8470 10684 8472 10704
rect 8472 10684 8524 10704
rect 8524 10684 8526 10704
rect 8470 10648 8526 10684
rect 8378 9832 8434 9888
rect 6446 9016 6502 9072
rect 5986 8880 6042 8936
rect 5802 8744 5858 8800
rect 5150 3290 5206 3292
rect 5230 3290 5286 3292
rect 5310 3290 5366 3292
rect 5390 3290 5446 3292
rect 5150 3238 5176 3290
rect 5176 3238 5206 3290
rect 5230 3238 5240 3290
rect 5240 3238 5286 3290
rect 5310 3238 5356 3290
rect 5356 3238 5366 3290
rect 5390 3238 5420 3290
rect 5420 3238 5446 3290
rect 5150 3236 5206 3238
rect 5230 3236 5286 3238
rect 5310 3236 5366 3238
rect 5390 3236 5446 3238
rect 4882 3032 4938 3088
rect 5342 2388 5344 2408
rect 5344 2388 5396 2408
rect 5396 2388 5398 2408
rect 5342 2352 5398 2388
rect 5150 2202 5206 2204
rect 5230 2202 5286 2204
rect 5310 2202 5366 2204
rect 5390 2202 5446 2204
rect 5150 2150 5176 2202
rect 5176 2150 5206 2202
rect 5230 2150 5240 2202
rect 5240 2150 5286 2202
rect 5310 2150 5356 2202
rect 5356 2150 5366 2202
rect 5390 2150 5420 2202
rect 5420 2150 5446 2202
rect 5150 2148 5206 2150
rect 5230 2148 5286 2150
rect 5310 2148 5366 2150
rect 5390 2148 5446 2150
rect 5710 3712 5766 3768
rect 5802 3188 5858 3224
rect 5802 3168 5804 3188
rect 5804 3168 5856 3188
rect 5856 3168 5858 3188
rect 6446 6976 6502 7032
rect 6538 6452 6594 6488
rect 6538 6432 6540 6452
rect 6540 6432 6592 6452
rect 6592 6432 6594 6452
rect 6078 3732 6134 3768
rect 6078 3712 6080 3732
rect 6080 3712 6132 3732
rect 6132 3712 6134 3732
rect 5894 2760 5950 2816
rect 5802 1808 5858 1864
rect 5618 992 5674 1048
rect 6446 5364 6502 5400
rect 6446 5344 6448 5364
rect 6448 5344 6500 5364
rect 6500 5344 6502 5364
rect 6538 5228 6594 5264
rect 6538 5208 6540 5228
rect 6540 5208 6592 5228
rect 6592 5208 6594 5228
rect 6538 4120 6594 4176
rect 6906 3304 6962 3360
rect 7182 2932 7184 2952
rect 7184 2932 7236 2952
rect 7236 2932 7238 2952
rect 7182 2896 7238 2932
rect 7182 2760 7238 2816
rect 6722 2488 6778 2544
rect 8378 9560 8434 9616
rect 7826 9424 7882 9480
rect 7734 7792 7790 7848
rect 8194 7948 8250 7984
rect 8194 7928 8196 7948
rect 8196 7928 8248 7948
rect 8248 7928 8250 7948
rect 8286 7828 8288 7848
rect 8288 7828 8340 7848
rect 8340 7828 8342 7848
rect 8286 7792 8342 7828
rect 8102 7248 8158 7304
rect 7826 7112 7882 7168
rect 8102 6316 8158 6352
rect 8102 6296 8104 6316
rect 8104 6296 8156 6316
rect 8156 6296 8158 6316
rect 7734 6180 7790 6216
rect 7734 6160 7736 6180
rect 7736 6160 7788 6180
rect 7788 6160 7790 6180
rect 8194 5772 8250 5808
rect 8194 5752 8196 5772
rect 8196 5752 8248 5772
rect 8248 5752 8250 5772
rect 7734 5636 7790 5672
rect 7734 5616 7736 5636
rect 7736 5616 7788 5636
rect 7788 5616 7790 5636
rect 8194 5092 8250 5128
rect 8194 5072 8196 5092
rect 8196 5072 8248 5092
rect 8248 5072 8250 5092
rect 8102 4392 8158 4448
rect 8930 8356 8986 8392
rect 8930 8336 8932 8356
rect 8932 8336 8984 8356
rect 8984 8336 8986 8356
rect 8654 7656 8710 7712
rect 8470 3984 8526 4040
rect 7550 1536 7606 1592
rect 7734 2760 7790 2816
rect 7642 856 7698 912
rect 9817 11450 9873 11452
rect 9897 11450 9953 11452
rect 9977 11450 10033 11452
rect 10057 11450 10113 11452
rect 9817 11398 9843 11450
rect 9843 11398 9873 11450
rect 9897 11398 9907 11450
rect 9907 11398 9953 11450
rect 9977 11398 10023 11450
rect 10023 11398 10033 11450
rect 10057 11398 10087 11450
rect 10087 11398 10113 11450
rect 9817 11396 9873 11398
rect 9897 11396 9953 11398
rect 9977 11396 10033 11398
rect 10057 11396 10113 11398
rect 9482 10104 9538 10160
rect 9817 10362 9873 10364
rect 9897 10362 9953 10364
rect 9977 10362 10033 10364
rect 10057 10362 10113 10364
rect 9817 10310 9843 10362
rect 9843 10310 9873 10362
rect 9897 10310 9907 10362
rect 9907 10310 9953 10362
rect 9977 10310 10023 10362
rect 10023 10310 10033 10362
rect 10057 10310 10087 10362
rect 10087 10310 10113 10362
rect 9817 10308 9873 10310
rect 9897 10308 9953 10310
rect 9977 10308 10033 10310
rect 10057 10308 10113 10310
rect 9666 9968 9722 10024
rect 11598 17040 11654 17096
rect 10678 11464 10734 11520
rect 10678 10512 10734 10568
rect 9666 9696 9722 9752
rect 9482 8200 9538 8256
rect 9298 7384 9354 7440
rect 8838 3052 8894 3088
rect 8838 3032 8840 3052
rect 8840 3032 8892 3052
rect 8892 3032 8894 3052
rect 8746 2252 8748 2272
rect 8748 2252 8800 2272
rect 8800 2252 8802 2272
rect 8746 2216 8802 2252
rect 9574 4800 9630 4856
rect 9482 4684 9538 4720
rect 9482 4664 9484 4684
rect 9484 4664 9536 4684
rect 9536 4664 9538 4684
rect 9114 4256 9170 4312
rect 9022 3984 9078 4040
rect 9298 4120 9354 4176
rect 9574 4120 9630 4176
rect 9817 9274 9873 9276
rect 9897 9274 9953 9276
rect 9977 9274 10033 9276
rect 10057 9274 10113 9276
rect 9817 9222 9843 9274
rect 9843 9222 9873 9274
rect 9897 9222 9907 9274
rect 9907 9222 9953 9274
rect 9977 9222 10023 9274
rect 10023 9222 10033 9274
rect 10057 9222 10087 9274
rect 10087 9222 10113 9274
rect 9817 9220 9873 9222
rect 9897 9220 9953 9222
rect 9977 9220 10033 9222
rect 10057 9220 10113 9222
rect 9817 8186 9873 8188
rect 9897 8186 9953 8188
rect 9977 8186 10033 8188
rect 10057 8186 10113 8188
rect 9817 8134 9843 8186
rect 9843 8134 9873 8186
rect 9897 8134 9907 8186
rect 9907 8134 9953 8186
rect 9977 8134 10023 8186
rect 10023 8134 10033 8186
rect 10057 8134 10087 8186
rect 10087 8134 10113 8186
rect 9817 8132 9873 8134
rect 9897 8132 9953 8134
rect 9977 8132 10033 8134
rect 10057 8132 10113 8134
rect 10218 8064 10274 8120
rect 10218 7656 10274 7712
rect 10402 8608 10458 8664
rect 9817 7098 9873 7100
rect 9897 7098 9953 7100
rect 9977 7098 10033 7100
rect 10057 7098 10113 7100
rect 9817 7046 9843 7098
rect 9843 7046 9873 7098
rect 9897 7046 9907 7098
rect 9907 7046 9953 7098
rect 9977 7046 10023 7098
rect 10023 7046 10033 7098
rect 10057 7046 10087 7098
rect 10087 7046 10113 7098
rect 9817 7044 9873 7046
rect 9897 7044 9953 7046
rect 9977 7044 10033 7046
rect 10057 7044 10113 7046
rect 10402 7112 10458 7168
rect 10218 6976 10274 7032
rect 10402 6024 10458 6080
rect 9817 6010 9873 6012
rect 9897 6010 9953 6012
rect 9977 6010 10033 6012
rect 10057 6010 10113 6012
rect 9817 5958 9843 6010
rect 9843 5958 9873 6010
rect 9897 5958 9907 6010
rect 9907 5958 9953 6010
rect 9977 5958 10023 6010
rect 10023 5958 10033 6010
rect 10057 5958 10087 6010
rect 10087 5958 10113 6010
rect 9817 5956 9873 5958
rect 9897 5956 9953 5958
rect 9977 5956 10033 5958
rect 10057 5956 10113 5958
rect 10218 5344 10274 5400
rect 9817 4922 9873 4924
rect 9897 4922 9953 4924
rect 9977 4922 10033 4924
rect 10057 4922 10113 4924
rect 9817 4870 9843 4922
rect 9843 4870 9873 4922
rect 9897 4870 9907 4922
rect 9907 4870 9953 4922
rect 9977 4870 10023 4922
rect 10023 4870 10033 4922
rect 10057 4870 10087 4922
rect 10087 4870 10113 4922
rect 9817 4868 9873 4870
rect 9897 4868 9953 4870
rect 9977 4868 10033 4870
rect 10057 4868 10113 4870
rect 9817 3834 9873 3836
rect 9897 3834 9953 3836
rect 9977 3834 10033 3836
rect 10057 3834 10113 3836
rect 9817 3782 9843 3834
rect 9843 3782 9873 3834
rect 9897 3782 9907 3834
rect 9907 3782 9953 3834
rect 9977 3782 10023 3834
rect 10023 3782 10033 3834
rect 10057 3782 10087 3834
rect 10087 3782 10113 3834
rect 9817 3780 9873 3782
rect 9897 3780 9953 3782
rect 9977 3780 10033 3782
rect 10057 3780 10113 3782
rect 10770 8200 10826 8256
rect 11414 12180 11416 12200
rect 11416 12180 11468 12200
rect 11468 12180 11470 12200
rect 11414 12144 11470 12180
rect 11138 11892 11194 11928
rect 11138 11872 11140 11892
rect 11140 11872 11192 11892
rect 11192 11872 11194 11892
rect 10862 7384 10918 7440
rect 10862 6704 10918 6760
rect 10862 6296 10918 6352
rect 8930 1264 8986 1320
rect 9298 2760 9354 2816
rect 9114 1128 9170 1184
rect 9817 2746 9873 2748
rect 9897 2746 9953 2748
rect 9977 2746 10033 2748
rect 10057 2746 10113 2748
rect 9817 2694 9843 2746
rect 9843 2694 9873 2746
rect 9897 2694 9907 2746
rect 9907 2694 9953 2746
rect 9977 2694 10023 2746
rect 10023 2694 10033 2746
rect 10057 2694 10087 2746
rect 10087 2694 10113 2746
rect 9817 2692 9873 2694
rect 9897 2692 9953 2694
rect 9977 2692 10033 2694
rect 10057 2692 10113 2694
rect 9390 2624 9446 2680
rect 10402 2760 10458 2816
rect 14484 25050 14540 25052
rect 14564 25050 14620 25052
rect 14644 25050 14700 25052
rect 14724 25050 14780 25052
rect 14484 24998 14510 25050
rect 14510 24998 14540 25050
rect 14564 24998 14574 25050
rect 14574 24998 14620 25050
rect 14644 24998 14690 25050
rect 14690 24998 14700 25050
rect 14724 24998 14754 25050
rect 14754 24998 14780 25050
rect 14484 24996 14540 24998
rect 14564 24996 14620 24998
rect 14644 24996 14700 24998
rect 14724 24996 14780 24998
rect 14484 23962 14540 23964
rect 14564 23962 14620 23964
rect 14644 23962 14700 23964
rect 14724 23962 14780 23964
rect 14484 23910 14510 23962
rect 14510 23910 14540 23962
rect 14564 23910 14574 23962
rect 14574 23910 14620 23962
rect 14644 23910 14690 23962
rect 14690 23910 14700 23962
rect 14724 23910 14754 23962
rect 14754 23910 14780 23962
rect 14484 23908 14540 23910
rect 14564 23908 14620 23910
rect 14644 23908 14700 23910
rect 14724 23908 14780 23910
rect 14484 22874 14540 22876
rect 14564 22874 14620 22876
rect 14644 22874 14700 22876
rect 14724 22874 14780 22876
rect 14484 22822 14510 22874
rect 14510 22822 14540 22874
rect 14564 22822 14574 22874
rect 14574 22822 14620 22874
rect 14644 22822 14690 22874
rect 14690 22822 14700 22874
rect 14724 22822 14754 22874
rect 14754 22822 14780 22874
rect 14484 22820 14540 22822
rect 14564 22820 14620 22822
rect 14644 22820 14700 22822
rect 14724 22820 14780 22822
rect 14484 21786 14540 21788
rect 14564 21786 14620 21788
rect 14644 21786 14700 21788
rect 14724 21786 14780 21788
rect 14484 21734 14510 21786
rect 14510 21734 14540 21786
rect 14564 21734 14574 21786
rect 14574 21734 14620 21786
rect 14644 21734 14690 21786
rect 14690 21734 14700 21786
rect 14724 21734 14754 21786
rect 14754 21734 14780 21786
rect 14484 21732 14540 21734
rect 14564 21732 14620 21734
rect 14644 21732 14700 21734
rect 14724 21732 14780 21734
rect 14484 20698 14540 20700
rect 14564 20698 14620 20700
rect 14644 20698 14700 20700
rect 14724 20698 14780 20700
rect 14484 20646 14510 20698
rect 14510 20646 14540 20698
rect 14564 20646 14574 20698
rect 14574 20646 14620 20698
rect 14644 20646 14690 20698
rect 14690 20646 14700 20698
rect 14724 20646 14754 20698
rect 14754 20646 14780 20698
rect 14484 20644 14540 20646
rect 14564 20644 14620 20646
rect 14644 20644 14700 20646
rect 14724 20644 14780 20646
rect 14484 19610 14540 19612
rect 14564 19610 14620 19612
rect 14644 19610 14700 19612
rect 14724 19610 14780 19612
rect 14484 19558 14510 19610
rect 14510 19558 14540 19610
rect 14564 19558 14574 19610
rect 14574 19558 14620 19610
rect 14644 19558 14690 19610
rect 14690 19558 14700 19610
rect 14724 19558 14754 19610
rect 14754 19558 14780 19610
rect 14484 19556 14540 19558
rect 14564 19556 14620 19558
rect 14644 19556 14700 19558
rect 14724 19556 14780 19558
rect 13254 19216 13310 19272
rect 12426 16632 12482 16688
rect 11690 12824 11746 12880
rect 11874 12416 11930 12472
rect 12334 12144 12390 12200
rect 13070 15564 13126 15600
rect 13070 15544 13072 15564
rect 13072 15544 13124 15564
rect 13124 15544 13126 15564
rect 13070 12588 13072 12608
rect 13072 12588 13124 12608
rect 13124 12588 13126 12608
rect 13070 12552 13126 12588
rect 12518 12416 12574 12472
rect 14484 18522 14540 18524
rect 14564 18522 14620 18524
rect 14644 18522 14700 18524
rect 14724 18522 14780 18524
rect 14484 18470 14510 18522
rect 14510 18470 14540 18522
rect 14564 18470 14574 18522
rect 14574 18470 14620 18522
rect 14644 18470 14690 18522
rect 14690 18470 14700 18522
rect 14724 18470 14754 18522
rect 14754 18470 14780 18522
rect 14484 18468 14540 18470
rect 14564 18468 14620 18470
rect 14644 18468 14700 18470
rect 14724 18468 14780 18470
rect 14484 17434 14540 17436
rect 14564 17434 14620 17436
rect 14644 17434 14700 17436
rect 14724 17434 14780 17436
rect 14484 17382 14510 17434
rect 14510 17382 14540 17434
rect 14564 17382 14574 17434
rect 14574 17382 14620 17434
rect 14644 17382 14690 17434
rect 14690 17382 14700 17434
rect 14724 17382 14754 17434
rect 14754 17382 14780 17434
rect 14484 17380 14540 17382
rect 14564 17380 14620 17382
rect 14644 17380 14700 17382
rect 14724 17380 14780 17382
rect 16014 18264 16070 18320
rect 17854 17312 17910 17368
rect 14484 16346 14540 16348
rect 14564 16346 14620 16348
rect 14644 16346 14700 16348
rect 14724 16346 14780 16348
rect 14484 16294 14510 16346
rect 14510 16294 14540 16346
rect 14564 16294 14574 16346
rect 14574 16294 14620 16346
rect 14644 16294 14690 16346
rect 14690 16294 14700 16346
rect 14724 16294 14754 16346
rect 14754 16294 14780 16346
rect 14484 16292 14540 16294
rect 14564 16292 14620 16294
rect 14644 16292 14700 16294
rect 14724 16292 14780 16294
rect 12702 8880 12758 8936
rect 12610 8608 12666 8664
rect 12334 8472 12390 8528
rect 12150 7384 12206 7440
rect 11782 6704 11838 6760
rect 12058 6976 12114 7032
rect 12518 7112 12574 7168
rect 12150 4004 12206 4040
rect 12150 3984 12152 4004
rect 12152 3984 12204 4004
rect 12204 3984 12206 4004
rect 11966 3712 12022 3768
rect 13438 12280 13494 12336
rect 13254 11192 13310 11248
rect 13346 10512 13402 10568
rect 14484 15258 14540 15260
rect 14564 15258 14620 15260
rect 14644 15258 14700 15260
rect 14724 15258 14780 15260
rect 14484 15206 14510 15258
rect 14510 15206 14540 15258
rect 14564 15206 14574 15258
rect 14574 15206 14620 15258
rect 14644 15206 14690 15258
rect 14690 15206 14700 15258
rect 14724 15206 14754 15258
rect 14754 15206 14780 15258
rect 14484 15204 14540 15206
rect 14564 15204 14620 15206
rect 14644 15204 14700 15206
rect 14724 15204 14780 15206
rect 14174 14728 14230 14784
rect 13806 13932 13862 13968
rect 13806 13912 13808 13932
rect 13808 13912 13860 13932
rect 13860 13912 13862 13932
rect 13990 12960 14046 13016
rect 13622 12008 13678 12064
rect 13898 11736 13954 11792
rect 13438 9832 13494 9888
rect 13254 9560 13310 9616
rect 13346 8916 13348 8936
rect 13348 8916 13400 8936
rect 13400 8916 13402 8936
rect 13346 8880 13402 8916
rect 14484 14170 14540 14172
rect 14564 14170 14620 14172
rect 14644 14170 14700 14172
rect 14724 14170 14780 14172
rect 14484 14118 14510 14170
rect 14510 14118 14540 14170
rect 14564 14118 14574 14170
rect 14574 14118 14620 14170
rect 14644 14118 14690 14170
rect 14690 14118 14700 14170
rect 14724 14118 14754 14170
rect 14754 14118 14780 14170
rect 14484 14116 14540 14118
rect 14564 14116 14620 14118
rect 14644 14116 14700 14118
rect 14724 14116 14780 14118
rect 16842 16088 16898 16144
rect 14484 13082 14540 13084
rect 14564 13082 14620 13084
rect 14644 13082 14700 13084
rect 14724 13082 14780 13084
rect 14484 13030 14510 13082
rect 14510 13030 14540 13082
rect 14564 13030 14574 13082
rect 14574 13030 14620 13082
rect 14644 13030 14690 13082
rect 14690 13030 14700 13082
rect 14724 13030 14754 13082
rect 14754 13030 14780 13082
rect 14484 13028 14540 13030
rect 14564 13028 14620 13030
rect 14644 13028 14700 13030
rect 14724 13028 14780 13030
rect 14266 12144 14322 12200
rect 14542 12164 14598 12200
rect 14542 12144 14544 12164
rect 14544 12144 14596 12164
rect 14596 12144 14598 12164
rect 14484 11994 14540 11996
rect 14564 11994 14620 11996
rect 14644 11994 14700 11996
rect 14724 11994 14780 11996
rect 14484 11942 14510 11994
rect 14510 11942 14540 11994
rect 14564 11942 14574 11994
rect 14574 11942 14620 11994
rect 14644 11942 14690 11994
rect 14690 11942 14700 11994
rect 14724 11942 14754 11994
rect 14754 11942 14780 11994
rect 14484 11940 14540 11942
rect 14564 11940 14620 11942
rect 14644 11940 14700 11942
rect 14724 11940 14780 11942
rect 13806 10804 13862 10840
rect 13806 10784 13808 10804
rect 13808 10784 13860 10804
rect 13860 10784 13862 10804
rect 15002 11620 15058 11656
rect 15002 11600 15004 11620
rect 15004 11600 15056 11620
rect 15056 11600 15058 11620
rect 14484 10906 14540 10908
rect 14564 10906 14620 10908
rect 14644 10906 14700 10908
rect 14724 10906 14780 10908
rect 14484 10854 14510 10906
rect 14510 10854 14540 10906
rect 14564 10854 14574 10906
rect 14574 10854 14620 10906
rect 14644 10854 14690 10906
rect 14690 10854 14700 10906
rect 14724 10854 14754 10906
rect 14754 10854 14780 10906
rect 14484 10852 14540 10854
rect 14564 10852 14620 10854
rect 14644 10852 14700 10854
rect 14724 10852 14780 10854
rect 14634 10240 14690 10296
rect 13990 10124 14046 10160
rect 13990 10104 13992 10124
rect 13992 10104 14044 10124
rect 14044 10104 14046 10124
rect 14484 9818 14540 9820
rect 14564 9818 14620 9820
rect 14644 9818 14700 9820
rect 14724 9818 14780 9820
rect 14484 9766 14510 9818
rect 14510 9766 14540 9818
rect 14564 9766 14574 9818
rect 14574 9766 14620 9818
rect 14644 9766 14690 9818
rect 14690 9766 14700 9818
rect 14724 9766 14754 9818
rect 14754 9766 14780 9818
rect 14484 9764 14540 9766
rect 14564 9764 14620 9766
rect 14644 9764 14700 9766
rect 14724 9764 14780 9766
rect 14484 8730 14540 8732
rect 14564 8730 14620 8732
rect 14644 8730 14700 8732
rect 14724 8730 14780 8732
rect 14484 8678 14510 8730
rect 14510 8678 14540 8730
rect 14564 8678 14574 8730
rect 14574 8678 14620 8730
rect 14644 8678 14690 8730
rect 14690 8678 14700 8730
rect 14724 8678 14754 8730
rect 14754 8678 14780 8730
rect 14484 8676 14540 8678
rect 14564 8676 14620 8678
rect 14644 8676 14700 8678
rect 14724 8676 14780 8678
rect 13898 8200 13954 8256
rect 13898 7384 13954 7440
rect 13346 6876 13348 6896
rect 13348 6876 13400 6896
rect 13400 6876 13402 6896
rect 13346 6840 13402 6876
rect 13254 6452 13310 6488
rect 13254 6432 13256 6452
rect 13256 6432 13308 6452
rect 13308 6432 13310 6452
rect 14634 8200 14690 8256
rect 16382 13912 16438 13968
rect 15186 12280 15242 12336
rect 15370 10104 15426 10160
rect 15094 8880 15150 8936
rect 14484 7642 14540 7644
rect 14564 7642 14620 7644
rect 14644 7642 14700 7644
rect 14724 7642 14780 7644
rect 14484 7590 14510 7642
rect 14510 7590 14540 7642
rect 14564 7590 14574 7642
rect 14574 7590 14620 7642
rect 14644 7590 14690 7642
rect 14690 7590 14700 7642
rect 14724 7590 14754 7642
rect 14754 7590 14780 7642
rect 14484 7588 14540 7590
rect 14564 7588 14620 7590
rect 14644 7588 14700 7590
rect 14724 7588 14780 7590
rect 14484 6554 14540 6556
rect 14564 6554 14620 6556
rect 14644 6554 14700 6556
rect 14724 6554 14780 6556
rect 14484 6502 14510 6554
rect 14510 6502 14540 6554
rect 14564 6502 14574 6554
rect 14574 6502 14620 6554
rect 14644 6502 14690 6554
rect 14690 6502 14700 6554
rect 14724 6502 14754 6554
rect 14754 6502 14780 6554
rect 14484 6500 14540 6502
rect 14564 6500 14620 6502
rect 14644 6500 14700 6502
rect 14724 6500 14780 6502
rect 12426 4528 12482 4584
rect 14484 5466 14540 5468
rect 14564 5466 14620 5468
rect 14644 5466 14700 5468
rect 14724 5466 14780 5468
rect 14484 5414 14510 5466
rect 14510 5414 14540 5466
rect 14564 5414 14574 5466
rect 14574 5414 14620 5466
rect 14644 5414 14690 5466
rect 14690 5414 14700 5466
rect 14724 5414 14754 5466
rect 14754 5414 14780 5466
rect 14484 5412 14540 5414
rect 14564 5412 14620 5414
rect 14644 5412 14700 5414
rect 14724 5412 14780 5414
rect 14266 4800 14322 4856
rect 13714 4256 13770 4312
rect 13254 3440 13310 3496
rect 13162 3304 13218 3360
rect 12334 3168 12390 3224
rect 12242 2760 12298 2816
rect 11506 2388 11508 2408
rect 11508 2388 11560 2408
rect 11560 2388 11562 2408
rect 11506 2352 11562 2388
rect 11322 2216 11378 2272
rect 13438 3032 13494 3088
rect 12426 2760 12482 2816
rect 15554 9832 15610 9888
rect 16198 10260 16254 10296
rect 16198 10240 16200 10260
rect 16200 10240 16252 10260
rect 16252 10240 16254 10260
rect 16474 13368 16530 13424
rect 16658 12436 16714 12472
rect 16658 12416 16660 12436
rect 16660 12416 16712 12436
rect 16712 12416 16714 12436
rect 18038 15272 18094 15328
rect 17946 14764 17948 14784
rect 17948 14764 18000 14784
rect 18000 14764 18002 14784
rect 17946 14728 18002 14764
rect 17302 12860 17304 12880
rect 17304 12860 17356 12880
rect 17356 12860 17358 12880
rect 17302 12824 17358 12860
rect 17946 12688 18002 12744
rect 18314 12688 18370 12744
rect 17578 12280 17634 12336
rect 17302 12144 17358 12200
rect 16750 11500 16752 11520
rect 16752 11500 16804 11520
rect 16804 11500 16806 11520
rect 16750 11464 16806 11500
rect 17210 10532 17266 10568
rect 17210 10512 17212 10532
rect 17212 10512 17264 10532
rect 17264 10512 17266 10532
rect 17670 11736 17726 11792
rect 16106 6840 16162 6896
rect 17670 9580 17726 9616
rect 17670 9560 17672 9580
rect 17672 9560 17724 9580
rect 17724 9560 17726 9580
rect 16842 9052 16844 9072
rect 16844 9052 16896 9072
rect 16896 9052 16898 9072
rect 16842 9016 16898 9052
rect 18498 12280 18554 12336
rect 19150 25594 19206 25596
rect 19230 25594 19286 25596
rect 19310 25594 19366 25596
rect 19390 25594 19446 25596
rect 19150 25542 19176 25594
rect 19176 25542 19206 25594
rect 19230 25542 19240 25594
rect 19240 25542 19286 25594
rect 19310 25542 19356 25594
rect 19356 25542 19366 25594
rect 19390 25542 19420 25594
rect 19420 25542 19446 25594
rect 19150 25540 19206 25542
rect 19230 25540 19286 25542
rect 19310 25540 19366 25542
rect 19390 25540 19446 25542
rect 19150 24506 19206 24508
rect 19230 24506 19286 24508
rect 19310 24506 19366 24508
rect 19390 24506 19446 24508
rect 19150 24454 19176 24506
rect 19176 24454 19206 24506
rect 19230 24454 19240 24506
rect 19240 24454 19286 24506
rect 19310 24454 19356 24506
rect 19356 24454 19366 24506
rect 19390 24454 19420 24506
rect 19420 24454 19446 24506
rect 19150 24452 19206 24454
rect 19230 24452 19286 24454
rect 19310 24452 19366 24454
rect 19390 24452 19446 24454
rect 20890 23568 20946 23624
rect 19150 23418 19206 23420
rect 19230 23418 19286 23420
rect 19310 23418 19366 23420
rect 19390 23418 19446 23420
rect 19150 23366 19176 23418
rect 19176 23366 19206 23418
rect 19230 23366 19240 23418
rect 19240 23366 19286 23418
rect 19310 23366 19356 23418
rect 19356 23366 19366 23418
rect 19390 23366 19420 23418
rect 19420 23366 19446 23418
rect 19150 23364 19206 23366
rect 19230 23364 19286 23366
rect 19310 23364 19366 23366
rect 19390 23364 19446 23366
rect 19150 22330 19206 22332
rect 19230 22330 19286 22332
rect 19310 22330 19366 22332
rect 19390 22330 19446 22332
rect 19150 22278 19176 22330
rect 19176 22278 19206 22330
rect 19230 22278 19240 22330
rect 19240 22278 19286 22330
rect 19310 22278 19356 22330
rect 19356 22278 19366 22330
rect 19390 22278 19420 22330
rect 19420 22278 19446 22330
rect 19150 22276 19206 22278
rect 19230 22276 19286 22278
rect 19310 22276 19366 22278
rect 19390 22276 19446 22278
rect 19150 21242 19206 21244
rect 19230 21242 19286 21244
rect 19310 21242 19366 21244
rect 19390 21242 19446 21244
rect 19150 21190 19176 21242
rect 19176 21190 19206 21242
rect 19230 21190 19240 21242
rect 19240 21190 19286 21242
rect 19310 21190 19356 21242
rect 19356 21190 19366 21242
rect 19390 21190 19420 21242
rect 19420 21190 19446 21242
rect 19150 21188 19206 21190
rect 19230 21188 19286 21190
rect 19310 21188 19366 21190
rect 19390 21188 19446 21190
rect 19150 20154 19206 20156
rect 19230 20154 19286 20156
rect 19310 20154 19366 20156
rect 19390 20154 19446 20156
rect 19150 20102 19176 20154
rect 19176 20102 19206 20154
rect 19230 20102 19240 20154
rect 19240 20102 19286 20154
rect 19310 20102 19356 20154
rect 19356 20102 19366 20154
rect 19390 20102 19420 20154
rect 19420 20102 19446 20154
rect 19150 20100 19206 20102
rect 19230 20100 19286 20102
rect 19310 20100 19366 20102
rect 19390 20100 19446 20102
rect 19150 19066 19206 19068
rect 19230 19066 19286 19068
rect 19310 19066 19366 19068
rect 19390 19066 19446 19068
rect 19150 19014 19176 19066
rect 19176 19014 19206 19066
rect 19230 19014 19240 19066
rect 19240 19014 19286 19066
rect 19310 19014 19356 19066
rect 19356 19014 19366 19066
rect 19390 19014 19420 19066
rect 19420 19014 19446 19066
rect 19150 19012 19206 19014
rect 19230 19012 19286 19014
rect 19310 19012 19366 19014
rect 19390 19012 19446 19014
rect 19150 17978 19206 17980
rect 19230 17978 19286 17980
rect 19310 17978 19366 17980
rect 19390 17978 19446 17980
rect 19150 17926 19176 17978
rect 19176 17926 19206 17978
rect 19230 17926 19240 17978
rect 19240 17926 19286 17978
rect 19310 17926 19356 17978
rect 19356 17926 19366 17978
rect 19390 17926 19420 17978
rect 19420 17926 19446 17978
rect 19150 17924 19206 17926
rect 19230 17924 19286 17926
rect 19310 17924 19366 17926
rect 19390 17924 19446 17926
rect 19150 16890 19206 16892
rect 19230 16890 19286 16892
rect 19310 16890 19366 16892
rect 19390 16890 19446 16892
rect 19150 16838 19176 16890
rect 19176 16838 19206 16890
rect 19230 16838 19240 16890
rect 19240 16838 19286 16890
rect 19310 16838 19356 16890
rect 19356 16838 19366 16890
rect 19390 16838 19420 16890
rect 19420 16838 19446 16890
rect 19150 16836 19206 16838
rect 19230 16836 19286 16838
rect 19310 16836 19366 16838
rect 19390 16836 19446 16838
rect 19150 15802 19206 15804
rect 19230 15802 19286 15804
rect 19310 15802 19366 15804
rect 19390 15802 19446 15804
rect 19150 15750 19176 15802
rect 19176 15750 19206 15802
rect 19230 15750 19240 15802
rect 19240 15750 19286 15802
rect 19310 15750 19356 15802
rect 19356 15750 19366 15802
rect 19390 15750 19420 15802
rect 19420 15750 19446 15802
rect 19150 15748 19206 15750
rect 19230 15748 19286 15750
rect 19310 15748 19366 15750
rect 19390 15748 19446 15750
rect 18958 15544 19014 15600
rect 19150 14714 19206 14716
rect 19230 14714 19286 14716
rect 19310 14714 19366 14716
rect 19390 14714 19446 14716
rect 19150 14662 19176 14714
rect 19176 14662 19206 14714
rect 19230 14662 19240 14714
rect 19240 14662 19286 14714
rect 19310 14662 19356 14714
rect 19356 14662 19366 14714
rect 19390 14662 19420 14714
rect 19420 14662 19446 14714
rect 19150 14660 19206 14662
rect 19230 14660 19286 14662
rect 19310 14660 19366 14662
rect 19390 14660 19446 14662
rect 19150 13626 19206 13628
rect 19230 13626 19286 13628
rect 19310 13626 19366 13628
rect 19390 13626 19446 13628
rect 19150 13574 19176 13626
rect 19176 13574 19206 13626
rect 19230 13574 19240 13626
rect 19240 13574 19286 13626
rect 19310 13574 19356 13626
rect 19356 13574 19366 13626
rect 19390 13574 19420 13626
rect 19420 13574 19446 13626
rect 19150 13572 19206 13574
rect 19230 13572 19286 13574
rect 19310 13572 19366 13574
rect 19390 13572 19446 13574
rect 19602 13504 19658 13560
rect 18958 12552 19014 12608
rect 19150 12538 19206 12540
rect 19230 12538 19286 12540
rect 19310 12538 19366 12540
rect 19390 12538 19446 12540
rect 19150 12486 19176 12538
rect 19176 12486 19206 12538
rect 19230 12486 19240 12538
rect 19240 12486 19286 12538
rect 19310 12486 19356 12538
rect 19356 12486 19366 12538
rect 19390 12486 19420 12538
rect 19420 12486 19446 12538
rect 19150 12484 19206 12486
rect 19230 12484 19286 12486
rect 19310 12484 19366 12486
rect 19390 12484 19446 12486
rect 20246 15428 20302 15464
rect 20246 15408 20248 15428
rect 20248 15408 20300 15428
rect 20300 15408 20302 15428
rect 20798 20712 20854 20768
rect 20522 20032 20578 20088
rect 18222 11600 18278 11656
rect 18314 10532 18370 10568
rect 18314 10512 18316 10532
rect 18316 10512 18368 10532
rect 18368 10512 18370 10532
rect 20430 12708 20486 12744
rect 20430 12688 20432 12708
rect 20432 12688 20484 12708
rect 20484 12688 20486 12708
rect 20430 12280 20486 12336
rect 18774 11636 18776 11656
rect 18776 11636 18828 11656
rect 18828 11636 18830 11656
rect 18774 11600 18830 11636
rect 19150 11450 19206 11452
rect 19230 11450 19286 11452
rect 19310 11450 19366 11452
rect 19390 11450 19446 11452
rect 19150 11398 19176 11450
rect 19176 11398 19206 11450
rect 19230 11398 19240 11450
rect 19240 11398 19286 11450
rect 19310 11398 19356 11450
rect 19356 11398 19366 11450
rect 19390 11398 19420 11450
rect 19420 11398 19446 11450
rect 19150 11396 19206 11398
rect 19230 11396 19286 11398
rect 19310 11396 19366 11398
rect 19390 11396 19446 11398
rect 20338 11192 20394 11248
rect 17854 9868 17856 9888
rect 17856 9868 17908 9888
rect 17908 9868 17910 9888
rect 17854 9832 17910 9868
rect 17854 8916 17856 8936
rect 17856 8916 17908 8936
rect 17908 8916 17910 8936
rect 17854 8880 17910 8916
rect 16566 7928 16622 7984
rect 16566 7656 16622 7712
rect 16658 6976 16714 7032
rect 15462 5616 15518 5672
rect 14484 4378 14540 4380
rect 14564 4378 14620 4380
rect 14644 4378 14700 4380
rect 14724 4378 14780 4380
rect 14484 4326 14510 4378
rect 14510 4326 14540 4378
rect 14564 4326 14574 4378
rect 14574 4326 14620 4378
rect 14644 4326 14690 4378
rect 14690 4326 14700 4378
rect 14724 4326 14754 4378
rect 14754 4326 14780 4378
rect 14484 4324 14540 4326
rect 14564 4324 14620 4326
rect 14644 4324 14700 4326
rect 14724 4324 14780 4326
rect 13806 3304 13862 3360
rect 14818 3440 14874 3496
rect 14484 3290 14540 3292
rect 14564 3290 14620 3292
rect 14644 3290 14700 3292
rect 14724 3290 14780 3292
rect 14484 3238 14510 3290
rect 14510 3238 14540 3290
rect 14564 3238 14574 3290
rect 14574 3238 14620 3290
rect 14644 3238 14690 3290
rect 14690 3238 14700 3290
rect 14724 3238 14754 3290
rect 14754 3238 14780 3290
rect 14484 3236 14540 3238
rect 14564 3236 14620 3238
rect 14644 3236 14700 3238
rect 14724 3236 14780 3238
rect 14358 2896 14414 2952
rect 16290 6316 16346 6352
rect 16290 6296 16292 6316
rect 16292 6296 16344 6316
rect 16344 6296 16346 6316
rect 16198 5616 16254 5672
rect 17762 8200 17818 8256
rect 17854 7404 17910 7440
rect 17854 7384 17856 7404
rect 17856 7384 17908 7404
rect 17908 7384 17910 7404
rect 18130 7268 18186 7304
rect 18130 7248 18132 7268
rect 18132 7248 18184 7268
rect 18184 7248 18186 7268
rect 18406 7112 18462 7168
rect 17026 5344 17082 5400
rect 16842 4936 16898 4992
rect 16842 4664 16898 4720
rect 16106 4120 16162 4176
rect 15738 3848 15794 3904
rect 17578 3984 17634 4040
rect 15278 3168 15334 3224
rect 16198 3576 16254 3632
rect 16014 3032 16070 3088
rect 14818 2760 14874 2816
rect 14484 2202 14540 2204
rect 14564 2202 14620 2204
rect 14644 2202 14700 2204
rect 14724 2202 14780 2204
rect 14484 2150 14510 2202
rect 14510 2150 14540 2202
rect 14564 2150 14574 2202
rect 14574 2150 14620 2202
rect 14644 2150 14690 2202
rect 14690 2150 14700 2202
rect 14724 2150 14754 2202
rect 14754 2150 14780 2202
rect 14484 2148 14540 2150
rect 14564 2148 14620 2150
rect 14644 2148 14700 2150
rect 14724 2148 14780 2150
rect 13806 1808 13862 1864
rect 13990 1808 14046 1864
rect 15462 1944 15518 2000
rect 20430 11056 20486 11112
rect 19150 10362 19206 10364
rect 19230 10362 19286 10364
rect 19310 10362 19366 10364
rect 19390 10362 19446 10364
rect 19150 10310 19176 10362
rect 19176 10310 19206 10362
rect 19230 10310 19240 10362
rect 19240 10310 19286 10362
rect 19310 10310 19356 10362
rect 19356 10310 19366 10362
rect 19390 10310 19420 10362
rect 19420 10310 19446 10362
rect 19150 10308 19206 10310
rect 19230 10308 19286 10310
rect 19310 10308 19366 10310
rect 19390 10308 19446 10310
rect 19602 10376 19658 10432
rect 19150 9274 19206 9276
rect 19230 9274 19286 9276
rect 19310 9274 19366 9276
rect 19390 9274 19446 9276
rect 19150 9222 19176 9274
rect 19176 9222 19206 9274
rect 19230 9222 19240 9274
rect 19240 9222 19286 9274
rect 19310 9222 19356 9274
rect 19356 9222 19366 9274
rect 19390 9222 19420 9274
rect 19420 9222 19446 9274
rect 19150 9220 19206 9222
rect 19230 9220 19286 9222
rect 19310 9220 19366 9222
rect 19390 9220 19446 9222
rect 19050 8744 19106 8800
rect 19150 8186 19206 8188
rect 19230 8186 19286 8188
rect 19310 8186 19366 8188
rect 19390 8186 19446 8188
rect 19150 8134 19176 8186
rect 19176 8134 19206 8186
rect 19230 8134 19240 8186
rect 19240 8134 19286 8186
rect 19310 8134 19356 8186
rect 19356 8134 19366 8186
rect 19390 8134 19420 8186
rect 19420 8134 19446 8186
rect 19150 8132 19206 8134
rect 19230 8132 19286 8134
rect 19310 8132 19366 8134
rect 19390 8132 19446 8134
rect 19150 7098 19206 7100
rect 19230 7098 19286 7100
rect 19310 7098 19366 7100
rect 19390 7098 19446 7100
rect 19150 7046 19176 7098
rect 19176 7046 19206 7098
rect 19230 7046 19240 7098
rect 19240 7046 19286 7098
rect 19310 7046 19356 7098
rect 19356 7046 19366 7098
rect 19390 7046 19420 7098
rect 19420 7046 19446 7098
rect 19150 7044 19206 7046
rect 19230 7044 19286 7046
rect 19310 7044 19366 7046
rect 19390 7044 19446 7046
rect 18958 6024 19014 6080
rect 19150 6010 19206 6012
rect 19230 6010 19286 6012
rect 19310 6010 19366 6012
rect 19390 6010 19446 6012
rect 19150 5958 19176 6010
rect 19176 5958 19206 6010
rect 19230 5958 19240 6010
rect 19240 5958 19286 6010
rect 19310 5958 19356 6010
rect 19356 5958 19366 6010
rect 19390 5958 19420 6010
rect 19420 5958 19446 6010
rect 19150 5956 19206 5958
rect 19230 5956 19286 5958
rect 19310 5956 19366 5958
rect 19390 5956 19446 5958
rect 18958 5616 19014 5672
rect 19150 4922 19206 4924
rect 19230 4922 19286 4924
rect 19310 4922 19366 4924
rect 19390 4922 19446 4924
rect 19150 4870 19176 4922
rect 19176 4870 19206 4922
rect 19230 4870 19240 4922
rect 19240 4870 19286 4922
rect 19310 4870 19356 4922
rect 19356 4870 19366 4922
rect 19390 4870 19420 4922
rect 19420 4870 19446 4922
rect 19150 4868 19206 4870
rect 19230 4868 19286 4870
rect 19310 4868 19366 4870
rect 19390 4868 19446 4870
rect 17670 3052 17726 3088
rect 17670 3032 17672 3052
rect 17672 3032 17724 3052
rect 17724 3032 17726 3052
rect 17486 2488 17542 2544
rect 16658 1672 16714 1728
rect 18498 1536 18554 1592
rect 17578 1400 17634 1456
rect 18682 2896 18738 2952
rect 20430 8608 20486 8664
rect 19150 3834 19206 3836
rect 19230 3834 19286 3836
rect 19310 3834 19366 3836
rect 19390 3834 19446 3836
rect 19150 3782 19176 3834
rect 19176 3782 19206 3834
rect 19230 3782 19240 3834
rect 19240 3782 19286 3834
rect 19310 3782 19356 3834
rect 19356 3782 19366 3834
rect 19390 3782 19420 3834
rect 19420 3782 19446 3834
rect 19150 3780 19206 3782
rect 19230 3780 19286 3782
rect 19310 3780 19366 3782
rect 19390 3780 19446 3782
rect 19150 2746 19206 2748
rect 19230 2746 19286 2748
rect 19310 2746 19366 2748
rect 19390 2746 19446 2748
rect 19150 2694 19176 2746
rect 19176 2694 19206 2746
rect 19230 2694 19240 2746
rect 19240 2694 19286 2746
rect 19310 2694 19356 2746
rect 19356 2694 19366 2746
rect 19390 2694 19420 2746
rect 19420 2694 19446 2746
rect 19150 2692 19206 2694
rect 19230 2692 19286 2694
rect 19310 2692 19366 2694
rect 19390 2692 19446 2694
rect 21534 23432 21590 23488
rect 20982 19352 21038 19408
rect 22914 27376 22970 27432
rect 24294 26288 24350 26344
rect 23817 25050 23873 25052
rect 23897 25050 23953 25052
rect 23977 25050 24033 25052
rect 24057 25050 24113 25052
rect 23817 24998 23843 25050
rect 23843 24998 23873 25050
rect 23897 24998 23907 25050
rect 23907 24998 23953 25050
rect 23977 24998 24023 25050
rect 24023 24998 24033 25050
rect 24057 24998 24087 25050
rect 24087 24998 24113 25050
rect 23817 24996 23873 24998
rect 23897 24996 23953 24998
rect 23977 24996 24033 24998
rect 24057 24996 24113 24998
rect 23190 24248 23246 24304
rect 23006 23468 23008 23488
rect 23008 23468 23060 23488
rect 23060 23468 23062 23488
rect 23006 23432 23062 23468
rect 21994 13504 22050 13560
rect 20614 10668 20670 10704
rect 20614 10648 20616 10668
rect 20616 10648 20668 10668
rect 20668 10648 20670 10668
rect 21442 12724 21444 12744
rect 21444 12724 21496 12744
rect 21496 12724 21498 12744
rect 21442 12688 21498 12724
rect 22270 15680 22326 15736
rect 22270 13368 22326 13424
rect 20890 8780 20892 8800
rect 20892 8780 20944 8800
rect 20944 8780 20946 8800
rect 20890 8744 20946 8780
rect 20614 7248 20670 7304
rect 21626 7928 21682 7984
rect 23817 23962 23873 23964
rect 23897 23962 23953 23964
rect 23977 23962 24033 23964
rect 24057 23962 24113 23964
rect 23817 23910 23843 23962
rect 23843 23910 23873 23962
rect 23897 23910 23907 23962
rect 23907 23910 23953 23962
rect 23977 23910 24023 23962
rect 24023 23910 24033 23962
rect 24057 23910 24087 23962
rect 24087 23910 24113 23962
rect 23817 23908 23873 23910
rect 23897 23908 23953 23910
rect 23977 23908 24033 23910
rect 24057 23908 24113 23910
rect 24938 25336 24994 25392
rect 24294 23160 24350 23216
rect 23817 22874 23873 22876
rect 23897 22874 23953 22876
rect 23977 22874 24033 22876
rect 24057 22874 24113 22876
rect 23817 22822 23843 22874
rect 23843 22822 23873 22874
rect 23897 22822 23907 22874
rect 23907 22822 23953 22874
rect 23977 22822 24023 22874
rect 24023 22822 24033 22874
rect 24057 22822 24087 22874
rect 24087 22822 24113 22874
rect 23817 22820 23873 22822
rect 23897 22820 23953 22822
rect 23977 22820 24033 22822
rect 24057 22820 24113 22822
rect 24202 22208 24258 22264
rect 23817 21786 23873 21788
rect 23897 21786 23953 21788
rect 23977 21786 24033 21788
rect 24057 21786 24113 21788
rect 23817 21734 23843 21786
rect 23843 21734 23873 21786
rect 23897 21734 23907 21786
rect 23907 21734 23953 21786
rect 23977 21734 24023 21786
rect 24023 21734 24033 21786
rect 24057 21734 24087 21786
rect 24087 21734 24113 21786
rect 23817 21732 23873 21734
rect 23897 21732 23953 21734
rect 23977 21732 24033 21734
rect 24057 21732 24113 21734
rect 23190 20712 23246 20768
rect 23006 19352 23062 19408
rect 23006 19236 23062 19272
rect 23006 19216 23008 19236
rect 23008 19216 23060 19236
rect 23060 19216 23062 19236
rect 23006 18692 23062 18728
rect 23006 18672 23008 18692
rect 23008 18672 23060 18692
rect 23060 18672 23062 18692
rect 23098 18264 23154 18320
rect 22638 18028 22640 18048
rect 22640 18028 22692 18048
rect 22692 18028 22694 18048
rect 22638 17992 22694 18028
rect 22638 12280 22694 12336
rect 23817 20698 23873 20700
rect 23897 20698 23953 20700
rect 23977 20698 24033 20700
rect 24057 20698 24113 20700
rect 23817 20646 23843 20698
rect 23843 20646 23873 20698
rect 23897 20646 23907 20698
rect 23907 20646 23953 20698
rect 23977 20646 24023 20698
rect 24023 20646 24033 20698
rect 24057 20646 24087 20698
rect 24087 20646 24113 20698
rect 23817 20644 23873 20646
rect 23897 20644 23953 20646
rect 23977 20644 24033 20646
rect 24057 20644 24113 20646
rect 23817 19610 23873 19612
rect 23897 19610 23953 19612
rect 23977 19610 24033 19612
rect 24057 19610 24113 19612
rect 23817 19558 23843 19610
rect 23843 19558 23873 19610
rect 23897 19558 23907 19610
rect 23907 19558 23953 19610
rect 23977 19558 24023 19610
rect 24023 19558 24033 19610
rect 24057 19558 24087 19610
rect 24087 19558 24113 19610
rect 23817 19556 23873 19558
rect 23897 19556 23953 19558
rect 23977 19556 24033 19558
rect 24057 19556 24113 19558
rect 24202 19080 24258 19136
rect 23817 18522 23873 18524
rect 23897 18522 23953 18524
rect 23977 18522 24033 18524
rect 24057 18522 24113 18524
rect 23817 18470 23843 18522
rect 23843 18470 23873 18522
rect 23897 18470 23907 18522
rect 23907 18470 23953 18522
rect 23977 18470 24023 18522
rect 24023 18470 24033 18522
rect 24057 18470 24087 18522
rect 24087 18470 24113 18522
rect 23817 18468 23873 18470
rect 23897 18468 23953 18470
rect 23977 18468 24033 18470
rect 24057 18468 24113 18470
rect 23558 18128 23614 18184
rect 23466 17312 23522 17368
rect 23006 15272 23062 15328
rect 23282 15988 23284 16008
rect 23284 15988 23336 16008
rect 23336 15988 23338 16008
rect 23282 15952 23338 15988
rect 22914 14356 22916 14376
rect 22916 14356 22968 14376
rect 22968 14356 22970 14376
rect 22914 14320 22970 14356
rect 22822 12552 22878 12608
rect 22822 12416 22878 12472
rect 23282 12552 23338 12608
rect 22546 10532 22602 10568
rect 22546 10512 22548 10532
rect 22548 10512 22600 10532
rect 22600 10512 22602 10532
rect 22454 9968 22510 10024
rect 23817 17434 23873 17436
rect 23897 17434 23953 17436
rect 23977 17434 24033 17436
rect 24057 17434 24113 17436
rect 23817 17382 23843 17434
rect 23843 17382 23873 17434
rect 23897 17382 23907 17434
rect 23907 17382 23953 17434
rect 23977 17382 24023 17434
rect 24023 17382 24033 17434
rect 24057 17382 24087 17434
rect 24087 17382 24113 17434
rect 23817 17380 23873 17382
rect 23897 17380 23953 17382
rect 23977 17380 24033 17382
rect 24057 17380 24113 17382
rect 24386 17060 24442 17096
rect 24386 17040 24388 17060
rect 24388 17040 24440 17060
rect 24440 17040 24442 17060
rect 23650 15952 23706 16008
rect 23817 16346 23873 16348
rect 23897 16346 23953 16348
rect 23977 16346 24033 16348
rect 24057 16346 24113 16348
rect 23817 16294 23843 16346
rect 23843 16294 23873 16346
rect 23897 16294 23907 16346
rect 23907 16294 23953 16346
rect 23977 16294 24023 16346
rect 24023 16294 24033 16346
rect 24057 16294 24087 16346
rect 24087 16294 24113 16346
rect 23817 16292 23873 16294
rect 23897 16292 23953 16294
rect 23977 16292 24033 16294
rect 24057 16292 24113 16294
rect 23466 13368 23522 13424
rect 23817 15258 23873 15260
rect 23897 15258 23953 15260
rect 23977 15258 24033 15260
rect 24057 15258 24113 15260
rect 23817 15206 23843 15258
rect 23843 15206 23873 15258
rect 23897 15206 23907 15258
rect 23907 15206 23953 15258
rect 23977 15206 24023 15258
rect 24023 15206 24033 15258
rect 24057 15206 24087 15258
rect 24087 15206 24113 15258
rect 23817 15204 23873 15206
rect 23897 15204 23953 15206
rect 23977 15204 24033 15206
rect 24057 15204 24113 15206
rect 23817 14170 23873 14172
rect 23897 14170 23953 14172
rect 23977 14170 24033 14172
rect 24057 14170 24113 14172
rect 23817 14118 23843 14170
rect 23843 14118 23873 14170
rect 23897 14118 23907 14170
rect 23907 14118 23953 14170
rect 23977 14118 24023 14170
rect 24023 14118 24033 14170
rect 24057 14118 24087 14170
rect 24087 14118 24113 14170
rect 23817 14116 23873 14118
rect 23897 14116 23953 14118
rect 23977 14116 24033 14118
rect 24057 14116 24113 14118
rect 24386 16668 24388 16688
rect 24388 16668 24440 16688
rect 24440 16668 24442 16688
rect 24386 16632 24442 16668
rect 24294 14864 24350 14920
rect 24018 13504 24074 13560
rect 24478 13504 24534 13560
rect 24294 13368 24350 13424
rect 23558 12552 23614 12608
rect 23817 13082 23873 13084
rect 23897 13082 23953 13084
rect 23977 13082 24033 13084
rect 24057 13082 24113 13084
rect 23817 13030 23843 13082
rect 23843 13030 23873 13082
rect 23897 13030 23907 13082
rect 23907 13030 23953 13082
rect 23977 13030 24023 13082
rect 24023 13030 24033 13082
rect 24057 13030 24087 13082
rect 24087 13030 24113 13082
rect 23817 13028 23873 13030
rect 23897 13028 23953 13030
rect 23977 13028 24033 13030
rect 24057 13028 24113 13030
rect 24754 15680 24810 15736
rect 25766 23568 25822 23624
rect 25030 21120 25086 21176
rect 25122 18164 25124 18184
rect 25124 18164 25176 18184
rect 25176 18164 25178 18184
rect 25122 18128 25178 18164
rect 25030 17040 25086 17096
rect 24846 14320 24902 14376
rect 24662 12824 24718 12880
rect 23374 12144 23430 12200
rect 24478 12688 24534 12744
rect 23817 11994 23873 11996
rect 23897 11994 23953 11996
rect 23977 11994 24033 11996
rect 24057 11994 24113 11996
rect 23817 11942 23843 11994
rect 23843 11942 23873 11994
rect 23897 11942 23907 11994
rect 23907 11942 23953 11994
rect 23977 11942 24023 11994
rect 24023 11942 24033 11994
rect 24057 11942 24087 11994
rect 24087 11942 24113 11994
rect 23817 11940 23873 11942
rect 23897 11940 23953 11942
rect 23977 11940 24033 11942
rect 24057 11940 24113 11942
rect 23650 11756 23706 11792
rect 23650 11736 23652 11756
rect 23652 11736 23704 11756
rect 23704 11736 23706 11756
rect 21350 7692 21352 7712
rect 21352 7692 21404 7712
rect 21404 7692 21406 7712
rect 21350 7656 21406 7692
rect 21258 7384 21314 7440
rect 20706 5772 20762 5808
rect 20706 5752 20708 5772
rect 20708 5752 20760 5772
rect 20760 5752 20762 5772
rect 20614 5616 20670 5672
rect 21350 4820 21406 4856
rect 21350 4800 21352 4820
rect 21352 4800 21404 4820
rect 21404 4800 21406 4820
rect 21626 7792 21682 7848
rect 23190 8608 23246 8664
rect 23282 8356 23338 8392
rect 23282 8336 23284 8356
rect 23284 8336 23336 8356
rect 23336 8336 23338 8356
rect 22270 5888 22326 5944
rect 23098 6840 23154 6896
rect 23190 5788 23192 5808
rect 23192 5788 23244 5808
rect 23244 5788 23246 5808
rect 23190 5752 23246 5788
rect 21902 5072 21958 5128
rect 21534 4256 21590 4312
rect 19602 1400 19658 1456
rect 19418 992 19474 1048
rect 20706 1808 20762 1864
rect 20062 856 20118 912
rect 22178 5072 22234 5128
rect 23190 5344 23246 5400
rect 23190 5072 23246 5128
rect 22086 4528 22142 4584
rect 23006 4392 23062 4448
rect 22730 4120 22786 4176
rect 22362 3576 22418 3632
rect 22270 2352 22326 2408
rect 22454 1400 22510 1456
rect 23817 10906 23873 10908
rect 23897 10906 23953 10908
rect 23977 10906 24033 10908
rect 24057 10906 24113 10908
rect 23817 10854 23843 10906
rect 23843 10854 23873 10906
rect 23897 10854 23907 10906
rect 23907 10854 23953 10906
rect 23977 10854 24023 10906
rect 24023 10854 24033 10906
rect 24057 10854 24087 10906
rect 24087 10854 24113 10906
rect 23817 10852 23873 10854
rect 23897 10852 23953 10854
rect 23977 10852 24033 10854
rect 24057 10852 24113 10854
rect 24202 10784 24258 10840
rect 23817 9818 23873 9820
rect 23897 9818 23953 9820
rect 23977 9818 24033 9820
rect 24057 9818 24113 9820
rect 23817 9766 23843 9818
rect 23843 9766 23873 9818
rect 23897 9766 23907 9818
rect 23907 9766 23953 9818
rect 23977 9766 24023 9818
rect 24023 9766 24033 9818
rect 24057 9766 24087 9818
rect 24087 9766 24113 9818
rect 23817 9764 23873 9766
rect 23897 9764 23953 9766
rect 23977 9764 24033 9766
rect 24057 9764 24113 9766
rect 23926 9444 23982 9480
rect 23926 9424 23928 9444
rect 23928 9424 23980 9444
rect 23980 9424 23982 9444
rect 24386 10684 24388 10704
rect 24388 10684 24440 10704
rect 24440 10684 24442 10704
rect 24386 10648 24442 10684
rect 23742 8880 23798 8936
rect 23817 8730 23873 8732
rect 23897 8730 23953 8732
rect 23977 8730 24033 8732
rect 24057 8730 24113 8732
rect 23817 8678 23843 8730
rect 23843 8678 23873 8730
rect 23897 8678 23907 8730
rect 23907 8678 23953 8730
rect 23977 8678 24023 8730
rect 24023 8678 24033 8730
rect 24057 8678 24087 8730
rect 24087 8678 24113 8730
rect 23817 8676 23873 8678
rect 23897 8676 23953 8678
rect 23977 8676 24033 8678
rect 24057 8676 24113 8678
rect 23817 7642 23873 7644
rect 23897 7642 23953 7644
rect 23977 7642 24033 7644
rect 24057 7642 24113 7644
rect 23817 7590 23843 7642
rect 23843 7590 23873 7642
rect 23897 7590 23907 7642
rect 23907 7590 23953 7642
rect 23977 7590 24023 7642
rect 24023 7590 24033 7642
rect 24057 7590 24087 7642
rect 24087 7590 24113 7642
rect 23817 7588 23873 7590
rect 23897 7588 23953 7590
rect 23977 7588 24033 7590
rect 24057 7588 24113 7590
rect 23742 7384 23798 7440
rect 23558 6740 23560 6760
rect 23560 6740 23612 6760
rect 23612 6740 23614 6760
rect 23558 6704 23614 6740
rect 23817 6554 23873 6556
rect 23897 6554 23953 6556
rect 23977 6554 24033 6556
rect 24057 6554 24113 6556
rect 23817 6502 23843 6554
rect 23843 6502 23873 6554
rect 23897 6502 23907 6554
rect 23907 6502 23953 6554
rect 23977 6502 24023 6554
rect 24023 6502 24033 6554
rect 24057 6502 24087 6554
rect 24087 6502 24113 6554
rect 23817 6500 23873 6502
rect 23897 6500 23953 6502
rect 23977 6500 24033 6502
rect 24057 6500 24113 6502
rect 23650 4800 23706 4856
rect 23650 4700 23652 4720
rect 23652 4700 23704 4720
rect 23704 4700 23706 4720
rect 23650 4664 23706 4700
rect 23558 4256 23614 4312
rect 23282 3984 23338 4040
rect 23098 3168 23154 3224
rect 23006 2916 23062 2952
rect 23006 2896 23008 2916
rect 23008 2896 23060 2916
rect 23060 2896 23062 2916
rect 23098 2488 23154 2544
rect 23558 1400 23614 1456
rect 23374 1264 23430 1320
rect 23190 1128 23246 1184
rect 23817 5466 23873 5468
rect 23897 5466 23953 5468
rect 23977 5466 24033 5468
rect 24057 5466 24113 5468
rect 23817 5414 23843 5466
rect 23843 5414 23873 5466
rect 23897 5414 23907 5466
rect 23907 5414 23953 5466
rect 23977 5414 24023 5466
rect 24023 5414 24033 5466
rect 24057 5414 24087 5466
rect 24087 5414 24113 5466
rect 23817 5412 23873 5414
rect 23897 5412 23953 5414
rect 23977 5412 24033 5414
rect 24057 5412 24113 5414
rect 23817 4378 23873 4380
rect 23897 4378 23953 4380
rect 23977 4378 24033 4380
rect 24057 4378 24113 4380
rect 23817 4326 23843 4378
rect 23843 4326 23873 4378
rect 23897 4326 23907 4378
rect 23907 4326 23953 4378
rect 23977 4326 24023 4378
rect 24023 4326 24033 4378
rect 24057 4326 24087 4378
rect 24087 4326 24113 4378
rect 23817 4324 23873 4326
rect 23897 4324 23953 4326
rect 23977 4324 24033 4326
rect 24057 4324 24113 4326
rect 23817 3290 23873 3292
rect 23897 3290 23953 3292
rect 23977 3290 24033 3292
rect 24057 3290 24113 3292
rect 23817 3238 23843 3290
rect 23843 3238 23873 3290
rect 23897 3238 23907 3290
rect 23907 3238 23953 3290
rect 23977 3238 24023 3290
rect 24023 3238 24033 3290
rect 24057 3238 24087 3290
rect 24087 3238 24113 3290
rect 23817 3236 23873 3238
rect 23897 3236 23953 3238
rect 23977 3236 24033 3238
rect 24057 3236 24113 3238
rect 24846 11636 24848 11656
rect 24848 11636 24900 11656
rect 24900 11636 24902 11656
rect 24846 11600 24902 11636
rect 24938 10376 24994 10432
rect 24938 9696 24994 9752
rect 24846 9460 24848 9480
rect 24848 9460 24900 9480
rect 24900 9460 24902 9480
rect 24846 9424 24902 9460
rect 25214 9016 25270 9072
rect 24754 8472 24810 8528
rect 24754 7284 24756 7304
rect 24756 7284 24808 7304
rect 24808 7284 24810 7304
rect 24754 7248 24810 7284
rect 24294 6568 24350 6624
rect 24570 6452 24626 6488
rect 24570 6432 24572 6452
rect 24572 6432 24624 6452
rect 24624 6432 24626 6452
rect 24754 6196 24756 6216
rect 24756 6196 24808 6216
rect 24808 6196 24810 6216
rect 24754 6160 24810 6196
rect 24938 5616 24994 5672
rect 25030 5208 25086 5264
rect 24846 5072 24902 5128
rect 24754 3440 24810 3496
rect 23817 2202 23873 2204
rect 23897 2202 23953 2204
rect 23977 2202 24033 2204
rect 24057 2202 24113 2204
rect 23817 2150 23843 2202
rect 23843 2150 23873 2202
rect 23897 2150 23907 2202
rect 23907 2150 23953 2202
rect 23977 2150 24023 2202
rect 24023 2150 24033 2202
rect 24057 2150 24087 2202
rect 24087 2150 24113 2202
rect 23817 2148 23873 2150
rect 23897 2148 23953 2150
rect 23977 2148 24033 2150
rect 24057 2148 24113 2150
rect 24938 4528 24994 4584
rect 24938 3440 24994 3496
rect 25398 13912 25454 13968
rect 25490 11736 25546 11792
rect 25306 7656 25362 7712
rect 25214 4120 25270 4176
rect 25122 448 25178 504
rect 26870 1672 26926 1728
<< metal3 >>
rect 22909 27434 22975 27437
rect 27048 27434 27528 27464
rect 22909 27432 27528 27434
rect 22909 27376 22914 27432
rect 22970 27376 27528 27432
rect 22909 27374 27528 27376
rect 22909 27371 22975 27374
rect 27048 27344 27528 27374
rect 24289 26346 24355 26349
rect 27048 26346 27528 26376
rect 24289 26344 27528 26346
rect 24289 26288 24294 26344
rect 24350 26288 27528 26344
rect 24289 26286 27528 26288
rect 24289 26283 24355 26286
rect 27048 26256 27528 26286
rect 9805 25600 10125 25601
rect 9805 25536 9813 25600
rect 9877 25536 9893 25600
rect 9957 25536 9973 25600
rect 10037 25536 10053 25600
rect 10117 25536 10125 25600
rect 9805 25535 10125 25536
rect 19138 25600 19458 25601
rect 19138 25536 19146 25600
rect 19210 25536 19226 25600
rect 19290 25536 19306 25600
rect 19370 25536 19386 25600
rect 19450 25536 19458 25600
rect 19138 25535 19458 25536
rect 24933 25394 24999 25397
rect 27048 25394 27528 25424
rect 24933 25392 27528 25394
rect 24933 25336 24938 25392
rect 24994 25336 27528 25392
rect 24933 25334 27528 25336
rect 24933 25331 24999 25334
rect 27048 25304 27528 25334
rect 5138 25056 5458 25057
rect 5138 24992 5146 25056
rect 5210 24992 5226 25056
rect 5290 24992 5306 25056
rect 5370 24992 5386 25056
rect 5450 24992 5458 25056
rect 5138 24991 5458 24992
rect 14472 25056 14792 25057
rect 14472 24992 14480 25056
rect 14544 24992 14560 25056
rect 14624 24992 14640 25056
rect 14704 24992 14720 25056
rect 14784 24992 14792 25056
rect 14472 24991 14792 24992
rect 23805 25056 24125 25057
rect 23805 24992 23813 25056
rect 23877 24992 23893 25056
rect 23957 24992 23973 25056
rect 24037 24992 24053 25056
rect 24117 24992 24125 25056
rect 23805 24991 24125 24992
rect 9805 24512 10125 24513
rect 9805 24448 9813 24512
rect 9877 24448 9893 24512
rect 9957 24448 9973 24512
rect 10037 24448 10053 24512
rect 10117 24448 10125 24512
rect 9805 24447 10125 24448
rect 19138 24512 19458 24513
rect 19138 24448 19146 24512
rect 19210 24448 19226 24512
rect 19290 24448 19306 24512
rect 19370 24448 19386 24512
rect 19450 24448 19458 24512
rect 19138 24447 19458 24448
rect 23185 24306 23251 24309
rect 27048 24306 27528 24336
rect 23185 24304 27528 24306
rect 23185 24248 23190 24304
rect 23246 24248 27528 24304
rect 23185 24246 27528 24248
rect 23185 24243 23251 24246
rect 27048 24216 27528 24246
rect 5138 23968 5458 23969
rect 5138 23904 5146 23968
rect 5210 23904 5226 23968
rect 5290 23904 5306 23968
rect 5370 23904 5386 23968
rect 5450 23904 5458 23968
rect 5138 23903 5458 23904
rect 14472 23968 14792 23969
rect 14472 23904 14480 23968
rect 14544 23904 14560 23968
rect 14624 23904 14640 23968
rect 14704 23904 14720 23968
rect 14784 23904 14792 23968
rect 14472 23903 14792 23904
rect 23805 23968 24125 23969
rect 23805 23904 23813 23968
rect 23877 23904 23893 23968
rect 23957 23904 23973 23968
rect 24037 23904 24053 23968
rect 24117 23904 24125 23968
rect 23805 23903 24125 23904
rect 20885 23626 20951 23629
rect 25761 23626 25827 23629
rect 20885 23624 25827 23626
rect 20885 23568 20890 23624
rect 20946 23568 25766 23624
rect 25822 23568 25827 23624
rect 20885 23566 25827 23568
rect 20885 23563 20951 23566
rect 25761 23563 25827 23566
rect 21529 23490 21595 23493
rect 23001 23490 23067 23493
rect 21529 23488 23067 23490
rect 21529 23432 21534 23488
rect 21590 23432 23006 23488
rect 23062 23432 23067 23488
rect 21529 23430 23067 23432
rect 21529 23427 21595 23430
rect 23001 23427 23067 23430
rect 9805 23424 10125 23425
rect 9805 23360 9813 23424
rect 9877 23360 9893 23424
rect 9957 23360 9973 23424
rect 10037 23360 10053 23424
rect 10117 23360 10125 23424
rect 9805 23359 10125 23360
rect 19138 23424 19458 23425
rect 19138 23360 19146 23424
rect 19210 23360 19226 23424
rect 19290 23360 19306 23424
rect 19370 23360 19386 23424
rect 19450 23360 19458 23424
rect 19138 23359 19458 23360
rect 24289 23218 24355 23221
rect 27048 23218 27528 23248
rect 24289 23216 27528 23218
rect 24289 23160 24294 23216
rect 24350 23160 27528 23216
rect 24289 23158 27528 23160
rect 24289 23155 24355 23158
rect 27048 23128 27528 23158
rect 5138 22880 5458 22881
rect 5138 22816 5146 22880
rect 5210 22816 5226 22880
rect 5290 22816 5306 22880
rect 5370 22816 5386 22880
rect 5450 22816 5458 22880
rect 5138 22815 5458 22816
rect 14472 22880 14792 22881
rect 14472 22816 14480 22880
rect 14544 22816 14560 22880
rect 14624 22816 14640 22880
rect 14704 22816 14720 22880
rect 14784 22816 14792 22880
rect 14472 22815 14792 22816
rect 23805 22880 24125 22881
rect 23805 22816 23813 22880
rect 23877 22816 23893 22880
rect 23957 22816 23973 22880
rect 24037 22816 24053 22880
rect 24117 22816 24125 22880
rect 23805 22815 24125 22816
rect 9805 22336 10125 22337
rect 9805 22272 9813 22336
rect 9877 22272 9893 22336
rect 9957 22272 9973 22336
rect 10037 22272 10053 22336
rect 10117 22272 10125 22336
rect 9805 22271 10125 22272
rect 19138 22336 19458 22337
rect 19138 22272 19146 22336
rect 19210 22272 19226 22336
rect 19290 22272 19306 22336
rect 19370 22272 19386 22336
rect 19450 22272 19458 22336
rect 19138 22271 19458 22272
rect 24197 22266 24263 22269
rect 27048 22266 27528 22296
rect 24197 22264 27528 22266
rect 24197 22208 24202 22264
rect 24258 22208 27528 22264
rect 24197 22206 27528 22208
rect 24197 22203 24263 22206
rect 27048 22176 27528 22206
rect 5138 21792 5458 21793
rect 5138 21728 5146 21792
rect 5210 21728 5226 21792
rect 5290 21728 5306 21792
rect 5370 21728 5386 21792
rect 5450 21728 5458 21792
rect 5138 21727 5458 21728
rect 14472 21792 14792 21793
rect 14472 21728 14480 21792
rect 14544 21728 14560 21792
rect 14624 21728 14640 21792
rect 14704 21728 14720 21792
rect 14784 21728 14792 21792
rect 14472 21727 14792 21728
rect 23805 21792 24125 21793
rect 23805 21728 23813 21792
rect 23877 21728 23893 21792
rect 23957 21728 23973 21792
rect 24037 21728 24053 21792
rect 24117 21728 24125 21792
rect 23805 21727 24125 21728
rect 9805 21248 10125 21249
rect 9805 21184 9813 21248
rect 9877 21184 9893 21248
rect 9957 21184 9973 21248
rect 10037 21184 10053 21248
rect 10117 21184 10125 21248
rect 9805 21183 10125 21184
rect 19138 21248 19458 21249
rect 19138 21184 19146 21248
rect 19210 21184 19226 21248
rect 19290 21184 19306 21248
rect 19370 21184 19386 21248
rect 19450 21184 19458 21248
rect 19138 21183 19458 21184
rect 25025 21178 25091 21181
rect 27048 21178 27528 21208
rect 25025 21176 27528 21178
rect 25025 21120 25030 21176
rect 25086 21120 27528 21176
rect 25025 21118 27528 21120
rect 25025 21115 25091 21118
rect 27048 21088 27528 21118
rect 20793 20770 20859 20773
rect 23185 20770 23251 20773
rect 20793 20768 23251 20770
rect 20793 20712 20798 20768
rect 20854 20712 23190 20768
rect 23246 20712 23251 20768
rect 20793 20710 23251 20712
rect 20793 20707 20859 20710
rect 23185 20707 23251 20710
rect 5138 20704 5458 20705
rect 5138 20640 5146 20704
rect 5210 20640 5226 20704
rect 5290 20640 5306 20704
rect 5370 20640 5386 20704
rect 5450 20640 5458 20704
rect 5138 20639 5458 20640
rect 14472 20704 14792 20705
rect 14472 20640 14480 20704
rect 14544 20640 14560 20704
rect 14624 20640 14640 20704
rect 14704 20640 14720 20704
rect 14784 20640 14792 20704
rect 14472 20639 14792 20640
rect 23805 20704 24125 20705
rect 23805 20640 23813 20704
rect 23877 20640 23893 20704
rect 23957 20640 23973 20704
rect 24037 20640 24053 20704
rect 24117 20640 24125 20704
rect 23805 20639 24125 20640
rect 9805 20160 10125 20161
rect 9805 20096 9813 20160
rect 9877 20096 9893 20160
rect 9957 20096 9973 20160
rect 10037 20096 10053 20160
rect 10117 20096 10125 20160
rect 9805 20095 10125 20096
rect 19138 20160 19458 20161
rect 19138 20096 19146 20160
rect 19210 20096 19226 20160
rect 19290 20096 19306 20160
rect 19370 20096 19386 20160
rect 19450 20096 19458 20160
rect 19138 20095 19458 20096
rect 20517 20090 20583 20093
rect 27048 20090 27528 20120
rect 20517 20088 27528 20090
rect 20517 20032 20522 20088
rect 20578 20032 27528 20088
rect 20517 20030 27528 20032
rect 20517 20027 20583 20030
rect 27048 20000 27528 20030
rect 5138 19616 5458 19617
rect 5138 19552 5146 19616
rect 5210 19552 5226 19616
rect 5290 19552 5306 19616
rect 5370 19552 5386 19616
rect 5450 19552 5458 19616
rect 5138 19551 5458 19552
rect 14472 19616 14792 19617
rect 14472 19552 14480 19616
rect 14544 19552 14560 19616
rect 14624 19552 14640 19616
rect 14704 19552 14720 19616
rect 14784 19552 14792 19616
rect 14472 19551 14792 19552
rect 23805 19616 24125 19617
rect 23805 19552 23813 19616
rect 23877 19552 23893 19616
rect 23957 19552 23973 19616
rect 24037 19552 24053 19616
rect 24117 19552 24125 19616
rect 23805 19551 24125 19552
rect 20977 19410 21043 19413
rect 23001 19410 23067 19413
rect 20977 19408 23067 19410
rect 20977 19352 20982 19408
rect 21038 19352 23006 19408
rect 23062 19352 23067 19408
rect 20977 19350 23067 19352
rect 20977 19347 21043 19350
rect 23001 19347 23067 19350
rect 13249 19274 13315 19277
rect 23001 19274 23067 19277
rect 13249 19272 23067 19274
rect 13249 19216 13254 19272
rect 13310 19216 23006 19272
rect 23062 19216 23067 19272
rect 13249 19214 23067 19216
rect 13249 19211 13315 19214
rect 23001 19211 23067 19214
rect 24197 19138 24263 19141
rect 27048 19138 27528 19168
rect 24197 19136 27528 19138
rect 24197 19080 24202 19136
rect 24258 19080 27528 19136
rect 24197 19078 27528 19080
rect 24197 19075 24263 19078
rect 9805 19072 10125 19073
rect 9805 19008 9813 19072
rect 9877 19008 9893 19072
rect 9957 19008 9973 19072
rect 10037 19008 10053 19072
rect 10117 19008 10125 19072
rect 9805 19007 10125 19008
rect 19138 19072 19458 19073
rect 19138 19008 19146 19072
rect 19210 19008 19226 19072
rect 19290 19008 19306 19072
rect 19370 19008 19386 19072
rect 19450 19008 19458 19072
rect 27048 19048 27528 19078
rect 19138 19007 19458 19008
rect 10397 18730 10463 18733
rect 23001 18730 23067 18733
rect 10397 18728 23067 18730
rect 10397 18672 10402 18728
rect 10458 18672 23006 18728
rect 23062 18672 23067 18728
rect 10397 18670 23067 18672
rect 10397 18667 10463 18670
rect 23001 18667 23067 18670
rect 5138 18528 5458 18529
rect 5138 18464 5146 18528
rect 5210 18464 5226 18528
rect 5290 18464 5306 18528
rect 5370 18464 5386 18528
rect 5450 18464 5458 18528
rect 5138 18463 5458 18464
rect 14472 18528 14792 18529
rect 14472 18464 14480 18528
rect 14544 18464 14560 18528
rect 14624 18464 14640 18528
rect 14704 18464 14720 18528
rect 14784 18464 14792 18528
rect 14472 18463 14792 18464
rect 23805 18528 24125 18529
rect 23805 18464 23813 18528
rect 23877 18464 23893 18528
rect 23957 18464 23973 18528
rect 24037 18464 24053 18528
rect 24117 18464 24125 18528
rect 23805 18463 24125 18464
rect 16009 18322 16075 18325
rect 23093 18322 23159 18325
rect 16009 18320 23159 18322
rect 16009 18264 16014 18320
rect 16070 18264 23098 18320
rect 23154 18264 23159 18320
rect 16009 18262 23159 18264
rect 16009 18259 16075 18262
rect 23093 18259 23159 18262
rect 23553 18186 23619 18189
rect 25117 18186 25183 18189
rect 23553 18184 25183 18186
rect 23553 18128 23558 18184
rect 23614 18128 25122 18184
rect 25178 18128 25183 18184
rect 23553 18126 25183 18128
rect 23553 18123 23619 18126
rect 25117 18123 25183 18126
rect 8281 18050 8347 18053
rect 9569 18050 9635 18053
rect 8281 18048 9635 18050
rect 8281 17992 8286 18048
rect 8342 17992 9574 18048
rect 9630 17992 9635 18048
rect 8281 17990 9635 17992
rect 8281 17987 8347 17990
rect 9569 17987 9635 17990
rect 22633 18050 22699 18053
rect 27048 18050 27528 18080
rect 22633 18048 27528 18050
rect 22633 17992 22638 18048
rect 22694 17992 27528 18048
rect 22633 17990 27528 17992
rect 22633 17987 22699 17990
rect 9805 17984 10125 17985
rect 9805 17920 9813 17984
rect 9877 17920 9893 17984
rect 9957 17920 9973 17984
rect 10037 17920 10053 17984
rect 10117 17920 10125 17984
rect 9805 17919 10125 17920
rect 19138 17984 19458 17985
rect 19138 17920 19146 17984
rect 19210 17920 19226 17984
rect 19290 17920 19306 17984
rect 19370 17920 19386 17984
rect 19450 17920 19458 17984
rect 27048 17960 27528 17990
rect 19138 17919 19458 17920
rect 5138 17440 5458 17441
rect 5138 17376 5146 17440
rect 5210 17376 5226 17440
rect 5290 17376 5306 17440
rect 5370 17376 5386 17440
rect 5450 17376 5458 17440
rect 5138 17375 5458 17376
rect 14472 17440 14792 17441
rect 14472 17376 14480 17440
rect 14544 17376 14560 17440
rect 14624 17376 14640 17440
rect 14704 17376 14720 17440
rect 14784 17376 14792 17440
rect 14472 17375 14792 17376
rect 23805 17440 24125 17441
rect 23805 17376 23813 17440
rect 23877 17376 23893 17440
rect 23957 17376 23973 17440
rect 24037 17376 24053 17440
rect 24117 17376 24125 17440
rect 23805 17375 24125 17376
rect 17849 17370 17915 17373
rect 23461 17370 23527 17373
rect 17849 17368 23527 17370
rect 17849 17312 17854 17368
rect 17910 17312 23466 17368
rect 23522 17312 23527 17368
rect 17849 17310 23527 17312
rect 17849 17307 17915 17310
rect 23461 17307 23527 17310
rect 11593 17098 11659 17101
rect 24381 17098 24447 17101
rect 11593 17096 24447 17098
rect 11593 17040 11598 17096
rect 11654 17040 24386 17096
rect 24442 17040 24447 17096
rect 11593 17038 24447 17040
rect 11593 17035 11659 17038
rect 24381 17035 24447 17038
rect 25025 17098 25091 17101
rect 27048 17098 27528 17128
rect 25025 17096 27528 17098
rect 25025 17040 25030 17096
rect 25086 17040 27528 17096
rect 25025 17038 27528 17040
rect 25025 17035 25091 17038
rect 27048 17008 27528 17038
rect 9805 16896 10125 16897
rect 9805 16832 9813 16896
rect 9877 16832 9893 16896
rect 9957 16832 9973 16896
rect 10037 16832 10053 16896
rect 10117 16832 10125 16896
rect 9805 16831 10125 16832
rect 19138 16896 19458 16897
rect 19138 16832 19146 16896
rect 19210 16832 19226 16896
rect 19290 16832 19306 16896
rect 19370 16832 19386 16896
rect 19450 16832 19458 16896
rect 19138 16831 19458 16832
rect 12421 16690 12487 16693
rect 24381 16690 24447 16693
rect 12421 16688 24447 16690
rect 12421 16632 12426 16688
rect 12482 16632 24386 16688
rect 24442 16632 24447 16688
rect 12421 16630 24447 16632
rect 12421 16627 12487 16630
rect 24381 16627 24447 16630
rect 5138 16352 5458 16353
rect 5138 16288 5146 16352
rect 5210 16288 5226 16352
rect 5290 16288 5306 16352
rect 5370 16288 5386 16352
rect 5450 16288 5458 16352
rect 5138 16287 5458 16288
rect 14472 16352 14792 16353
rect 14472 16288 14480 16352
rect 14544 16288 14560 16352
rect 14624 16288 14640 16352
rect 14704 16288 14720 16352
rect 14784 16288 14792 16352
rect 14472 16287 14792 16288
rect 23805 16352 24125 16353
rect 23805 16288 23813 16352
rect 23877 16288 23893 16352
rect 23957 16288 23973 16352
rect 24037 16288 24053 16352
rect 24117 16288 24125 16352
rect 23805 16287 24125 16288
rect 5521 16146 5587 16149
rect 16837 16146 16903 16149
rect 5521 16144 16903 16146
rect 5521 16088 5526 16144
rect 5582 16088 16842 16144
rect 16898 16088 16903 16144
rect 5521 16086 16903 16088
rect 5521 16083 5587 16086
rect 16837 16083 16903 16086
rect 23277 16012 23343 16013
rect 23277 16010 23324 16012
rect 23232 16008 23324 16010
rect 23232 15952 23282 16008
rect 23232 15950 23324 15952
rect 23277 15948 23324 15950
rect 23388 15948 23394 16012
rect 23645 16010 23711 16013
rect 27048 16010 27528 16040
rect 23645 16008 27528 16010
rect 23645 15952 23650 16008
rect 23706 15952 27528 16008
rect 23645 15950 27528 15952
rect 23277 15947 23343 15948
rect 23645 15947 23711 15950
rect 27048 15920 27528 15950
rect 9805 15808 10125 15809
rect 9805 15744 9813 15808
rect 9877 15744 9893 15808
rect 9957 15744 9973 15808
rect 10037 15744 10053 15808
rect 10117 15744 10125 15808
rect 9805 15743 10125 15744
rect 19138 15808 19458 15809
rect 19138 15744 19146 15808
rect 19210 15744 19226 15808
rect 19290 15744 19306 15808
rect 19370 15744 19386 15808
rect 19450 15744 19458 15808
rect 19138 15743 19458 15744
rect 22265 15738 22331 15741
rect 24749 15738 24815 15741
rect 22265 15736 24815 15738
rect 22265 15680 22270 15736
rect 22326 15680 24754 15736
rect 24810 15680 24815 15736
rect 22265 15678 24815 15680
rect 22265 15675 22331 15678
rect 24749 15675 24815 15678
rect 13065 15602 13131 15605
rect 18953 15602 19019 15605
rect 13065 15600 19019 15602
rect 13065 15544 13070 15600
rect 13126 15544 18958 15600
rect 19014 15544 19019 15600
rect 13065 15542 19019 15544
rect 13065 15539 13131 15542
rect 18953 15539 19019 15542
rect 8189 15466 8255 15469
rect 20241 15466 20307 15469
rect 8189 15464 20307 15466
rect 8189 15408 8194 15464
rect 8250 15408 20246 15464
rect 20302 15408 20307 15464
rect 8189 15406 20307 15408
rect 8189 15403 8255 15406
rect 20241 15403 20307 15406
rect 18033 15330 18099 15333
rect 23001 15330 23067 15333
rect 18033 15328 23067 15330
rect 18033 15272 18038 15328
rect 18094 15272 23006 15328
rect 23062 15272 23067 15328
rect 18033 15270 23067 15272
rect 18033 15267 18099 15270
rect 23001 15267 23067 15270
rect 5138 15264 5458 15265
rect 5138 15200 5146 15264
rect 5210 15200 5226 15264
rect 5290 15200 5306 15264
rect 5370 15200 5386 15264
rect 5450 15200 5458 15264
rect 5138 15199 5458 15200
rect 14472 15264 14792 15265
rect 14472 15200 14480 15264
rect 14544 15200 14560 15264
rect 14624 15200 14640 15264
rect 14704 15200 14720 15264
rect 14784 15200 14792 15264
rect 14472 15199 14792 15200
rect 23805 15264 24125 15265
rect 23805 15200 23813 15264
rect 23877 15200 23893 15264
rect 23957 15200 23973 15264
rect 24037 15200 24053 15264
rect 24117 15200 24125 15264
rect 23805 15199 24125 15200
rect 24289 14922 24355 14925
rect 27048 14922 27528 14952
rect 24289 14920 27528 14922
rect 24289 14864 24294 14920
rect 24350 14864 27528 14920
rect 24289 14862 27528 14864
rect 24289 14859 24355 14862
rect 27048 14832 27528 14862
rect 14169 14786 14235 14789
rect 17941 14786 18007 14789
rect 14169 14784 18007 14786
rect 14169 14728 14174 14784
rect 14230 14728 17946 14784
rect 18002 14728 18007 14784
rect 14169 14726 18007 14728
rect 14169 14723 14235 14726
rect 17941 14723 18007 14726
rect 9805 14720 10125 14721
rect 9805 14656 9813 14720
rect 9877 14656 9893 14720
rect 9957 14656 9973 14720
rect 10037 14656 10053 14720
rect 10117 14656 10125 14720
rect 9805 14655 10125 14656
rect 19138 14720 19458 14721
rect 19138 14656 19146 14720
rect 19210 14656 19226 14720
rect 19290 14656 19306 14720
rect 19370 14656 19386 14720
rect 19450 14656 19458 14720
rect 19138 14655 19458 14656
rect 1013 14378 1079 14381
rect 8925 14378 8991 14381
rect 1013 14376 8991 14378
rect 1013 14320 1018 14376
rect 1074 14320 8930 14376
rect 8986 14320 8991 14376
rect 1013 14318 8991 14320
rect 1013 14315 1079 14318
rect 8925 14315 8991 14318
rect 22909 14378 22975 14381
rect 24841 14378 24907 14381
rect 22909 14376 24907 14378
rect 22909 14320 22914 14376
rect 22970 14320 24846 14376
rect 24902 14320 24907 14376
rect 22909 14318 24907 14320
rect 22909 14315 22975 14318
rect 24841 14315 24907 14318
rect 5138 14176 5458 14177
rect 5138 14112 5146 14176
rect 5210 14112 5226 14176
rect 5290 14112 5306 14176
rect 5370 14112 5386 14176
rect 5450 14112 5458 14176
rect 5138 14111 5458 14112
rect 14472 14176 14792 14177
rect 14472 14112 14480 14176
rect 14544 14112 14560 14176
rect 14624 14112 14640 14176
rect 14704 14112 14720 14176
rect 14784 14112 14792 14176
rect 14472 14111 14792 14112
rect 23805 14176 24125 14177
rect 23805 14112 23813 14176
rect 23877 14112 23893 14176
rect 23957 14112 23973 14176
rect 24037 14112 24053 14176
rect 24117 14112 24125 14176
rect 23805 14111 24125 14112
rect 13801 13970 13867 13973
rect 16377 13970 16443 13973
rect 13801 13968 16443 13970
rect 13801 13912 13806 13968
rect 13862 13912 16382 13968
rect 16438 13912 16443 13968
rect 13801 13910 16443 13912
rect 13801 13907 13867 13910
rect 16377 13907 16443 13910
rect 25393 13970 25459 13973
rect 27048 13970 27528 14000
rect 25393 13968 27528 13970
rect 25393 13912 25398 13968
rect 25454 13912 27528 13968
rect 25393 13910 27528 13912
rect 25393 13907 25459 13910
rect 27048 13880 27528 13910
rect 9805 13632 10125 13633
rect 9805 13568 9813 13632
rect 9877 13568 9893 13632
rect 9957 13568 9973 13632
rect 10037 13568 10053 13632
rect 10117 13568 10125 13632
rect 9805 13567 10125 13568
rect 19138 13632 19458 13633
rect 19138 13568 19146 13632
rect 19210 13568 19226 13632
rect 19290 13568 19306 13632
rect 19370 13568 19386 13632
rect 19450 13568 19458 13632
rect 19138 13567 19458 13568
rect 19597 13562 19663 13565
rect 21989 13562 22055 13565
rect 19597 13560 22055 13562
rect 19597 13504 19602 13560
rect 19658 13504 21994 13560
rect 22050 13504 22055 13560
rect 19597 13502 22055 13504
rect 19597 13499 19663 13502
rect 21989 13499 22055 13502
rect 24013 13562 24079 13565
rect 24473 13562 24539 13565
rect 24013 13560 24539 13562
rect 24013 13504 24018 13560
rect 24074 13504 24478 13560
rect 24534 13504 24539 13560
rect 24013 13502 24539 13504
rect 24013 13499 24079 13502
rect 24473 13499 24539 13502
rect 16469 13426 16535 13429
rect 22265 13426 22331 13429
rect 16469 13424 22331 13426
rect 16469 13368 16474 13424
rect 16530 13368 22270 13424
rect 22326 13368 22331 13424
rect 16469 13366 22331 13368
rect 16469 13363 16535 13366
rect 22265 13363 22331 13366
rect 23461 13426 23527 13429
rect 24289 13426 24355 13429
rect 23461 13424 24355 13426
rect 23461 13368 23466 13424
rect 23522 13368 24294 13424
rect 24350 13368 24355 13424
rect 23461 13366 24355 13368
rect 23461 13363 23527 13366
rect 24289 13363 24355 13366
rect 5138 13088 5458 13089
rect 5138 13024 5146 13088
rect 5210 13024 5226 13088
rect 5290 13024 5306 13088
rect 5370 13024 5386 13088
rect 5450 13024 5458 13088
rect 5138 13023 5458 13024
rect 14472 13088 14792 13089
rect 14472 13024 14480 13088
rect 14544 13024 14560 13088
rect 14624 13024 14640 13088
rect 14704 13024 14720 13088
rect 14784 13024 14792 13088
rect 14472 13023 14792 13024
rect 23805 13088 24125 13089
rect 23805 13024 23813 13088
rect 23877 13024 23893 13088
rect 23957 13024 23973 13088
rect 24037 13024 24053 13088
rect 24117 13024 24125 13088
rect 23805 13023 24125 13024
rect 9477 13018 9543 13021
rect 13985 13018 14051 13021
rect 9477 13016 14051 13018
rect 9477 12960 9482 13016
rect 9538 12960 13990 13016
rect 14046 12960 14051 13016
rect 9477 12958 14051 12960
rect 9477 12955 9543 12958
rect 13985 12955 14051 12958
rect 11685 12882 11751 12885
rect 17297 12882 17363 12885
rect 11685 12880 17363 12882
rect 11685 12824 11690 12880
rect 11746 12824 17302 12880
rect 17358 12824 17363 12880
rect 11685 12822 17363 12824
rect 11685 12819 11751 12822
rect 17297 12819 17363 12822
rect 24657 12882 24723 12885
rect 27048 12882 27528 12912
rect 24657 12880 27528 12882
rect 24657 12824 24662 12880
rect 24718 12824 27528 12880
rect 24657 12822 27528 12824
rect 24657 12819 24723 12822
rect 27048 12792 27528 12822
rect 5061 12746 5127 12749
rect 17941 12746 18007 12749
rect 5061 12744 18007 12746
rect 5061 12688 5066 12744
rect 5122 12688 17946 12744
rect 18002 12688 18007 12744
rect 5061 12686 18007 12688
rect 5061 12683 5127 12686
rect 17941 12683 18007 12686
rect 18309 12746 18375 12749
rect 20425 12746 20491 12749
rect 18309 12744 20491 12746
rect 18309 12688 18314 12744
rect 18370 12688 20430 12744
rect 20486 12688 20491 12744
rect 18309 12686 20491 12688
rect 18309 12683 18375 12686
rect 20425 12683 20491 12686
rect 21437 12746 21503 12749
rect 24473 12746 24539 12749
rect 21437 12744 24539 12746
rect 21437 12688 21442 12744
rect 21498 12688 24478 12744
rect 24534 12688 24539 12744
rect 21437 12686 24539 12688
rect 21437 12683 21503 12686
rect 24473 12683 24539 12686
rect 13065 12610 13131 12613
rect 18953 12610 19019 12613
rect 13065 12608 19019 12610
rect 13065 12552 13070 12608
rect 13126 12552 18958 12608
rect 19014 12552 19019 12608
rect 13065 12550 19019 12552
rect 13065 12547 13131 12550
rect 18953 12547 19019 12550
rect 22817 12610 22883 12613
rect 23277 12610 23343 12613
rect 23553 12610 23619 12613
rect 22817 12608 23343 12610
rect 22817 12552 22822 12608
rect 22878 12552 23282 12608
rect 23338 12552 23343 12608
rect 22817 12550 23343 12552
rect 22817 12547 22883 12550
rect 23277 12547 23343 12550
rect 23510 12608 23619 12610
rect 23510 12552 23558 12608
rect 23614 12552 23619 12608
rect 23510 12547 23619 12552
rect 9805 12544 10125 12545
rect 9805 12480 9813 12544
rect 9877 12480 9893 12544
rect 9957 12480 9973 12544
rect 10037 12480 10053 12544
rect 10117 12480 10125 12544
rect 9805 12479 10125 12480
rect 19138 12544 19458 12545
rect 19138 12480 19146 12544
rect 19210 12480 19226 12544
rect 19290 12480 19306 12544
rect 19370 12480 19386 12544
rect 19450 12480 19458 12544
rect 19138 12479 19458 12480
rect 11869 12474 11935 12477
rect 12513 12474 12579 12477
rect 16653 12474 16719 12477
rect 11869 12472 16719 12474
rect 11869 12416 11874 12472
rect 11930 12416 12518 12472
rect 12574 12416 16658 12472
rect 16714 12416 16719 12472
rect 11869 12414 16719 12416
rect 11869 12411 11935 12414
rect 12513 12411 12579 12414
rect 16653 12411 16719 12414
rect 22817 12474 22883 12477
rect 23510 12474 23570 12547
rect 22817 12472 23570 12474
rect 22817 12416 22822 12472
rect 22878 12416 23570 12472
rect 22817 12414 23570 12416
rect 22817 12411 22883 12414
rect 9385 12338 9451 12341
rect 13433 12338 13499 12341
rect 15181 12338 15247 12341
rect 17573 12338 17639 12341
rect 18493 12338 18559 12341
rect 9385 12336 18559 12338
rect 9385 12280 9390 12336
rect 9446 12280 13438 12336
rect 13494 12280 15186 12336
rect 15242 12280 17578 12336
rect 17634 12280 18498 12336
rect 18554 12280 18559 12336
rect 9385 12278 18559 12280
rect 9385 12275 9451 12278
rect 13433 12275 13499 12278
rect 15181 12275 15247 12278
rect 17573 12275 17639 12278
rect 18493 12275 18559 12278
rect 20425 12338 20491 12341
rect 22633 12338 22699 12341
rect 20425 12336 22699 12338
rect 20425 12280 20430 12336
rect 20486 12280 22638 12336
rect 22694 12280 22699 12336
rect 20425 12278 22699 12280
rect 20425 12275 20491 12278
rect 22633 12275 22699 12278
rect 11409 12202 11475 12205
rect 12329 12202 12395 12205
rect 14261 12202 14327 12205
rect 14537 12202 14603 12205
rect 17297 12202 17363 12205
rect 23369 12204 23435 12205
rect 23318 12202 23324 12204
rect 11409 12200 17363 12202
rect 11409 12144 11414 12200
rect 11470 12144 12334 12200
rect 12390 12144 14266 12200
rect 14322 12144 14542 12200
rect 14598 12144 17302 12200
rect 17358 12144 17363 12200
rect 11409 12142 17363 12144
rect 23278 12142 23324 12202
rect 23388 12200 23435 12204
rect 23430 12144 23435 12200
rect 11409 12139 11475 12142
rect 12329 12139 12395 12142
rect 14261 12139 14327 12142
rect 14537 12139 14603 12142
rect 17297 12139 17363 12142
rect 23318 12140 23324 12142
rect 23388 12140 23435 12144
rect 23369 12139 23435 12140
rect 7729 12066 7795 12069
rect 13617 12066 13683 12069
rect 7729 12064 13683 12066
rect 7729 12008 7734 12064
rect 7790 12008 13622 12064
rect 13678 12008 13683 12064
rect 7729 12006 13683 12008
rect 7729 12003 7795 12006
rect 13617 12003 13683 12006
rect 5138 12000 5458 12001
rect 5138 11936 5146 12000
rect 5210 11936 5226 12000
rect 5290 11936 5306 12000
rect 5370 11936 5386 12000
rect 5450 11936 5458 12000
rect 5138 11935 5458 11936
rect 14472 12000 14792 12001
rect 14472 11936 14480 12000
rect 14544 11936 14560 12000
rect 14624 11936 14640 12000
rect 14704 11936 14720 12000
rect 14784 11936 14792 12000
rect 14472 11935 14792 11936
rect 23805 12000 24125 12001
rect 23805 11936 23813 12000
rect 23877 11936 23893 12000
rect 23957 11936 23973 12000
rect 24037 11936 24053 12000
rect 24117 11936 24125 12000
rect 23805 11935 24125 11936
rect 8649 11930 8715 11933
rect 11133 11930 11199 11933
rect 8649 11928 11199 11930
rect 8649 11872 8654 11928
rect 8710 11872 11138 11928
rect 11194 11872 11199 11928
rect 8649 11870 11199 11872
rect 8649 11867 8715 11870
rect 11133 11867 11199 11870
rect 8281 11794 8347 11797
rect 13893 11794 13959 11797
rect 8281 11792 13959 11794
rect 8281 11736 8286 11792
rect 8342 11736 13898 11792
rect 13954 11736 13959 11792
rect 8281 11734 13959 11736
rect 8281 11731 8347 11734
rect 13893 11731 13959 11734
rect 17665 11794 17731 11797
rect 23645 11794 23711 11797
rect 17665 11792 23711 11794
rect 17665 11736 17670 11792
rect 17726 11736 23650 11792
rect 23706 11736 23711 11792
rect 17665 11734 23711 11736
rect 17665 11731 17731 11734
rect 23645 11731 23711 11734
rect 25485 11794 25551 11797
rect 27048 11794 27528 11824
rect 25485 11792 27528 11794
rect 25485 11736 25490 11792
rect 25546 11736 27528 11792
rect 25485 11734 27528 11736
rect 25485 11731 25551 11734
rect 27048 11704 27528 11734
rect 14997 11658 15063 11661
rect 18217 11658 18283 11661
rect 14997 11656 18283 11658
rect 14997 11600 15002 11656
rect 15058 11600 18222 11656
rect 18278 11600 18283 11656
rect 14997 11598 18283 11600
rect 14997 11595 15063 11598
rect 18217 11595 18283 11598
rect 18769 11658 18835 11661
rect 24841 11658 24907 11661
rect 18769 11656 24907 11658
rect 18769 11600 18774 11656
rect 18830 11600 24846 11656
rect 24902 11600 24907 11656
rect 18769 11598 24907 11600
rect 18769 11595 18835 11598
rect 24841 11595 24907 11598
rect 10673 11522 10739 11525
rect 16745 11522 16811 11525
rect 10673 11520 16811 11522
rect 10673 11464 10678 11520
rect 10734 11464 16750 11520
rect 16806 11464 16811 11520
rect 10673 11462 16811 11464
rect 10673 11459 10739 11462
rect 16745 11459 16811 11462
rect 9805 11456 10125 11457
rect 9805 11392 9813 11456
rect 9877 11392 9893 11456
rect 9957 11392 9973 11456
rect 10037 11392 10053 11456
rect 10117 11392 10125 11456
rect 9805 11391 10125 11392
rect 19138 11456 19458 11457
rect 19138 11392 19146 11456
rect 19210 11392 19226 11456
rect 19290 11392 19306 11456
rect 19370 11392 19386 11456
rect 19450 11392 19458 11456
rect 19138 11391 19458 11392
rect 3681 11250 3747 11253
rect 8097 11250 8163 11253
rect 3681 11248 8163 11250
rect 3681 11192 3686 11248
rect 3742 11192 8102 11248
rect 8158 11192 8163 11248
rect 3681 11190 8163 11192
rect 3681 11187 3747 11190
rect 8097 11187 8163 11190
rect 13249 11250 13315 11253
rect 20333 11250 20399 11253
rect 13249 11248 20399 11250
rect 13249 11192 13254 11248
rect 13310 11192 20338 11248
rect 20394 11192 20399 11248
rect 13249 11190 20399 11192
rect 13249 11187 13315 11190
rect 20333 11187 20399 11190
rect 8281 11114 8347 11117
rect 20425 11114 20491 11117
rect 8281 11112 20491 11114
rect 8281 11056 8286 11112
rect 8342 11056 20430 11112
rect 20486 11056 20491 11112
rect 8281 11054 20491 11056
rect 8281 11051 8347 11054
rect 20425 11051 20491 11054
rect 5138 10912 5458 10913
rect 5138 10848 5146 10912
rect 5210 10848 5226 10912
rect 5290 10848 5306 10912
rect 5370 10848 5386 10912
rect 5450 10848 5458 10912
rect 5138 10847 5458 10848
rect 14472 10912 14792 10913
rect 14472 10848 14480 10912
rect 14544 10848 14560 10912
rect 14624 10848 14640 10912
rect 14704 10848 14720 10912
rect 14784 10848 14792 10912
rect 14472 10847 14792 10848
rect 23805 10912 24125 10913
rect 23805 10848 23813 10912
rect 23877 10848 23893 10912
rect 23957 10848 23973 10912
rect 24037 10848 24053 10912
rect 24117 10848 24125 10912
rect 23805 10847 24125 10848
rect 7361 10842 7427 10845
rect 13801 10842 13867 10845
rect 7361 10840 13867 10842
rect 7361 10784 7366 10840
rect 7422 10784 13806 10840
rect 13862 10784 13867 10840
rect 7361 10782 13867 10784
rect 7361 10779 7427 10782
rect 13801 10779 13867 10782
rect 24197 10842 24263 10845
rect 27048 10842 27528 10872
rect 24197 10840 27528 10842
rect 24197 10784 24202 10840
rect 24258 10784 27528 10840
rect 24197 10782 27528 10784
rect 24197 10779 24263 10782
rect 27048 10752 27528 10782
rect 8465 10706 8531 10709
rect 20609 10706 20675 10709
rect 24381 10706 24447 10709
rect 8465 10704 24447 10706
rect 8465 10648 8470 10704
rect 8526 10648 20614 10704
rect 20670 10648 24386 10704
rect 24442 10648 24447 10704
rect 8465 10646 24447 10648
rect 8465 10643 8531 10646
rect 20609 10643 20675 10646
rect 24381 10643 24447 10646
rect 4417 10570 4483 10573
rect 10673 10570 10739 10573
rect 4417 10568 10739 10570
rect 4417 10512 4422 10568
rect 4478 10512 10678 10568
rect 10734 10512 10739 10568
rect 4417 10510 10739 10512
rect 4417 10507 4483 10510
rect 10673 10507 10739 10510
rect 13341 10570 13407 10573
rect 17205 10570 17271 10573
rect 13341 10568 17271 10570
rect 13341 10512 13346 10568
rect 13402 10512 17210 10568
rect 17266 10512 17271 10568
rect 13341 10510 17271 10512
rect 13341 10507 13407 10510
rect 17205 10507 17271 10510
rect 18309 10570 18375 10573
rect 22541 10570 22607 10573
rect 18309 10568 22607 10570
rect 18309 10512 18314 10568
rect 18370 10512 22546 10568
rect 22602 10512 22607 10568
rect 18309 10510 22607 10512
rect 18309 10507 18375 10510
rect 22541 10507 22607 10510
rect 19597 10434 19663 10437
rect 24933 10434 24999 10437
rect 19597 10432 24999 10434
rect 19597 10376 19602 10432
rect 19658 10376 24938 10432
rect 24994 10376 24999 10432
rect 19597 10374 24999 10376
rect 19597 10371 19663 10374
rect 24933 10371 24999 10374
rect 9805 10368 10125 10369
rect 9805 10304 9813 10368
rect 9877 10304 9893 10368
rect 9957 10304 9973 10368
rect 10037 10304 10053 10368
rect 10117 10304 10125 10368
rect 9805 10303 10125 10304
rect 19138 10368 19458 10369
rect 19138 10304 19146 10368
rect 19210 10304 19226 10368
rect 19290 10304 19306 10368
rect 19370 10304 19386 10368
rect 19450 10304 19458 10368
rect 19138 10303 19458 10304
rect 14629 10298 14695 10301
rect 16193 10298 16259 10301
rect 14629 10296 16259 10298
rect 14629 10240 14634 10296
rect 14690 10240 16198 10296
rect 16254 10240 16259 10296
rect 14629 10238 16259 10240
rect 14629 10235 14695 10238
rect 16193 10235 16259 10238
rect 9477 10162 9543 10165
rect 13985 10162 14051 10165
rect 15365 10162 15431 10165
rect 9477 10160 14051 10162
rect 9477 10104 9482 10160
rect 9538 10104 13990 10160
rect 14046 10104 14051 10160
rect 9477 10102 14051 10104
rect 9477 10099 9543 10102
rect 13985 10099 14051 10102
rect 14126 10160 15431 10162
rect 14126 10104 15370 10160
rect 15426 10104 15431 10160
rect 14126 10102 15431 10104
rect 9661 10026 9727 10029
rect 14126 10026 14186 10102
rect 15365 10099 15431 10102
rect 22449 10026 22515 10029
rect 9661 10024 14186 10026
rect 9661 9968 9666 10024
rect 9722 9968 14186 10024
rect 9661 9966 14186 9968
rect 14310 10024 22515 10026
rect 14310 9968 22454 10024
rect 22510 9968 22515 10024
rect 14310 9966 22515 9968
rect 9661 9963 9727 9966
rect 8373 9890 8439 9893
rect 13433 9890 13499 9893
rect 8373 9888 13499 9890
rect 8373 9832 8378 9888
rect 8434 9832 13438 9888
rect 13494 9832 13499 9888
rect 8373 9830 13499 9832
rect 8373 9827 8439 9830
rect 13433 9827 13499 9830
rect 5138 9824 5458 9825
rect 5138 9760 5146 9824
rect 5210 9760 5226 9824
rect 5290 9760 5306 9824
rect 5370 9760 5386 9824
rect 5450 9760 5458 9824
rect 5138 9759 5458 9760
rect 9661 9754 9727 9757
rect 14310 9754 14370 9966
rect 22449 9963 22515 9966
rect 15549 9890 15615 9893
rect 17849 9890 17915 9893
rect 15549 9888 17915 9890
rect 15549 9832 15554 9888
rect 15610 9832 17854 9888
rect 17910 9832 17915 9888
rect 15549 9830 17915 9832
rect 15549 9827 15615 9830
rect 17849 9827 17915 9830
rect 14472 9824 14792 9825
rect 14472 9760 14480 9824
rect 14544 9760 14560 9824
rect 14624 9760 14640 9824
rect 14704 9760 14720 9824
rect 14784 9760 14792 9824
rect 14472 9759 14792 9760
rect 23805 9824 24125 9825
rect 23805 9760 23813 9824
rect 23877 9760 23893 9824
rect 23957 9760 23973 9824
rect 24037 9760 24053 9824
rect 24117 9760 24125 9824
rect 23805 9759 24125 9760
rect 9661 9752 14370 9754
rect 9661 9696 9666 9752
rect 9722 9696 14370 9752
rect 9661 9694 14370 9696
rect 24933 9754 24999 9757
rect 27048 9754 27528 9784
rect 24933 9752 27528 9754
rect 24933 9696 24938 9752
rect 24994 9696 27528 9752
rect 24933 9694 27528 9696
rect 9661 9691 9727 9694
rect 24933 9691 24999 9694
rect 27048 9664 27528 9694
rect 8373 9618 8439 9621
rect 13249 9618 13315 9621
rect 8373 9616 13315 9618
rect 8373 9560 8378 9616
rect 8434 9560 13254 9616
rect 13310 9560 13315 9616
rect 8373 9558 13315 9560
rect 8373 9555 8439 9558
rect 13249 9555 13315 9558
rect 17665 9618 17731 9621
rect 17665 9616 24674 9618
rect 17665 9560 17670 9616
rect 17726 9560 24674 9616
rect 17665 9558 24674 9560
rect 17665 9555 17731 9558
rect 7821 9482 7887 9485
rect 23921 9482 23987 9485
rect 7821 9480 23987 9482
rect 7821 9424 7826 9480
rect 7882 9424 23926 9480
rect 23982 9424 23987 9480
rect 7821 9422 23987 9424
rect 24614 9482 24674 9558
rect 24841 9482 24907 9485
rect 24614 9480 24907 9482
rect 24614 9424 24846 9480
rect 24902 9424 24907 9480
rect 24614 9422 24907 9424
rect 7821 9419 7887 9422
rect 23921 9419 23987 9422
rect 24841 9419 24907 9422
rect 9805 9280 10125 9281
rect 9805 9216 9813 9280
rect 9877 9216 9893 9280
rect 9957 9216 9973 9280
rect 10037 9216 10053 9280
rect 10117 9216 10125 9280
rect 9805 9215 10125 9216
rect 19138 9280 19458 9281
rect 19138 9216 19146 9280
rect 19210 9216 19226 9280
rect 19290 9216 19306 9280
rect 19370 9216 19386 9280
rect 19450 9216 19458 9280
rect 19138 9215 19458 9216
rect 6441 9074 6507 9077
rect 16837 9074 16903 9077
rect 25209 9074 25275 9077
rect 6441 9072 15612 9074
rect 6441 9016 6446 9072
rect 6502 9016 15612 9072
rect 6441 9014 15612 9016
rect 6441 9011 6507 9014
rect 5981 8938 6047 8941
rect 12697 8938 12763 8941
rect 13341 8938 13407 8941
rect 15089 8938 15155 8941
rect 5981 8936 13407 8938
rect 5981 8880 5986 8936
rect 6042 8880 12702 8936
rect 12758 8880 13346 8936
rect 13402 8880 13407 8936
rect 5981 8878 13407 8880
rect 5981 8875 6047 8878
rect 12697 8875 12763 8878
rect 13341 8875 13407 8878
rect 13574 8936 15155 8938
rect 13574 8880 15094 8936
rect 15150 8880 15155 8936
rect 13574 8878 15155 8880
rect 15552 8938 15612 9014
rect 16837 9072 25275 9074
rect 16837 9016 16842 9072
rect 16898 9016 25214 9072
rect 25270 9016 25275 9072
rect 16837 9014 25275 9016
rect 16837 9011 16903 9014
rect 25209 9011 25275 9014
rect 17849 8938 17915 8941
rect 15552 8936 17915 8938
rect 15552 8880 17854 8936
rect 17910 8880 17915 8936
rect 15552 8878 17915 8880
rect 5797 8802 5863 8805
rect 13574 8802 13634 8878
rect 15089 8875 15155 8878
rect 17849 8875 17915 8878
rect 23737 8938 23803 8941
rect 23737 8936 24306 8938
rect 23737 8880 23742 8936
rect 23798 8880 24306 8936
rect 23737 8878 24306 8880
rect 23737 8875 23803 8878
rect 5797 8800 13634 8802
rect 5797 8744 5802 8800
rect 5858 8744 13634 8800
rect 5797 8742 13634 8744
rect 19045 8802 19111 8805
rect 20885 8802 20951 8805
rect 19045 8800 20951 8802
rect 19045 8744 19050 8800
rect 19106 8744 20890 8800
rect 20946 8744 20951 8800
rect 19045 8742 20951 8744
rect 24246 8802 24306 8878
rect 27048 8802 27528 8832
rect 24246 8742 27528 8802
rect 5797 8739 5863 8742
rect 19045 8739 19111 8742
rect 20885 8739 20951 8742
rect 5138 8736 5458 8737
rect 5138 8672 5146 8736
rect 5210 8672 5226 8736
rect 5290 8672 5306 8736
rect 5370 8672 5386 8736
rect 5450 8672 5458 8736
rect 5138 8671 5458 8672
rect 14472 8736 14792 8737
rect 14472 8672 14480 8736
rect 14544 8672 14560 8736
rect 14624 8672 14640 8736
rect 14704 8672 14720 8736
rect 14784 8672 14792 8736
rect 14472 8671 14792 8672
rect 23805 8736 24125 8737
rect 23805 8672 23813 8736
rect 23877 8672 23893 8736
rect 23957 8672 23973 8736
rect 24037 8672 24053 8736
rect 24117 8672 24125 8736
rect 27048 8712 27528 8742
rect 23805 8671 24125 8672
rect 10397 8666 10463 8669
rect 12605 8666 12671 8669
rect 10397 8664 12671 8666
rect 10397 8608 10402 8664
rect 10458 8608 12610 8664
rect 12666 8608 12671 8664
rect 10397 8606 12671 8608
rect 10397 8603 10463 8606
rect 12605 8603 12671 8606
rect 20425 8666 20491 8669
rect 23185 8666 23251 8669
rect 20425 8664 23251 8666
rect 20425 8608 20430 8664
rect 20486 8608 23190 8664
rect 23246 8608 23251 8664
rect 20425 8606 23251 8608
rect 20425 8603 20491 8606
rect 23185 8603 23251 8606
rect 12329 8530 12395 8533
rect 24749 8530 24815 8533
rect 12329 8528 24815 8530
rect 12329 8472 12334 8528
rect 12390 8472 24754 8528
rect 24810 8472 24815 8528
rect 12329 8470 24815 8472
rect 12329 8467 12395 8470
rect 24749 8467 24815 8470
rect 8925 8394 8991 8397
rect 23277 8394 23343 8397
rect 8925 8392 23343 8394
rect 8925 8336 8930 8392
rect 8986 8336 23282 8392
rect 23338 8336 23343 8392
rect 8925 8334 23343 8336
rect 8925 8331 8991 8334
rect 23277 8331 23343 8334
rect 3313 8258 3379 8261
rect 9477 8258 9543 8261
rect 3313 8256 9543 8258
rect 3313 8200 3318 8256
rect 3374 8200 9482 8256
rect 9538 8200 9543 8256
rect 3313 8198 9543 8200
rect 3313 8195 3379 8198
rect 9477 8195 9543 8198
rect 10765 8258 10831 8261
rect 13893 8258 13959 8261
rect 10765 8256 13959 8258
rect 10765 8200 10770 8256
rect 10826 8200 13898 8256
rect 13954 8200 13959 8256
rect 10765 8198 13959 8200
rect 10765 8195 10831 8198
rect 13893 8195 13959 8198
rect 14629 8258 14695 8261
rect 17757 8258 17823 8261
rect 14629 8256 17823 8258
rect 14629 8200 14634 8256
rect 14690 8200 17762 8256
rect 17818 8200 17823 8256
rect 14629 8198 17823 8200
rect 14629 8195 14695 8198
rect 17757 8195 17823 8198
rect 9805 8192 10125 8193
rect 9805 8128 9813 8192
rect 9877 8128 9893 8192
rect 9957 8128 9973 8192
rect 10037 8128 10053 8192
rect 10117 8128 10125 8192
rect 9805 8127 10125 8128
rect 19138 8192 19458 8193
rect 19138 8128 19146 8192
rect 19210 8128 19226 8192
rect 19290 8128 19306 8192
rect 19370 8128 19386 8192
rect 19450 8128 19458 8192
rect 19138 8127 19458 8128
rect 10213 8122 10279 8125
rect 10213 8120 16762 8122
rect 10213 8064 10218 8120
rect 10274 8064 16762 8120
rect 10213 8062 16762 8064
rect 10213 8059 10279 8062
rect 8189 7986 8255 7989
rect 16561 7986 16627 7989
rect 8189 7984 16627 7986
rect 8189 7928 8194 7984
rect 8250 7928 16566 7984
rect 16622 7928 16627 7984
rect 8189 7926 16627 7928
rect 16702 7986 16762 8062
rect 21621 7986 21687 7989
rect 16702 7984 21687 7986
rect 16702 7928 21626 7984
rect 21682 7928 21687 7984
rect 16702 7926 21687 7928
rect 8189 7923 8255 7926
rect 16561 7923 16627 7926
rect 21621 7923 21687 7926
rect 7729 7852 7795 7853
rect 7678 7788 7684 7852
rect 7748 7850 7795 7852
rect 8281 7850 8347 7853
rect 21621 7850 21687 7853
rect 7748 7848 7840 7850
rect 7790 7792 7840 7848
rect 7748 7790 7840 7792
rect 8281 7848 21687 7850
rect 8281 7792 8286 7848
rect 8342 7792 21626 7848
rect 21682 7792 21687 7848
rect 8281 7790 21687 7792
rect 7748 7788 7795 7790
rect 7729 7787 7795 7788
rect 8281 7787 8347 7790
rect 21621 7787 21687 7790
rect 8649 7714 8715 7717
rect 10213 7714 10279 7717
rect 8649 7712 10279 7714
rect 8649 7656 8654 7712
rect 8710 7656 10218 7712
rect 10274 7656 10279 7712
rect 8649 7654 10279 7656
rect 8649 7651 8715 7654
rect 10213 7651 10279 7654
rect 16561 7714 16627 7717
rect 21345 7714 21411 7717
rect 16561 7712 21411 7714
rect 16561 7656 16566 7712
rect 16622 7656 21350 7712
rect 21406 7656 21411 7712
rect 16561 7654 21411 7656
rect 16561 7651 16627 7654
rect 21345 7651 21411 7654
rect 25301 7714 25367 7717
rect 27048 7714 27528 7744
rect 25301 7712 27528 7714
rect 25301 7656 25306 7712
rect 25362 7656 27528 7712
rect 25301 7654 27528 7656
rect 25301 7651 25367 7654
rect 5138 7648 5458 7649
rect 5138 7584 5146 7648
rect 5210 7584 5226 7648
rect 5290 7584 5306 7648
rect 5370 7584 5386 7648
rect 5450 7584 5458 7648
rect 5138 7583 5458 7584
rect 14472 7648 14792 7649
rect 14472 7584 14480 7648
rect 14544 7584 14560 7648
rect 14624 7584 14640 7648
rect 14704 7584 14720 7648
rect 14784 7584 14792 7648
rect 14472 7583 14792 7584
rect 23805 7648 24125 7649
rect 23805 7584 23813 7648
rect 23877 7584 23893 7648
rect 23957 7584 23973 7648
rect 24037 7584 24053 7648
rect 24117 7584 24125 7648
rect 27048 7624 27528 7654
rect 23805 7583 24125 7584
rect 9293 7442 9359 7445
rect 10857 7442 10923 7445
rect 12145 7442 12211 7445
rect 9293 7440 12211 7442
rect 9293 7384 9298 7440
rect 9354 7384 10862 7440
rect 10918 7384 12150 7440
rect 12206 7384 12211 7440
rect 9293 7382 12211 7384
rect 9293 7379 9359 7382
rect 10857 7379 10923 7382
rect 12145 7379 12211 7382
rect 13893 7442 13959 7445
rect 17849 7442 17915 7445
rect 13893 7440 17915 7442
rect 13893 7384 13898 7440
rect 13954 7384 17854 7440
rect 17910 7384 17915 7440
rect 13893 7382 17915 7384
rect 13893 7379 13959 7382
rect 17849 7379 17915 7382
rect 21253 7442 21319 7445
rect 23737 7442 23803 7445
rect 21253 7440 23803 7442
rect 21253 7384 21258 7440
rect 21314 7384 23742 7440
rect 23798 7384 23803 7440
rect 21253 7382 23803 7384
rect 21253 7379 21319 7382
rect 23737 7379 23803 7382
rect 8097 7306 8163 7309
rect 18125 7306 18191 7309
rect 8097 7304 18191 7306
rect 8097 7248 8102 7304
rect 8158 7248 18130 7304
rect 18186 7248 18191 7304
rect 8097 7246 18191 7248
rect 8097 7243 8163 7246
rect 18125 7243 18191 7246
rect 20609 7306 20675 7309
rect 24749 7306 24815 7309
rect 20609 7304 24815 7306
rect 20609 7248 20614 7304
rect 20670 7248 24754 7304
rect 24810 7248 24815 7304
rect 20609 7246 24815 7248
rect 20609 7243 20675 7246
rect 24749 7243 24815 7246
rect 1657 7170 1723 7173
rect 7821 7170 7887 7173
rect 1657 7168 7887 7170
rect 1657 7112 1662 7168
rect 1718 7112 7826 7168
rect 7882 7112 7887 7168
rect 1657 7110 7887 7112
rect 1657 7107 1723 7110
rect 7821 7107 7887 7110
rect 10397 7170 10463 7173
rect 12513 7170 12579 7173
rect 18401 7170 18467 7173
rect 10397 7168 12346 7170
rect 10397 7112 10402 7168
rect 10458 7112 12346 7168
rect 10397 7110 12346 7112
rect 10397 7107 10463 7110
rect 9805 7104 10125 7105
rect 9805 7040 9813 7104
rect 9877 7040 9893 7104
rect 9957 7040 9973 7104
rect 10037 7040 10053 7104
rect 10117 7040 10125 7104
rect 9805 7039 10125 7040
rect 2761 7034 2827 7037
rect 6441 7034 6507 7037
rect 2761 7032 6507 7034
rect 2761 6976 2766 7032
rect 2822 6976 6446 7032
rect 6502 6976 6507 7032
rect 2761 6974 6507 6976
rect 2761 6971 2827 6974
rect 6441 6971 6507 6974
rect 10213 7034 10279 7037
rect 12053 7034 12119 7037
rect 10213 7032 12119 7034
rect 10213 6976 10218 7032
rect 10274 6976 12058 7032
rect 12114 6976 12119 7032
rect 10213 6974 12119 6976
rect 12286 7034 12346 7110
rect 12513 7168 18467 7170
rect 12513 7112 12518 7168
rect 12574 7112 18406 7168
rect 18462 7112 18467 7168
rect 12513 7110 18467 7112
rect 12513 7107 12579 7110
rect 18401 7107 18467 7110
rect 19138 7104 19458 7105
rect 19138 7040 19146 7104
rect 19210 7040 19226 7104
rect 19290 7040 19306 7104
rect 19370 7040 19386 7104
rect 19450 7040 19458 7104
rect 19138 7039 19458 7040
rect 16653 7034 16719 7037
rect 12286 7032 16719 7034
rect 12286 6976 16658 7032
rect 16714 6976 16719 7032
rect 12286 6974 16719 6976
rect 10213 6971 10279 6974
rect 12053 6971 12119 6974
rect 16653 6971 16719 6974
rect 13341 6898 13407 6901
rect 16101 6898 16167 6901
rect 13341 6896 16167 6898
rect 13341 6840 13346 6896
rect 13402 6840 16106 6896
rect 16162 6840 16167 6896
rect 13341 6838 16167 6840
rect 13341 6835 13407 6838
rect 16101 6835 16167 6838
rect 22950 6836 22956 6900
rect 23020 6898 23026 6900
rect 23093 6898 23159 6901
rect 23020 6896 23159 6898
rect 23020 6840 23098 6896
rect 23154 6840 23159 6896
rect 23020 6838 23159 6840
rect 23020 6836 23026 6838
rect 23093 6835 23159 6838
rect 3773 6762 3839 6765
rect 10857 6762 10923 6765
rect 3773 6760 10923 6762
rect 3773 6704 3778 6760
rect 3834 6704 10862 6760
rect 10918 6704 10923 6760
rect 3773 6702 10923 6704
rect 3773 6699 3839 6702
rect 10857 6699 10923 6702
rect 11777 6762 11843 6765
rect 23553 6762 23619 6765
rect 11777 6760 23619 6762
rect 11777 6704 11782 6760
rect 11838 6704 23558 6760
rect 23614 6704 23619 6760
rect 11777 6702 23619 6704
rect 11777 6699 11843 6702
rect 23553 6699 23619 6702
rect 24289 6626 24355 6629
rect 27048 6626 27528 6656
rect 24289 6624 27528 6626
rect 24289 6568 24294 6624
rect 24350 6568 27528 6624
rect 24289 6566 27528 6568
rect 24289 6563 24355 6566
rect 5138 6560 5458 6561
rect 5138 6496 5146 6560
rect 5210 6496 5226 6560
rect 5290 6496 5306 6560
rect 5370 6496 5386 6560
rect 5450 6496 5458 6560
rect 5138 6495 5458 6496
rect 14472 6560 14792 6561
rect 14472 6496 14480 6560
rect 14544 6496 14560 6560
rect 14624 6496 14640 6560
rect 14704 6496 14720 6560
rect 14784 6496 14792 6560
rect 14472 6495 14792 6496
rect 23805 6560 24125 6561
rect 23805 6496 23813 6560
rect 23877 6496 23893 6560
rect 23957 6496 23973 6560
rect 24037 6496 24053 6560
rect 24117 6496 24125 6560
rect 27048 6536 27528 6566
rect 23805 6495 24125 6496
rect 4049 6490 4115 6493
rect 4182 6490 4188 6492
rect 4049 6488 4188 6490
rect 4049 6432 4054 6488
rect 4110 6432 4188 6488
rect 4049 6430 4188 6432
rect 4049 6427 4115 6430
rect 4182 6428 4188 6430
rect 4252 6428 4258 6492
rect 6533 6490 6599 6493
rect 13249 6490 13315 6493
rect 6533 6488 13315 6490
rect 6533 6432 6538 6488
rect 6594 6432 13254 6488
rect 13310 6432 13315 6488
rect 6533 6430 13315 6432
rect 6533 6427 6599 6430
rect 13249 6427 13315 6430
rect 24422 6428 24428 6492
rect 24492 6490 24498 6492
rect 24565 6490 24631 6493
rect 24492 6488 24631 6490
rect 24492 6432 24570 6488
rect 24626 6432 24631 6488
rect 24492 6430 24631 6432
rect 24492 6428 24498 6430
rect 24565 6427 24631 6430
rect 8097 6354 8163 6357
rect 10254 6354 10260 6356
rect 8097 6352 10260 6354
rect 8097 6296 8102 6352
rect 8158 6296 10260 6352
rect 8097 6294 10260 6296
rect 8097 6291 8163 6294
rect 10254 6292 10260 6294
rect 10324 6292 10330 6356
rect 10857 6354 10923 6357
rect 16285 6354 16351 6357
rect 10857 6352 16351 6354
rect 10857 6296 10862 6352
rect 10918 6296 16290 6352
rect 16346 6296 16351 6352
rect 10857 6294 16351 6296
rect 10857 6291 10923 6294
rect 16285 6291 16351 6294
rect 7729 6218 7795 6221
rect 24749 6218 24815 6221
rect 7729 6216 24815 6218
rect 7729 6160 7734 6216
rect 7790 6160 24754 6216
rect 24810 6160 24815 6216
rect 7729 6158 24815 6160
rect 7729 6155 7795 6158
rect 24749 6155 24815 6158
rect 10397 6082 10463 6085
rect 18953 6082 19019 6085
rect 10397 6080 19019 6082
rect 10397 6024 10402 6080
rect 10458 6024 18958 6080
rect 19014 6024 19019 6080
rect 10397 6022 19019 6024
rect 10397 6019 10463 6022
rect 18953 6019 19019 6022
rect 9805 6016 10125 6017
rect 9805 5952 9813 6016
rect 9877 5952 9893 6016
rect 9957 5952 9973 6016
rect 10037 5952 10053 6016
rect 10117 5952 10125 6016
rect 9805 5951 10125 5952
rect 19138 6016 19458 6017
rect 19138 5952 19146 6016
rect 19210 5952 19226 6016
rect 19290 5952 19306 6016
rect 19370 5952 19386 6016
rect 19450 5952 19458 6016
rect 19138 5951 19458 5952
rect 22265 5946 22331 5949
rect 19646 5944 22331 5946
rect 19646 5888 22270 5944
rect 22326 5888 22331 5944
rect 19646 5886 22331 5888
rect 8189 5810 8255 5813
rect 19646 5810 19706 5886
rect 22265 5883 22331 5886
rect 8189 5808 19706 5810
rect 8189 5752 8194 5808
rect 8250 5752 19706 5808
rect 8189 5750 19706 5752
rect 20701 5810 20767 5813
rect 23185 5810 23251 5813
rect 20701 5808 23251 5810
rect 20701 5752 20706 5808
rect 20762 5752 23190 5808
rect 23246 5752 23251 5808
rect 20701 5750 23251 5752
rect 8189 5747 8255 5750
rect 20701 5747 20767 5750
rect 23185 5747 23251 5750
rect 7729 5674 7795 5677
rect 15457 5674 15523 5677
rect 16193 5674 16259 5677
rect 7729 5672 11840 5674
rect 7729 5616 7734 5672
rect 7790 5640 11840 5672
rect 11918 5640 14922 5674
rect 7790 5616 14922 5640
rect 7729 5614 14922 5616
rect 7729 5611 7795 5614
rect 11780 5580 11978 5614
rect 14862 5538 14922 5614
rect 15457 5672 16259 5674
rect 15457 5616 15462 5672
rect 15518 5616 16198 5672
rect 16254 5616 16259 5672
rect 15457 5614 16259 5616
rect 15457 5611 15523 5614
rect 16193 5611 16259 5614
rect 18953 5674 19019 5677
rect 20609 5674 20675 5677
rect 18953 5672 20675 5674
rect 18953 5616 18958 5672
rect 19014 5616 20614 5672
rect 20670 5616 20675 5672
rect 18953 5614 20675 5616
rect 18953 5611 19019 5614
rect 20609 5611 20675 5614
rect 24933 5674 24999 5677
rect 27048 5674 27528 5704
rect 24933 5672 27528 5674
rect 24933 5616 24938 5672
rect 24994 5616 27528 5672
rect 24933 5614 27528 5616
rect 24933 5611 24999 5614
rect 27048 5584 27528 5614
rect 14862 5478 16900 5538
rect 5138 5472 5458 5473
rect 5138 5408 5146 5472
rect 5210 5408 5226 5472
rect 5290 5408 5306 5472
rect 5370 5408 5386 5472
rect 5450 5408 5458 5472
rect 5138 5407 5458 5408
rect 14472 5472 14792 5473
rect 14472 5408 14480 5472
rect 14544 5408 14560 5472
rect 14624 5408 14640 5472
rect 14704 5408 14720 5472
rect 14784 5408 14792 5472
rect 14472 5407 14792 5408
rect 6441 5402 6507 5405
rect 10213 5402 10279 5405
rect 6441 5400 10279 5402
rect 6441 5344 6446 5400
rect 6502 5344 10218 5400
rect 10274 5344 10279 5400
rect 6441 5342 10279 5344
rect 6441 5339 6507 5342
rect 10213 5339 10279 5342
rect 6533 5266 6599 5269
rect 16840 5266 16900 5478
rect 23805 5472 24125 5473
rect 23805 5408 23813 5472
rect 23877 5408 23893 5472
rect 23957 5408 23973 5472
rect 24037 5408 24053 5472
rect 24117 5408 24125 5472
rect 23805 5407 24125 5408
rect 17021 5402 17087 5405
rect 23185 5402 23251 5405
rect 17021 5400 23251 5402
rect 17021 5344 17026 5400
rect 17082 5344 23190 5400
rect 23246 5344 23251 5400
rect 17021 5342 23251 5344
rect 17021 5339 17087 5342
rect 23185 5339 23251 5342
rect 25025 5266 25091 5269
rect 6533 5264 14692 5266
rect 6533 5208 6538 5264
rect 6594 5208 14692 5264
rect 6533 5206 14692 5208
rect 16840 5264 25091 5266
rect 16840 5208 25030 5264
rect 25086 5208 25091 5264
rect 16840 5206 25091 5208
rect 6533 5203 6599 5206
rect 8189 5130 8255 5133
rect 14632 5130 14692 5206
rect 25025 5203 25091 5206
rect 21897 5130 21963 5133
rect 8189 5128 14048 5130
rect 8189 5072 8194 5128
rect 8250 5072 14048 5128
rect 8189 5070 14048 5072
rect 14632 5128 21963 5130
rect 14632 5072 21902 5128
rect 21958 5072 21963 5128
rect 14632 5070 21963 5072
rect 8189 5067 8255 5070
rect 13988 4994 14048 5070
rect 21897 5067 21963 5070
rect 22030 5068 22036 5132
rect 22100 5130 22106 5132
rect 22173 5130 22239 5133
rect 22100 5128 22239 5130
rect 22100 5072 22178 5128
rect 22234 5072 22239 5128
rect 22100 5070 22239 5072
rect 22100 5068 22106 5070
rect 22173 5067 22239 5070
rect 23185 5130 23251 5133
rect 24841 5130 24907 5133
rect 23185 5128 24907 5130
rect 23185 5072 23190 5128
rect 23246 5072 24846 5128
rect 24902 5072 24907 5128
rect 23185 5070 24907 5072
rect 23185 5067 23251 5070
rect 24841 5067 24907 5070
rect 16837 4994 16903 4997
rect 13988 4992 16903 4994
rect 13988 4936 16842 4992
rect 16898 4936 16903 4992
rect 13988 4934 16903 4936
rect 16837 4931 16903 4934
rect 9805 4928 10125 4929
rect 9805 4864 9813 4928
rect 9877 4864 9893 4928
rect 9957 4864 9973 4928
rect 10037 4864 10053 4928
rect 10117 4864 10125 4928
rect 9805 4863 10125 4864
rect 19138 4928 19458 4929
rect 19138 4864 19146 4928
rect 19210 4864 19226 4928
rect 19290 4864 19306 4928
rect 19370 4864 19386 4928
rect 19450 4864 19458 4928
rect 19138 4863 19458 4864
rect 3405 4858 3471 4861
rect 9569 4858 9635 4861
rect 3405 4856 9635 4858
rect 3405 4800 3410 4856
rect 3466 4800 9574 4856
rect 9630 4800 9635 4856
rect 3405 4798 9635 4800
rect 3405 4795 3471 4798
rect 9569 4795 9635 4798
rect 10254 4796 10260 4860
rect 10324 4858 10330 4860
rect 14261 4858 14327 4861
rect 10324 4856 14327 4858
rect 10324 4800 14266 4856
rect 14322 4800 14327 4856
rect 10324 4798 14327 4800
rect 10324 4796 10330 4798
rect 14261 4795 14327 4798
rect 21345 4858 21411 4861
rect 23645 4858 23711 4861
rect 21345 4856 23711 4858
rect 21345 4800 21350 4856
rect 21406 4800 23650 4856
rect 23706 4800 23711 4856
rect 21345 4798 23711 4800
rect 21345 4795 21411 4798
rect 23645 4795 23711 4798
rect 9477 4722 9543 4725
rect 16837 4722 16903 4725
rect 23645 4722 23711 4725
rect 9477 4720 16762 4722
rect 9477 4664 9482 4720
rect 9538 4664 16762 4720
rect 9477 4662 16762 4664
rect 9477 4659 9543 4662
rect 4969 4586 5035 4589
rect 12421 4586 12487 4589
rect 16702 4586 16762 4662
rect 16837 4720 23711 4722
rect 16837 4664 16842 4720
rect 16898 4664 23650 4720
rect 23706 4664 23711 4720
rect 16837 4662 23711 4664
rect 16837 4659 16903 4662
rect 23645 4659 23711 4662
rect 22081 4586 22147 4589
rect 4969 4584 12487 4586
rect 4969 4528 4974 4584
rect 5030 4528 12426 4584
rect 12482 4528 12487 4584
rect 4969 4526 12487 4528
rect 4969 4523 5035 4526
rect 12421 4523 12487 4526
rect 14310 4526 14922 4586
rect 16702 4584 22147 4586
rect 16702 4528 22086 4584
rect 22142 4528 22147 4584
rect 16702 4526 22147 4528
rect 8097 4450 8163 4453
rect 14310 4450 14370 4526
rect 8097 4448 14370 4450
rect 8097 4392 8102 4448
rect 8158 4392 14370 4448
rect 8097 4390 14370 4392
rect 14862 4450 14922 4526
rect 22081 4523 22147 4526
rect 24933 4586 24999 4589
rect 27048 4586 27528 4616
rect 24933 4584 27528 4586
rect 24933 4528 24938 4584
rect 24994 4528 27528 4584
rect 24933 4526 27528 4528
rect 24933 4523 24999 4526
rect 27048 4496 27528 4526
rect 23001 4450 23067 4453
rect 14862 4448 23067 4450
rect 14862 4392 23006 4448
rect 23062 4392 23067 4448
rect 14862 4390 23067 4392
rect 8097 4387 8163 4390
rect 23001 4387 23067 4390
rect 5138 4384 5458 4385
rect 5138 4320 5146 4384
rect 5210 4320 5226 4384
rect 5290 4320 5306 4384
rect 5370 4320 5386 4384
rect 5450 4320 5458 4384
rect 5138 4319 5458 4320
rect 14472 4384 14792 4385
rect 14472 4320 14480 4384
rect 14544 4320 14560 4384
rect 14624 4320 14640 4384
rect 14704 4320 14720 4384
rect 14784 4320 14792 4384
rect 14472 4319 14792 4320
rect 23805 4384 24125 4385
rect 23805 4320 23813 4384
rect 23877 4320 23893 4384
rect 23957 4320 23973 4384
rect 24037 4320 24053 4384
rect 24117 4320 24125 4384
rect 23805 4319 24125 4320
rect 9109 4314 9175 4317
rect 13709 4314 13775 4317
rect 9109 4312 13775 4314
rect 9109 4256 9114 4312
rect 9170 4256 13714 4312
rect 13770 4256 13775 4312
rect 9109 4254 13775 4256
rect 9109 4251 9175 4254
rect 13709 4251 13775 4254
rect 21529 4314 21595 4317
rect 23553 4314 23619 4317
rect 21529 4312 23619 4314
rect 21529 4256 21534 4312
rect 21590 4256 23558 4312
rect 23614 4256 23619 4312
rect 21529 4254 23619 4256
rect 21529 4251 21595 4254
rect 23553 4251 23619 4254
rect 6533 4178 6599 4181
rect 9293 4178 9359 4181
rect 6533 4176 9359 4178
rect 6533 4120 6538 4176
rect 6594 4120 9298 4176
rect 9354 4120 9359 4176
rect 6533 4118 9359 4120
rect 6533 4115 6599 4118
rect 9293 4115 9359 4118
rect 9569 4178 9635 4181
rect 16101 4178 16167 4181
rect 9569 4176 16167 4178
rect 9569 4120 9574 4176
rect 9630 4120 16106 4176
rect 16162 4120 16167 4176
rect 9569 4118 16167 4120
rect 9569 4115 9635 4118
rect 16101 4115 16167 4118
rect 22725 4178 22791 4181
rect 25209 4178 25275 4181
rect 22725 4176 25275 4178
rect 22725 4120 22730 4176
rect 22786 4120 25214 4176
rect 25270 4120 25275 4176
rect 22725 4118 25275 4120
rect 22725 4115 22791 4118
rect 25209 4115 25275 4118
rect 3589 4042 3655 4045
rect 8465 4042 8531 4045
rect 3589 4040 8531 4042
rect 3589 3984 3594 4040
rect 3650 3984 8470 4040
rect 8526 3984 8531 4040
rect 3589 3982 8531 3984
rect 3589 3979 3655 3982
rect 8465 3979 8531 3982
rect 9017 4042 9083 4045
rect 12145 4042 12211 4045
rect 9017 4040 12211 4042
rect 9017 3984 9022 4040
rect 9078 3984 12150 4040
rect 12206 3984 12211 4040
rect 9017 3982 12211 3984
rect 9017 3979 9083 3982
rect 12145 3979 12211 3982
rect 17573 4042 17639 4045
rect 23277 4042 23343 4045
rect 17573 4040 23343 4042
rect 17573 3984 17578 4040
rect 17634 3984 23282 4040
rect 23338 3984 23343 4040
rect 17573 3982 23343 3984
rect 17573 3979 17639 3982
rect 23277 3979 23343 3982
rect 15733 3906 15799 3909
rect 15733 3904 16578 3906
rect 15733 3848 15738 3904
rect 15794 3848 16578 3904
rect 15733 3846 16578 3848
rect 15733 3843 15799 3846
rect 9805 3840 10125 3841
rect 9805 3776 9813 3840
rect 9877 3776 9893 3840
rect 9957 3776 9973 3840
rect 10037 3776 10053 3840
rect 10117 3776 10125 3840
rect 9805 3775 10125 3776
rect 1 3770 67 3773
rect 5705 3770 5771 3773
rect 1 3768 5771 3770
rect 1 3712 6 3768
rect 62 3712 5710 3768
rect 5766 3712 5771 3768
rect 1 3710 5771 3712
rect 1 3707 67 3710
rect 5705 3707 5771 3710
rect 6073 3770 6139 3773
rect 6206 3770 6212 3772
rect 6073 3768 6212 3770
rect 6073 3712 6078 3768
rect 6134 3712 6212 3768
rect 6073 3710 6212 3712
rect 6073 3707 6139 3710
rect 6206 3708 6212 3710
rect 6276 3708 6282 3772
rect 11961 3770 12027 3773
rect 11961 3768 16394 3770
rect 11961 3712 11966 3768
rect 12022 3712 16394 3768
rect 11961 3710 16394 3712
rect 11961 3707 12027 3710
rect 3957 3634 4023 3637
rect 16193 3634 16259 3637
rect 3957 3632 16259 3634
rect 3957 3576 3962 3632
rect 4018 3576 16198 3632
rect 16254 3576 16259 3632
rect 3957 3574 16259 3576
rect 3957 3571 4023 3574
rect 16193 3571 16259 3574
rect 4601 3498 4667 3501
rect 13249 3498 13315 3501
rect 14813 3498 14879 3501
rect 4601 3496 14879 3498
rect 4601 3440 4606 3496
rect 4662 3440 13254 3496
rect 13310 3440 14818 3496
rect 14874 3440 14879 3496
rect 4601 3438 14879 3440
rect 4601 3435 4667 3438
rect 13249 3435 13315 3438
rect 14813 3435 14879 3438
rect 6901 3362 6967 3365
rect 13157 3362 13223 3365
rect 13801 3362 13867 3365
rect 6901 3360 13867 3362
rect 6901 3304 6906 3360
rect 6962 3304 13162 3360
rect 13218 3304 13806 3360
rect 13862 3304 13867 3360
rect 6901 3302 13867 3304
rect 16334 3362 16394 3710
rect 16518 3634 16578 3846
rect 19138 3840 19458 3841
rect 19138 3776 19146 3840
rect 19210 3776 19226 3840
rect 19290 3776 19306 3840
rect 19370 3776 19386 3840
rect 19450 3776 19458 3840
rect 19138 3775 19458 3776
rect 22357 3634 22423 3637
rect 16518 3632 22423 3634
rect 16518 3576 22362 3632
rect 22418 3576 22423 3632
rect 16518 3574 22423 3576
rect 22357 3571 22423 3574
rect 24749 3498 24815 3501
rect 23648 3496 24815 3498
rect 23648 3440 24754 3496
rect 24810 3440 24815 3496
rect 23648 3438 24815 3440
rect 23648 3362 23708 3438
rect 24749 3435 24815 3438
rect 24933 3498 24999 3501
rect 27048 3498 27528 3528
rect 24933 3496 27528 3498
rect 24933 3440 24938 3496
rect 24994 3440 27528 3496
rect 24933 3438 27528 3440
rect 24933 3435 24999 3438
rect 27048 3408 27528 3438
rect 16334 3302 23708 3362
rect 6901 3299 6967 3302
rect 13157 3299 13223 3302
rect 13801 3299 13867 3302
rect 5138 3296 5458 3297
rect 5138 3232 5146 3296
rect 5210 3232 5226 3296
rect 5290 3232 5306 3296
rect 5370 3232 5386 3296
rect 5450 3232 5458 3296
rect 5138 3231 5458 3232
rect 14472 3296 14792 3297
rect 14472 3232 14480 3296
rect 14544 3232 14560 3296
rect 14624 3232 14640 3296
rect 14704 3232 14720 3296
rect 14784 3232 14792 3296
rect 14472 3231 14792 3232
rect 23805 3296 24125 3297
rect 23805 3232 23813 3296
rect 23877 3232 23893 3296
rect 23957 3232 23973 3296
rect 24037 3232 24053 3296
rect 24117 3232 24125 3296
rect 23805 3231 24125 3232
rect 5797 3226 5863 3229
rect 12329 3226 12395 3229
rect 5797 3224 12395 3226
rect 5797 3168 5802 3224
rect 5858 3168 12334 3224
rect 12390 3168 12395 3224
rect 5797 3166 12395 3168
rect 5797 3163 5863 3166
rect 12329 3163 12395 3166
rect 15273 3226 15339 3229
rect 23093 3226 23159 3229
rect 15273 3224 23159 3226
rect 15273 3168 15278 3224
rect 15334 3168 23098 3224
rect 23154 3168 23159 3224
rect 15273 3166 23159 3168
rect 15273 3163 15339 3166
rect 23093 3163 23159 3166
rect 4877 3090 4943 3093
rect 7678 3090 7684 3092
rect 4877 3088 7684 3090
rect 4877 3032 4882 3088
rect 4938 3032 7684 3088
rect 4877 3030 7684 3032
rect 4877 3027 4943 3030
rect 7678 3028 7684 3030
rect 7748 3028 7754 3092
rect 8833 3090 8899 3093
rect 13433 3090 13499 3093
rect 8833 3088 13499 3090
rect 8833 3032 8838 3088
rect 8894 3032 13438 3088
rect 13494 3032 13499 3088
rect 8833 3030 13499 3032
rect 8833 3027 8899 3030
rect 13433 3027 13499 3030
rect 16009 3090 16075 3093
rect 17665 3090 17731 3093
rect 16009 3088 17731 3090
rect 16009 3032 16014 3088
rect 16070 3032 17670 3088
rect 17726 3032 17731 3088
rect 16009 3030 17731 3032
rect 16009 3027 16075 3030
rect 17665 3027 17731 3030
rect 1013 2954 1079 2957
rect 4233 2954 4299 2957
rect 1013 2952 4299 2954
rect 1013 2896 1018 2952
rect 1074 2896 4238 2952
rect 4294 2896 4299 2952
rect 1013 2894 4299 2896
rect 1013 2891 1079 2894
rect 4233 2891 4299 2894
rect 7177 2954 7243 2957
rect 14353 2954 14419 2957
rect 7177 2952 14419 2954
rect 7177 2896 7182 2952
rect 7238 2896 14358 2952
rect 14414 2896 14419 2952
rect 7177 2894 14419 2896
rect 7177 2891 7243 2894
rect 14353 2891 14419 2894
rect 18677 2954 18743 2957
rect 23001 2954 23067 2957
rect 18677 2952 23067 2954
rect 18677 2896 18682 2952
rect 18738 2896 23006 2952
rect 23062 2896 23067 2952
rect 18677 2894 23067 2896
rect 18677 2891 18743 2894
rect 23001 2891 23067 2894
rect 2025 2818 2091 2821
rect 4325 2818 4391 2821
rect 2025 2816 4391 2818
rect 2025 2760 2030 2816
rect 2086 2760 4330 2816
rect 4386 2760 4391 2816
rect 2025 2758 4391 2760
rect 2025 2755 2091 2758
rect 4325 2755 4391 2758
rect 5889 2818 5955 2821
rect 7177 2818 7243 2821
rect 5889 2816 7243 2818
rect 5889 2760 5894 2816
rect 5950 2760 7182 2816
rect 7238 2760 7243 2816
rect 5889 2758 7243 2760
rect 5889 2755 5955 2758
rect 7177 2755 7243 2758
rect 7729 2818 7795 2821
rect 9293 2818 9359 2821
rect 7729 2816 9359 2818
rect 7729 2760 7734 2816
rect 7790 2760 9298 2816
rect 9354 2760 9359 2816
rect 7729 2758 9359 2760
rect 7729 2755 7795 2758
rect 9293 2755 9359 2758
rect 10397 2818 10463 2821
rect 12237 2818 12303 2821
rect 10397 2816 12303 2818
rect 10397 2760 10402 2816
rect 10458 2760 12242 2816
rect 12298 2760 12303 2816
rect 10397 2758 12303 2760
rect 10397 2755 10463 2758
rect 12237 2755 12303 2758
rect 12421 2818 12487 2821
rect 14813 2818 14879 2821
rect 12421 2816 14879 2818
rect 12421 2760 12426 2816
rect 12482 2760 14818 2816
rect 14874 2760 14879 2816
rect 12421 2758 14879 2760
rect 12421 2755 12487 2758
rect 14813 2755 14879 2758
rect 9805 2752 10125 2753
rect 9805 2688 9813 2752
rect 9877 2688 9893 2752
rect 9957 2688 9973 2752
rect 10037 2688 10053 2752
rect 10117 2688 10125 2752
rect 9805 2687 10125 2688
rect 19138 2752 19458 2753
rect 19138 2688 19146 2752
rect 19210 2688 19226 2752
rect 19290 2688 19306 2752
rect 19370 2688 19386 2752
rect 19450 2688 19458 2752
rect 19138 2687 19458 2688
rect 4509 2682 4575 2685
rect 9385 2682 9451 2685
rect 4509 2680 9451 2682
rect 4509 2624 4514 2680
rect 4570 2624 9390 2680
rect 9446 2624 9451 2680
rect 4509 2622 9451 2624
rect 4509 2619 4575 2622
rect 9385 2619 9451 2622
rect 6717 2546 6783 2549
rect 17481 2546 17547 2549
rect 6717 2544 17547 2546
rect 6717 2488 6722 2544
rect 6778 2488 17486 2544
rect 17542 2488 17547 2544
rect 6717 2486 17547 2488
rect 6717 2483 6783 2486
rect 17481 2483 17547 2486
rect 23093 2546 23159 2549
rect 27048 2546 27528 2576
rect 23093 2544 27528 2546
rect 23093 2488 23098 2544
rect 23154 2488 27528 2544
rect 23093 2486 27528 2488
rect 23093 2483 23159 2486
rect 27048 2456 27528 2486
rect 5337 2410 5403 2413
rect 11501 2410 11567 2413
rect 22265 2412 22331 2413
rect 5337 2408 11567 2410
rect 5337 2352 5342 2408
rect 5398 2352 11506 2408
rect 11562 2352 11567 2408
rect 5337 2350 11567 2352
rect 5337 2347 5403 2350
rect 11501 2347 11567 2350
rect 22214 2348 22220 2412
rect 22284 2410 22331 2412
rect 22284 2408 22376 2410
rect 22326 2352 22376 2408
rect 22284 2350 22376 2352
rect 22284 2348 22331 2350
rect 22265 2347 22331 2348
rect 8741 2274 8807 2277
rect 11317 2274 11383 2277
rect 8741 2272 11383 2274
rect 8741 2216 8746 2272
rect 8802 2216 11322 2272
rect 11378 2216 11383 2272
rect 8741 2214 11383 2216
rect 8741 2211 8807 2214
rect 11317 2211 11383 2214
rect 5138 2208 5458 2209
rect 5138 2144 5146 2208
rect 5210 2144 5226 2208
rect 5290 2144 5306 2208
rect 5370 2144 5386 2208
rect 5450 2144 5458 2208
rect 5138 2143 5458 2144
rect 14472 2208 14792 2209
rect 14472 2144 14480 2208
rect 14544 2144 14560 2208
rect 14624 2144 14640 2208
rect 14704 2144 14720 2208
rect 14784 2144 14792 2208
rect 14472 2143 14792 2144
rect 23805 2208 24125 2209
rect 23805 2144 23813 2208
rect 23877 2144 23893 2208
rect 23957 2144 23973 2208
rect 24037 2144 24053 2208
rect 24117 2144 24125 2208
rect 23805 2143 24125 2144
rect 3037 2002 3103 2005
rect 15457 2002 15523 2005
rect 3037 2000 15523 2002
rect 3037 1944 3042 2000
rect 3098 1944 15462 2000
rect 15518 1944 15523 2000
rect 3037 1942 15523 1944
rect 3037 1939 3103 1942
rect 15457 1939 15523 1942
rect 5797 1866 5863 1869
rect 13801 1866 13867 1869
rect 5797 1864 13867 1866
rect 5797 1808 5802 1864
rect 5858 1808 13806 1864
rect 13862 1808 13867 1864
rect 5797 1806 13867 1808
rect 5797 1803 5863 1806
rect 13801 1803 13867 1806
rect 13985 1866 14051 1869
rect 20701 1866 20767 1869
rect 13985 1864 20767 1866
rect 13985 1808 13990 1864
rect 14046 1808 20706 1864
rect 20762 1808 20767 1864
rect 13985 1806 20767 1808
rect 13985 1803 14051 1806
rect 20701 1803 20767 1806
rect 2117 1732 2183 1733
rect 2117 1730 2164 1732
rect 2072 1728 2164 1730
rect 2072 1672 2122 1728
rect 2072 1670 2164 1672
rect 2117 1668 2164 1670
rect 2228 1668 2234 1732
rect 3221 1730 3287 1733
rect 16653 1730 16719 1733
rect 26865 1732 26931 1733
rect 26814 1730 26820 1732
rect 3221 1728 16719 1730
rect 3221 1672 3226 1728
rect 3282 1672 16658 1728
rect 16714 1672 16719 1728
rect 3221 1670 16719 1672
rect 26774 1670 26820 1730
rect 26884 1728 26931 1732
rect 26926 1672 26931 1728
rect 2117 1667 2183 1668
rect 3221 1667 3287 1670
rect 16653 1667 16719 1670
rect 26814 1668 26820 1670
rect 26884 1668 26931 1672
rect 26865 1667 26931 1668
rect 7545 1594 7611 1597
rect 18493 1594 18559 1597
rect 7545 1592 18559 1594
rect 7545 1536 7550 1592
rect 7606 1536 18498 1592
rect 18554 1536 18559 1592
rect 7545 1534 18559 1536
rect 7545 1531 7611 1534
rect 18493 1531 18559 1534
rect 2853 1458 2919 1461
rect 17573 1458 17639 1461
rect 2853 1456 17639 1458
rect 2853 1400 2858 1456
rect 2914 1400 17578 1456
rect 17634 1400 17639 1456
rect 2853 1398 17639 1400
rect 2853 1395 2919 1398
rect 17573 1395 17639 1398
rect 19597 1458 19663 1461
rect 22449 1458 22515 1461
rect 19597 1456 22515 1458
rect 19597 1400 19602 1456
rect 19658 1400 22454 1456
rect 22510 1400 22515 1456
rect 19597 1398 22515 1400
rect 19597 1395 19663 1398
rect 22449 1395 22515 1398
rect 23553 1458 23619 1461
rect 27048 1458 27528 1488
rect 23553 1456 27528 1458
rect 23553 1400 23558 1456
rect 23614 1400 27528 1456
rect 23553 1398 27528 1400
rect 23553 1395 23619 1398
rect 27048 1368 27528 1398
rect 8925 1322 8991 1325
rect 23369 1322 23435 1325
rect 8925 1320 23435 1322
rect 8925 1264 8930 1320
rect 8986 1264 23374 1320
rect 23430 1264 23435 1320
rect 8925 1262 23435 1264
rect 8925 1259 8991 1262
rect 23369 1259 23435 1262
rect 9109 1186 9175 1189
rect 23185 1186 23251 1189
rect 9109 1184 23251 1186
rect 9109 1128 9114 1184
rect 9170 1128 23190 1184
rect 23246 1128 23251 1184
rect 9109 1126 23251 1128
rect 9109 1123 9175 1126
rect 23185 1123 23251 1126
rect 5613 1050 5679 1053
rect 19413 1050 19479 1053
rect 5613 1048 19479 1050
rect 5613 992 5618 1048
rect 5674 992 19418 1048
rect 19474 992 19479 1048
rect 5613 990 19479 992
rect 5613 987 5679 990
rect 19413 987 19479 990
rect 7637 914 7703 917
rect 20057 914 20123 917
rect 7637 912 20123 914
rect 7637 856 7642 912
rect 7698 856 20062 912
rect 20118 856 20123 912
rect 7637 854 20123 856
rect 7637 851 7703 854
rect 20057 851 20123 854
rect 25117 506 25183 509
rect 27048 506 27528 536
rect 25117 504 27528 506
rect 25117 448 25122 504
rect 25178 448 27528 504
rect 25117 446 27528 448
rect 25117 443 25183 446
rect 27048 416 27528 446
<< via3 >>
rect 9813 25596 9877 25600
rect 9813 25540 9817 25596
rect 9817 25540 9873 25596
rect 9873 25540 9877 25596
rect 9813 25536 9877 25540
rect 9893 25596 9957 25600
rect 9893 25540 9897 25596
rect 9897 25540 9953 25596
rect 9953 25540 9957 25596
rect 9893 25536 9957 25540
rect 9973 25596 10037 25600
rect 9973 25540 9977 25596
rect 9977 25540 10033 25596
rect 10033 25540 10037 25596
rect 9973 25536 10037 25540
rect 10053 25596 10117 25600
rect 10053 25540 10057 25596
rect 10057 25540 10113 25596
rect 10113 25540 10117 25596
rect 10053 25536 10117 25540
rect 19146 25596 19210 25600
rect 19146 25540 19150 25596
rect 19150 25540 19206 25596
rect 19206 25540 19210 25596
rect 19146 25536 19210 25540
rect 19226 25596 19290 25600
rect 19226 25540 19230 25596
rect 19230 25540 19286 25596
rect 19286 25540 19290 25596
rect 19226 25536 19290 25540
rect 19306 25596 19370 25600
rect 19306 25540 19310 25596
rect 19310 25540 19366 25596
rect 19366 25540 19370 25596
rect 19306 25536 19370 25540
rect 19386 25596 19450 25600
rect 19386 25540 19390 25596
rect 19390 25540 19446 25596
rect 19446 25540 19450 25596
rect 19386 25536 19450 25540
rect 5146 25052 5210 25056
rect 5146 24996 5150 25052
rect 5150 24996 5206 25052
rect 5206 24996 5210 25052
rect 5146 24992 5210 24996
rect 5226 25052 5290 25056
rect 5226 24996 5230 25052
rect 5230 24996 5286 25052
rect 5286 24996 5290 25052
rect 5226 24992 5290 24996
rect 5306 25052 5370 25056
rect 5306 24996 5310 25052
rect 5310 24996 5366 25052
rect 5366 24996 5370 25052
rect 5306 24992 5370 24996
rect 5386 25052 5450 25056
rect 5386 24996 5390 25052
rect 5390 24996 5446 25052
rect 5446 24996 5450 25052
rect 5386 24992 5450 24996
rect 14480 25052 14544 25056
rect 14480 24996 14484 25052
rect 14484 24996 14540 25052
rect 14540 24996 14544 25052
rect 14480 24992 14544 24996
rect 14560 25052 14624 25056
rect 14560 24996 14564 25052
rect 14564 24996 14620 25052
rect 14620 24996 14624 25052
rect 14560 24992 14624 24996
rect 14640 25052 14704 25056
rect 14640 24996 14644 25052
rect 14644 24996 14700 25052
rect 14700 24996 14704 25052
rect 14640 24992 14704 24996
rect 14720 25052 14784 25056
rect 14720 24996 14724 25052
rect 14724 24996 14780 25052
rect 14780 24996 14784 25052
rect 14720 24992 14784 24996
rect 23813 25052 23877 25056
rect 23813 24996 23817 25052
rect 23817 24996 23873 25052
rect 23873 24996 23877 25052
rect 23813 24992 23877 24996
rect 23893 25052 23957 25056
rect 23893 24996 23897 25052
rect 23897 24996 23953 25052
rect 23953 24996 23957 25052
rect 23893 24992 23957 24996
rect 23973 25052 24037 25056
rect 23973 24996 23977 25052
rect 23977 24996 24033 25052
rect 24033 24996 24037 25052
rect 23973 24992 24037 24996
rect 24053 25052 24117 25056
rect 24053 24996 24057 25052
rect 24057 24996 24113 25052
rect 24113 24996 24117 25052
rect 24053 24992 24117 24996
rect 9813 24508 9877 24512
rect 9813 24452 9817 24508
rect 9817 24452 9873 24508
rect 9873 24452 9877 24508
rect 9813 24448 9877 24452
rect 9893 24508 9957 24512
rect 9893 24452 9897 24508
rect 9897 24452 9953 24508
rect 9953 24452 9957 24508
rect 9893 24448 9957 24452
rect 9973 24508 10037 24512
rect 9973 24452 9977 24508
rect 9977 24452 10033 24508
rect 10033 24452 10037 24508
rect 9973 24448 10037 24452
rect 10053 24508 10117 24512
rect 10053 24452 10057 24508
rect 10057 24452 10113 24508
rect 10113 24452 10117 24508
rect 10053 24448 10117 24452
rect 19146 24508 19210 24512
rect 19146 24452 19150 24508
rect 19150 24452 19206 24508
rect 19206 24452 19210 24508
rect 19146 24448 19210 24452
rect 19226 24508 19290 24512
rect 19226 24452 19230 24508
rect 19230 24452 19286 24508
rect 19286 24452 19290 24508
rect 19226 24448 19290 24452
rect 19306 24508 19370 24512
rect 19306 24452 19310 24508
rect 19310 24452 19366 24508
rect 19366 24452 19370 24508
rect 19306 24448 19370 24452
rect 19386 24508 19450 24512
rect 19386 24452 19390 24508
rect 19390 24452 19446 24508
rect 19446 24452 19450 24508
rect 19386 24448 19450 24452
rect 5146 23964 5210 23968
rect 5146 23908 5150 23964
rect 5150 23908 5206 23964
rect 5206 23908 5210 23964
rect 5146 23904 5210 23908
rect 5226 23964 5290 23968
rect 5226 23908 5230 23964
rect 5230 23908 5286 23964
rect 5286 23908 5290 23964
rect 5226 23904 5290 23908
rect 5306 23964 5370 23968
rect 5306 23908 5310 23964
rect 5310 23908 5366 23964
rect 5366 23908 5370 23964
rect 5306 23904 5370 23908
rect 5386 23964 5450 23968
rect 5386 23908 5390 23964
rect 5390 23908 5446 23964
rect 5446 23908 5450 23964
rect 5386 23904 5450 23908
rect 14480 23964 14544 23968
rect 14480 23908 14484 23964
rect 14484 23908 14540 23964
rect 14540 23908 14544 23964
rect 14480 23904 14544 23908
rect 14560 23964 14624 23968
rect 14560 23908 14564 23964
rect 14564 23908 14620 23964
rect 14620 23908 14624 23964
rect 14560 23904 14624 23908
rect 14640 23964 14704 23968
rect 14640 23908 14644 23964
rect 14644 23908 14700 23964
rect 14700 23908 14704 23964
rect 14640 23904 14704 23908
rect 14720 23964 14784 23968
rect 14720 23908 14724 23964
rect 14724 23908 14780 23964
rect 14780 23908 14784 23964
rect 14720 23904 14784 23908
rect 23813 23964 23877 23968
rect 23813 23908 23817 23964
rect 23817 23908 23873 23964
rect 23873 23908 23877 23964
rect 23813 23904 23877 23908
rect 23893 23964 23957 23968
rect 23893 23908 23897 23964
rect 23897 23908 23953 23964
rect 23953 23908 23957 23964
rect 23893 23904 23957 23908
rect 23973 23964 24037 23968
rect 23973 23908 23977 23964
rect 23977 23908 24033 23964
rect 24033 23908 24037 23964
rect 23973 23904 24037 23908
rect 24053 23964 24117 23968
rect 24053 23908 24057 23964
rect 24057 23908 24113 23964
rect 24113 23908 24117 23964
rect 24053 23904 24117 23908
rect 9813 23420 9877 23424
rect 9813 23364 9817 23420
rect 9817 23364 9873 23420
rect 9873 23364 9877 23420
rect 9813 23360 9877 23364
rect 9893 23420 9957 23424
rect 9893 23364 9897 23420
rect 9897 23364 9953 23420
rect 9953 23364 9957 23420
rect 9893 23360 9957 23364
rect 9973 23420 10037 23424
rect 9973 23364 9977 23420
rect 9977 23364 10033 23420
rect 10033 23364 10037 23420
rect 9973 23360 10037 23364
rect 10053 23420 10117 23424
rect 10053 23364 10057 23420
rect 10057 23364 10113 23420
rect 10113 23364 10117 23420
rect 10053 23360 10117 23364
rect 19146 23420 19210 23424
rect 19146 23364 19150 23420
rect 19150 23364 19206 23420
rect 19206 23364 19210 23420
rect 19146 23360 19210 23364
rect 19226 23420 19290 23424
rect 19226 23364 19230 23420
rect 19230 23364 19286 23420
rect 19286 23364 19290 23420
rect 19226 23360 19290 23364
rect 19306 23420 19370 23424
rect 19306 23364 19310 23420
rect 19310 23364 19366 23420
rect 19366 23364 19370 23420
rect 19306 23360 19370 23364
rect 19386 23420 19450 23424
rect 19386 23364 19390 23420
rect 19390 23364 19446 23420
rect 19446 23364 19450 23420
rect 19386 23360 19450 23364
rect 5146 22876 5210 22880
rect 5146 22820 5150 22876
rect 5150 22820 5206 22876
rect 5206 22820 5210 22876
rect 5146 22816 5210 22820
rect 5226 22876 5290 22880
rect 5226 22820 5230 22876
rect 5230 22820 5286 22876
rect 5286 22820 5290 22876
rect 5226 22816 5290 22820
rect 5306 22876 5370 22880
rect 5306 22820 5310 22876
rect 5310 22820 5366 22876
rect 5366 22820 5370 22876
rect 5306 22816 5370 22820
rect 5386 22876 5450 22880
rect 5386 22820 5390 22876
rect 5390 22820 5446 22876
rect 5446 22820 5450 22876
rect 5386 22816 5450 22820
rect 14480 22876 14544 22880
rect 14480 22820 14484 22876
rect 14484 22820 14540 22876
rect 14540 22820 14544 22876
rect 14480 22816 14544 22820
rect 14560 22876 14624 22880
rect 14560 22820 14564 22876
rect 14564 22820 14620 22876
rect 14620 22820 14624 22876
rect 14560 22816 14624 22820
rect 14640 22876 14704 22880
rect 14640 22820 14644 22876
rect 14644 22820 14700 22876
rect 14700 22820 14704 22876
rect 14640 22816 14704 22820
rect 14720 22876 14784 22880
rect 14720 22820 14724 22876
rect 14724 22820 14780 22876
rect 14780 22820 14784 22876
rect 14720 22816 14784 22820
rect 23813 22876 23877 22880
rect 23813 22820 23817 22876
rect 23817 22820 23873 22876
rect 23873 22820 23877 22876
rect 23813 22816 23877 22820
rect 23893 22876 23957 22880
rect 23893 22820 23897 22876
rect 23897 22820 23953 22876
rect 23953 22820 23957 22876
rect 23893 22816 23957 22820
rect 23973 22876 24037 22880
rect 23973 22820 23977 22876
rect 23977 22820 24033 22876
rect 24033 22820 24037 22876
rect 23973 22816 24037 22820
rect 24053 22876 24117 22880
rect 24053 22820 24057 22876
rect 24057 22820 24113 22876
rect 24113 22820 24117 22876
rect 24053 22816 24117 22820
rect 9813 22332 9877 22336
rect 9813 22276 9817 22332
rect 9817 22276 9873 22332
rect 9873 22276 9877 22332
rect 9813 22272 9877 22276
rect 9893 22332 9957 22336
rect 9893 22276 9897 22332
rect 9897 22276 9953 22332
rect 9953 22276 9957 22332
rect 9893 22272 9957 22276
rect 9973 22332 10037 22336
rect 9973 22276 9977 22332
rect 9977 22276 10033 22332
rect 10033 22276 10037 22332
rect 9973 22272 10037 22276
rect 10053 22332 10117 22336
rect 10053 22276 10057 22332
rect 10057 22276 10113 22332
rect 10113 22276 10117 22332
rect 10053 22272 10117 22276
rect 19146 22332 19210 22336
rect 19146 22276 19150 22332
rect 19150 22276 19206 22332
rect 19206 22276 19210 22332
rect 19146 22272 19210 22276
rect 19226 22332 19290 22336
rect 19226 22276 19230 22332
rect 19230 22276 19286 22332
rect 19286 22276 19290 22332
rect 19226 22272 19290 22276
rect 19306 22332 19370 22336
rect 19306 22276 19310 22332
rect 19310 22276 19366 22332
rect 19366 22276 19370 22332
rect 19306 22272 19370 22276
rect 19386 22332 19450 22336
rect 19386 22276 19390 22332
rect 19390 22276 19446 22332
rect 19446 22276 19450 22332
rect 19386 22272 19450 22276
rect 5146 21788 5210 21792
rect 5146 21732 5150 21788
rect 5150 21732 5206 21788
rect 5206 21732 5210 21788
rect 5146 21728 5210 21732
rect 5226 21788 5290 21792
rect 5226 21732 5230 21788
rect 5230 21732 5286 21788
rect 5286 21732 5290 21788
rect 5226 21728 5290 21732
rect 5306 21788 5370 21792
rect 5306 21732 5310 21788
rect 5310 21732 5366 21788
rect 5366 21732 5370 21788
rect 5306 21728 5370 21732
rect 5386 21788 5450 21792
rect 5386 21732 5390 21788
rect 5390 21732 5446 21788
rect 5446 21732 5450 21788
rect 5386 21728 5450 21732
rect 14480 21788 14544 21792
rect 14480 21732 14484 21788
rect 14484 21732 14540 21788
rect 14540 21732 14544 21788
rect 14480 21728 14544 21732
rect 14560 21788 14624 21792
rect 14560 21732 14564 21788
rect 14564 21732 14620 21788
rect 14620 21732 14624 21788
rect 14560 21728 14624 21732
rect 14640 21788 14704 21792
rect 14640 21732 14644 21788
rect 14644 21732 14700 21788
rect 14700 21732 14704 21788
rect 14640 21728 14704 21732
rect 14720 21788 14784 21792
rect 14720 21732 14724 21788
rect 14724 21732 14780 21788
rect 14780 21732 14784 21788
rect 14720 21728 14784 21732
rect 23813 21788 23877 21792
rect 23813 21732 23817 21788
rect 23817 21732 23873 21788
rect 23873 21732 23877 21788
rect 23813 21728 23877 21732
rect 23893 21788 23957 21792
rect 23893 21732 23897 21788
rect 23897 21732 23953 21788
rect 23953 21732 23957 21788
rect 23893 21728 23957 21732
rect 23973 21788 24037 21792
rect 23973 21732 23977 21788
rect 23977 21732 24033 21788
rect 24033 21732 24037 21788
rect 23973 21728 24037 21732
rect 24053 21788 24117 21792
rect 24053 21732 24057 21788
rect 24057 21732 24113 21788
rect 24113 21732 24117 21788
rect 24053 21728 24117 21732
rect 9813 21244 9877 21248
rect 9813 21188 9817 21244
rect 9817 21188 9873 21244
rect 9873 21188 9877 21244
rect 9813 21184 9877 21188
rect 9893 21244 9957 21248
rect 9893 21188 9897 21244
rect 9897 21188 9953 21244
rect 9953 21188 9957 21244
rect 9893 21184 9957 21188
rect 9973 21244 10037 21248
rect 9973 21188 9977 21244
rect 9977 21188 10033 21244
rect 10033 21188 10037 21244
rect 9973 21184 10037 21188
rect 10053 21244 10117 21248
rect 10053 21188 10057 21244
rect 10057 21188 10113 21244
rect 10113 21188 10117 21244
rect 10053 21184 10117 21188
rect 19146 21244 19210 21248
rect 19146 21188 19150 21244
rect 19150 21188 19206 21244
rect 19206 21188 19210 21244
rect 19146 21184 19210 21188
rect 19226 21244 19290 21248
rect 19226 21188 19230 21244
rect 19230 21188 19286 21244
rect 19286 21188 19290 21244
rect 19226 21184 19290 21188
rect 19306 21244 19370 21248
rect 19306 21188 19310 21244
rect 19310 21188 19366 21244
rect 19366 21188 19370 21244
rect 19306 21184 19370 21188
rect 19386 21244 19450 21248
rect 19386 21188 19390 21244
rect 19390 21188 19446 21244
rect 19446 21188 19450 21244
rect 19386 21184 19450 21188
rect 5146 20700 5210 20704
rect 5146 20644 5150 20700
rect 5150 20644 5206 20700
rect 5206 20644 5210 20700
rect 5146 20640 5210 20644
rect 5226 20700 5290 20704
rect 5226 20644 5230 20700
rect 5230 20644 5286 20700
rect 5286 20644 5290 20700
rect 5226 20640 5290 20644
rect 5306 20700 5370 20704
rect 5306 20644 5310 20700
rect 5310 20644 5366 20700
rect 5366 20644 5370 20700
rect 5306 20640 5370 20644
rect 5386 20700 5450 20704
rect 5386 20644 5390 20700
rect 5390 20644 5446 20700
rect 5446 20644 5450 20700
rect 5386 20640 5450 20644
rect 14480 20700 14544 20704
rect 14480 20644 14484 20700
rect 14484 20644 14540 20700
rect 14540 20644 14544 20700
rect 14480 20640 14544 20644
rect 14560 20700 14624 20704
rect 14560 20644 14564 20700
rect 14564 20644 14620 20700
rect 14620 20644 14624 20700
rect 14560 20640 14624 20644
rect 14640 20700 14704 20704
rect 14640 20644 14644 20700
rect 14644 20644 14700 20700
rect 14700 20644 14704 20700
rect 14640 20640 14704 20644
rect 14720 20700 14784 20704
rect 14720 20644 14724 20700
rect 14724 20644 14780 20700
rect 14780 20644 14784 20700
rect 14720 20640 14784 20644
rect 23813 20700 23877 20704
rect 23813 20644 23817 20700
rect 23817 20644 23873 20700
rect 23873 20644 23877 20700
rect 23813 20640 23877 20644
rect 23893 20700 23957 20704
rect 23893 20644 23897 20700
rect 23897 20644 23953 20700
rect 23953 20644 23957 20700
rect 23893 20640 23957 20644
rect 23973 20700 24037 20704
rect 23973 20644 23977 20700
rect 23977 20644 24033 20700
rect 24033 20644 24037 20700
rect 23973 20640 24037 20644
rect 24053 20700 24117 20704
rect 24053 20644 24057 20700
rect 24057 20644 24113 20700
rect 24113 20644 24117 20700
rect 24053 20640 24117 20644
rect 9813 20156 9877 20160
rect 9813 20100 9817 20156
rect 9817 20100 9873 20156
rect 9873 20100 9877 20156
rect 9813 20096 9877 20100
rect 9893 20156 9957 20160
rect 9893 20100 9897 20156
rect 9897 20100 9953 20156
rect 9953 20100 9957 20156
rect 9893 20096 9957 20100
rect 9973 20156 10037 20160
rect 9973 20100 9977 20156
rect 9977 20100 10033 20156
rect 10033 20100 10037 20156
rect 9973 20096 10037 20100
rect 10053 20156 10117 20160
rect 10053 20100 10057 20156
rect 10057 20100 10113 20156
rect 10113 20100 10117 20156
rect 10053 20096 10117 20100
rect 19146 20156 19210 20160
rect 19146 20100 19150 20156
rect 19150 20100 19206 20156
rect 19206 20100 19210 20156
rect 19146 20096 19210 20100
rect 19226 20156 19290 20160
rect 19226 20100 19230 20156
rect 19230 20100 19286 20156
rect 19286 20100 19290 20156
rect 19226 20096 19290 20100
rect 19306 20156 19370 20160
rect 19306 20100 19310 20156
rect 19310 20100 19366 20156
rect 19366 20100 19370 20156
rect 19306 20096 19370 20100
rect 19386 20156 19450 20160
rect 19386 20100 19390 20156
rect 19390 20100 19446 20156
rect 19446 20100 19450 20156
rect 19386 20096 19450 20100
rect 5146 19612 5210 19616
rect 5146 19556 5150 19612
rect 5150 19556 5206 19612
rect 5206 19556 5210 19612
rect 5146 19552 5210 19556
rect 5226 19612 5290 19616
rect 5226 19556 5230 19612
rect 5230 19556 5286 19612
rect 5286 19556 5290 19612
rect 5226 19552 5290 19556
rect 5306 19612 5370 19616
rect 5306 19556 5310 19612
rect 5310 19556 5366 19612
rect 5366 19556 5370 19612
rect 5306 19552 5370 19556
rect 5386 19612 5450 19616
rect 5386 19556 5390 19612
rect 5390 19556 5446 19612
rect 5446 19556 5450 19612
rect 5386 19552 5450 19556
rect 14480 19612 14544 19616
rect 14480 19556 14484 19612
rect 14484 19556 14540 19612
rect 14540 19556 14544 19612
rect 14480 19552 14544 19556
rect 14560 19612 14624 19616
rect 14560 19556 14564 19612
rect 14564 19556 14620 19612
rect 14620 19556 14624 19612
rect 14560 19552 14624 19556
rect 14640 19612 14704 19616
rect 14640 19556 14644 19612
rect 14644 19556 14700 19612
rect 14700 19556 14704 19612
rect 14640 19552 14704 19556
rect 14720 19612 14784 19616
rect 14720 19556 14724 19612
rect 14724 19556 14780 19612
rect 14780 19556 14784 19612
rect 14720 19552 14784 19556
rect 23813 19612 23877 19616
rect 23813 19556 23817 19612
rect 23817 19556 23873 19612
rect 23873 19556 23877 19612
rect 23813 19552 23877 19556
rect 23893 19612 23957 19616
rect 23893 19556 23897 19612
rect 23897 19556 23953 19612
rect 23953 19556 23957 19612
rect 23893 19552 23957 19556
rect 23973 19612 24037 19616
rect 23973 19556 23977 19612
rect 23977 19556 24033 19612
rect 24033 19556 24037 19612
rect 23973 19552 24037 19556
rect 24053 19612 24117 19616
rect 24053 19556 24057 19612
rect 24057 19556 24113 19612
rect 24113 19556 24117 19612
rect 24053 19552 24117 19556
rect 9813 19068 9877 19072
rect 9813 19012 9817 19068
rect 9817 19012 9873 19068
rect 9873 19012 9877 19068
rect 9813 19008 9877 19012
rect 9893 19068 9957 19072
rect 9893 19012 9897 19068
rect 9897 19012 9953 19068
rect 9953 19012 9957 19068
rect 9893 19008 9957 19012
rect 9973 19068 10037 19072
rect 9973 19012 9977 19068
rect 9977 19012 10033 19068
rect 10033 19012 10037 19068
rect 9973 19008 10037 19012
rect 10053 19068 10117 19072
rect 10053 19012 10057 19068
rect 10057 19012 10113 19068
rect 10113 19012 10117 19068
rect 10053 19008 10117 19012
rect 19146 19068 19210 19072
rect 19146 19012 19150 19068
rect 19150 19012 19206 19068
rect 19206 19012 19210 19068
rect 19146 19008 19210 19012
rect 19226 19068 19290 19072
rect 19226 19012 19230 19068
rect 19230 19012 19286 19068
rect 19286 19012 19290 19068
rect 19226 19008 19290 19012
rect 19306 19068 19370 19072
rect 19306 19012 19310 19068
rect 19310 19012 19366 19068
rect 19366 19012 19370 19068
rect 19306 19008 19370 19012
rect 19386 19068 19450 19072
rect 19386 19012 19390 19068
rect 19390 19012 19446 19068
rect 19446 19012 19450 19068
rect 19386 19008 19450 19012
rect 5146 18524 5210 18528
rect 5146 18468 5150 18524
rect 5150 18468 5206 18524
rect 5206 18468 5210 18524
rect 5146 18464 5210 18468
rect 5226 18524 5290 18528
rect 5226 18468 5230 18524
rect 5230 18468 5286 18524
rect 5286 18468 5290 18524
rect 5226 18464 5290 18468
rect 5306 18524 5370 18528
rect 5306 18468 5310 18524
rect 5310 18468 5366 18524
rect 5366 18468 5370 18524
rect 5306 18464 5370 18468
rect 5386 18524 5450 18528
rect 5386 18468 5390 18524
rect 5390 18468 5446 18524
rect 5446 18468 5450 18524
rect 5386 18464 5450 18468
rect 14480 18524 14544 18528
rect 14480 18468 14484 18524
rect 14484 18468 14540 18524
rect 14540 18468 14544 18524
rect 14480 18464 14544 18468
rect 14560 18524 14624 18528
rect 14560 18468 14564 18524
rect 14564 18468 14620 18524
rect 14620 18468 14624 18524
rect 14560 18464 14624 18468
rect 14640 18524 14704 18528
rect 14640 18468 14644 18524
rect 14644 18468 14700 18524
rect 14700 18468 14704 18524
rect 14640 18464 14704 18468
rect 14720 18524 14784 18528
rect 14720 18468 14724 18524
rect 14724 18468 14780 18524
rect 14780 18468 14784 18524
rect 14720 18464 14784 18468
rect 23813 18524 23877 18528
rect 23813 18468 23817 18524
rect 23817 18468 23873 18524
rect 23873 18468 23877 18524
rect 23813 18464 23877 18468
rect 23893 18524 23957 18528
rect 23893 18468 23897 18524
rect 23897 18468 23953 18524
rect 23953 18468 23957 18524
rect 23893 18464 23957 18468
rect 23973 18524 24037 18528
rect 23973 18468 23977 18524
rect 23977 18468 24033 18524
rect 24033 18468 24037 18524
rect 23973 18464 24037 18468
rect 24053 18524 24117 18528
rect 24053 18468 24057 18524
rect 24057 18468 24113 18524
rect 24113 18468 24117 18524
rect 24053 18464 24117 18468
rect 9813 17980 9877 17984
rect 9813 17924 9817 17980
rect 9817 17924 9873 17980
rect 9873 17924 9877 17980
rect 9813 17920 9877 17924
rect 9893 17980 9957 17984
rect 9893 17924 9897 17980
rect 9897 17924 9953 17980
rect 9953 17924 9957 17980
rect 9893 17920 9957 17924
rect 9973 17980 10037 17984
rect 9973 17924 9977 17980
rect 9977 17924 10033 17980
rect 10033 17924 10037 17980
rect 9973 17920 10037 17924
rect 10053 17980 10117 17984
rect 10053 17924 10057 17980
rect 10057 17924 10113 17980
rect 10113 17924 10117 17980
rect 10053 17920 10117 17924
rect 19146 17980 19210 17984
rect 19146 17924 19150 17980
rect 19150 17924 19206 17980
rect 19206 17924 19210 17980
rect 19146 17920 19210 17924
rect 19226 17980 19290 17984
rect 19226 17924 19230 17980
rect 19230 17924 19286 17980
rect 19286 17924 19290 17980
rect 19226 17920 19290 17924
rect 19306 17980 19370 17984
rect 19306 17924 19310 17980
rect 19310 17924 19366 17980
rect 19366 17924 19370 17980
rect 19306 17920 19370 17924
rect 19386 17980 19450 17984
rect 19386 17924 19390 17980
rect 19390 17924 19446 17980
rect 19446 17924 19450 17980
rect 19386 17920 19450 17924
rect 5146 17436 5210 17440
rect 5146 17380 5150 17436
rect 5150 17380 5206 17436
rect 5206 17380 5210 17436
rect 5146 17376 5210 17380
rect 5226 17436 5290 17440
rect 5226 17380 5230 17436
rect 5230 17380 5286 17436
rect 5286 17380 5290 17436
rect 5226 17376 5290 17380
rect 5306 17436 5370 17440
rect 5306 17380 5310 17436
rect 5310 17380 5366 17436
rect 5366 17380 5370 17436
rect 5306 17376 5370 17380
rect 5386 17436 5450 17440
rect 5386 17380 5390 17436
rect 5390 17380 5446 17436
rect 5446 17380 5450 17436
rect 5386 17376 5450 17380
rect 14480 17436 14544 17440
rect 14480 17380 14484 17436
rect 14484 17380 14540 17436
rect 14540 17380 14544 17436
rect 14480 17376 14544 17380
rect 14560 17436 14624 17440
rect 14560 17380 14564 17436
rect 14564 17380 14620 17436
rect 14620 17380 14624 17436
rect 14560 17376 14624 17380
rect 14640 17436 14704 17440
rect 14640 17380 14644 17436
rect 14644 17380 14700 17436
rect 14700 17380 14704 17436
rect 14640 17376 14704 17380
rect 14720 17436 14784 17440
rect 14720 17380 14724 17436
rect 14724 17380 14780 17436
rect 14780 17380 14784 17436
rect 14720 17376 14784 17380
rect 23813 17436 23877 17440
rect 23813 17380 23817 17436
rect 23817 17380 23873 17436
rect 23873 17380 23877 17436
rect 23813 17376 23877 17380
rect 23893 17436 23957 17440
rect 23893 17380 23897 17436
rect 23897 17380 23953 17436
rect 23953 17380 23957 17436
rect 23893 17376 23957 17380
rect 23973 17436 24037 17440
rect 23973 17380 23977 17436
rect 23977 17380 24033 17436
rect 24033 17380 24037 17436
rect 23973 17376 24037 17380
rect 24053 17436 24117 17440
rect 24053 17380 24057 17436
rect 24057 17380 24113 17436
rect 24113 17380 24117 17436
rect 24053 17376 24117 17380
rect 9813 16892 9877 16896
rect 9813 16836 9817 16892
rect 9817 16836 9873 16892
rect 9873 16836 9877 16892
rect 9813 16832 9877 16836
rect 9893 16892 9957 16896
rect 9893 16836 9897 16892
rect 9897 16836 9953 16892
rect 9953 16836 9957 16892
rect 9893 16832 9957 16836
rect 9973 16892 10037 16896
rect 9973 16836 9977 16892
rect 9977 16836 10033 16892
rect 10033 16836 10037 16892
rect 9973 16832 10037 16836
rect 10053 16892 10117 16896
rect 10053 16836 10057 16892
rect 10057 16836 10113 16892
rect 10113 16836 10117 16892
rect 10053 16832 10117 16836
rect 19146 16892 19210 16896
rect 19146 16836 19150 16892
rect 19150 16836 19206 16892
rect 19206 16836 19210 16892
rect 19146 16832 19210 16836
rect 19226 16892 19290 16896
rect 19226 16836 19230 16892
rect 19230 16836 19286 16892
rect 19286 16836 19290 16892
rect 19226 16832 19290 16836
rect 19306 16892 19370 16896
rect 19306 16836 19310 16892
rect 19310 16836 19366 16892
rect 19366 16836 19370 16892
rect 19306 16832 19370 16836
rect 19386 16892 19450 16896
rect 19386 16836 19390 16892
rect 19390 16836 19446 16892
rect 19446 16836 19450 16892
rect 19386 16832 19450 16836
rect 5146 16348 5210 16352
rect 5146 16292 5150 16348
rect 5150 16292 5206 16348
rect 5206 16292 5210 16348
rect 5146 16288 5210 16292
rect 5226 16348 5290 16352
rect 5226 16292 5230 16348
rect 5230 16292 5286 16348
rect 5286 16292 5290 16348
rect 5226 16288 5290 16292
rect 5306 16348 5370 16352
rect 5306 16292 5310 16348
rect 5310 16292 5366 16348
rect 5366 16292 5370 16348
rect 5306 16288 5370 16292
rect 5386 16348 5450 16352
rect 5386 16292 5390 16348
rect 5390 16292 5446 16348
rect 5446 16292 5450 16348
rect 5386 16288 5450 16292
rect 14480 16348 14544 16352
rect 14480 16292 14484 16348
rect 14484 16292 14540 16348
rect 14540 16292 14544 16348
rect 14480 16288 14544 16292
rect 14560 16348 14624 16352
rect 14560 16292 14564 16348
rect 14564 16292 14620 16348
rect 14620 16292 14624 16348
rect 14560 16288 14624 16292
rect 14640 16348 14704 16352
rect 14640 16292 14644 16348
rect 14644 16292 14700 16348
rect 14700 16292 14704 16348
rect 14640 16288 14704 16292
rect 14720 16348 14784 16352
rect 14720 16292 14724 16348
rect 14724 16292 14780 16348
rect 14780 16292 14784 16348
rect 14720 16288 14784 16292
rect 23813 16348 23877 16352
rect 23813 16292 23817 16348
rect 23817 16292 23873 16348
rect 23873 16292 23877 16348
rect 23813 16288 23877 16292
rect 23893 16348 23957 16352
rect 23893 16292 23897 16348
rect 23897 16292 23953 16348
rect 23953 16292 23957 16348
rect 23893 16288 23957 16292
rect 23973 16348 24037 16352
rect 23973 16292 23977 16348
rect 23977 16292 24033 16348
rect 24033 16292 24037 16348
rect 23973 16288 24037 16292
rect 24053 16348 24117 16352
rect 24053 16292 24057 16348
rect 24057 16292 24113 16348
rect 24113 16292 24117 16348
rect 24053 16288 24117 16292
rect 23324 16008 23388 16012
rect 23324 15952 23338 16008
rect 23338 15952 23388 16008
rect 23324 15948 23388 15952
rect 9813 15804 9877 15808
rect 9813 15748 9817 15804
rect 9817 15748 9873 15804
rect 9873 15748 9877 15804
rect 9813 15744 9877 15748
rect 9893 15804 9957 15808
rect 9893 15748 9897 15804
rect 9897 15748 9953 15804
rect 9953 15748 9957 15804
rect 9893 15744 9957 15748
rect 9973 15804 10037 15808
rect 9973 15748 9977 15804
rect 9977 15748 10033 15804
rect 10033 15748 10037 15804
rect 9973 15744 10037 15748
rect 10053 15804 10117 15808
rect 10053 15748 10057 15804
rect 10057 15748 10113 15804
rect 10113 15748 10117 15804
rect 10053 15744 10117 15748
rect 19146 15804 19210 15808
rect 19146 15748 19150 15804
rect 19150 15748 19206 15804
rect 19206 15748 19210 15804
rect 19146 15744 19210 15748
rect 19226 15804 19290 15808
rect 19226 15748 19230 15804
rect 19230 15748 19286 15804
rect 19286 15748 19290 15804
rect 19226 15744 19290 15748
rect 19306 15804 19370 15808
rect 19306 15748 19310 15804
rect 19310 15748 19366 15804
rect 19366 15748 19370 15804
rect 19306 15744 19370 15748
rect 19386 15804 19450 15808
rect 19386 15748 19390 15804
rect 19390 15748 19446 15804
rect 19446 15748 19450 15804
rect 19386 15744 19450 15748
rect 5146 15260 5210 15264
rect 5146 15204 5150 15260
rect 5150 15204 5206 15260
rect 5206 15204 5210 15260
rect 5146 15200 5210 15204
rect 5226 15260 5290 15264
rect 5226 15204 5230 15260
rect 5230 15204 5286 15260
rect 5286 15204 5290 15260
rect 5226 15200 5290 15204
rect 5306 15260 5370 15264
rect 5306 15204 5310 15260
rect 5310 15204 5366 15260
rect 5366 15204 5370 15260
rect 5306 15200 5370 15204
rect 5386 15260 5450 15264
rect 5386 15204 5390 15260
rect 5390 15204 5446 15260
rect 5446 15204 5450 15260
rect 5386 15200 5450 15204
rect 14480 15260 14544 15264
rect 14480 15204 14484 15260
rect 14484 15204 14540 15260
rect 14540 15204 14544 15260
rect 14480 15200 14544 15204
rect 14560 15260 14624 15264
rect 14560 15204 14564 15260
rect 14564 15204 14620 15260
rect 14620 15204 14624 15260
rect 14560 15200 14624 15204
rect 14640 15260 14704 15264
rect 14640 15204 14644 15260
rect 14644 15204 14700 15260
rect 14700 15204 14704 15260
rect 14640 15200 14704 15204
rect 14720 15260 14784 15264
rect 14720 15204 14724 15260
rect 14724 15204 14780 15260
rect 14780 15204 14784 15260
rect 14720 15200 14784 15204
rect 23813 15260 23877 15264
rect 23813 15204 23817 15260
rect 23817 15204 23873 15260
rect 23873 15204 23877 15260
rect 23813 15200 23877 15204
rect 23893 15260 23957 15264
rect 23893 15204 23897 15260
rect 23897 15204 23953 15260
rect 23953 15204 23957 15260
rect 23893 15200 23957 15204
rect 23973 15260 24037 15264
rect 23973 15204 23977 15260
rect 23977 15204 24033 15260
rect 24033 15204 24037 15260
rect 23973 15200 24037 15204
rect 24053 15260 24117 15264
rect 24053 15204 24057 15260
rect 24057 15204 24113 15260
rect 24113 15204 24117 15260
rect 24053 15200 24117 15204
rect 9813 14716 9877 14720
rect 9813 14660 9817 14716
rect 9817 14660 9873 14716
rect 9873 14660 9877 14716
rect 9813 14656 9877 14660
rect 9893 14716 9957 14720
rect 9893 14660 9897 14716
rect 9897 14660 9953 14716
rect 9953 14660 9957 14716
rect 9893 14656 9957 14660
rect 9973 14716 10037 14720
rect 9973 14660 9977 14716
rect 9977 14660 10033 14716
rect 10033 14660 10037 14716
rect 9973 14656 10037 14660
rect 10053 14716 10117 14720
rect 10053 14660 10057 14716
rect 10057 14660 10113 14716
rect 10113 14660 10117 14716
rect 10053 14656 10117 14660
rect 19146 14716 19210 14720
rect 19146 14660 19150 14716
rect 19150 14660 19206 14716
rect 19206 14660 19210 14716
rect 19146 14656 19210 14660
rect 19226 14716 19290 14720
rect 19226 14660 19230 14716
rect 19230 14660 19286 14716
rect 19286 14660 19290 14716
rect 19226 14656 19290 14660
rect 19306 14716 19370 14720
rect 19306 14660 19310 14716
rect 19310 14660 19366 14716
rect 19366 14660 19370 14716
rect 19306 14656 19370 14660
rect 19386 14716 19450 14720
rect 19386 14660 19390 14716
rect 19390 14660 19446 14716
rect 19446 14660 19450 14716
rect 19386 14656 19450 14660
rect 5146 14172 5210 14176
rect 5146 14116 5150 14172
rect 5150 14116 5206 14172
rect 5206 14116 5210 14172
rect 5146 14112 5210 14116
rect 5226 14172 5290 14176
rect 5226 14116 5230 14172
rect 5230 14116 5286 14172
rect 5286 14116 5290 14172
rect 5226 14112 5290 14116
rect 5306 14172 5370 14176
rect 5306 14116 5310 14172
rect 5310 14116 5366 14172
rect 5366 14116 5370 14172
rect 5306 14112 5370 14116
rect 5386 14172 5450 14176
rect 5386 14116 5390 14172
rect 5390 14116 5446 14172
rect 5446 14116 5450 14172
rect 5386 14112 5450 14116
rect 14480 14172 14544 14176
rect 14480 14116 14484 14172
rect 14484 14116 14540 14172
rect 14540 14116 14544 14172
rect 14480 14112 14544 14116
rect 14560 14172 14624 14176
rect 14560 14116 14564 14172
rect 14564 14116 14620 14172
rect 14620 14116 14624 14172
rect 14560 14112 14624 14116
rect 14640 14172 14704 14176
rect 14640 14116 14644 14172
rect 14644 14116 14700 14172
rect 14700 14116 14704 14172
rect 14640 14112 14704 14116
rect 14720 14172 14784 14176
rect 14720 14116 14724 14172
rect 14724 14116 14780 14172
rect 14780 14116 14784 14172
rect 14720 14112 14784 14116
rect 23813 14172 23877 14176
rect 23813 14116 23817 14172
rect 23817 14116 23873 14172
rect 23873 14116 23877 14172
rect 23813 14112 23877 14116
rect 23893 14172 23957 14176
rect 23893 14116 23897 14172
rect 23897 14116 23953 14172
rect 23953 14116 23957 14172
rect 23893 14112 23957 14116
rect 23973 14172 24037 14176
rect 23973 14116 23977 14172
rect 23977 14116 24033 14172
rect 24033 14116 24037 14172
rect 23973 14112 24037 14116
rect 24053 14172 24117 14176
rect 24053 14116 24057 14172
rect 24057 14116 24113 14172
rect 24113 14116 24117 14172
rect 24053 14112 24117 14116
rect 9813 13628 9877 13632
rect 9813 13572 9817 13628
rect 9817 13572 9873 13628
rect 9873 13572 9877 13628
rect 9813 13568 9877 13572
rect 9893 13628 9957 13632
rect 9893 13572 9897 13628
rect 9897 13572 9953 13628
rect 9953 13572 9957 13628
rect 9893 13568 9957 13572
rect 9973 13628 10037 13632
rect 9973 13572 9977 13628
rect 9977 13572 10033 13628
rect 10033 13572 10037 13628
rect 9973 13568 10037 13572
rect 10053 13628 10117 13632
rect 10053 13572 10057 13628
rect 10057 13572 10113 13628
rect 10113 13572 10117 13628
rect 10053 13568 10117 13572
rect 19146 13628 19210 13632
rect 19146 13572 19150 13628
rect 19150 13572 19206 13628
rect 19206 13572 19210 13628
rect 19146 13568 19210 13572
rect 19226 13628 19290 13632
rect 19226 13572 19230 13628
rect 19230 13572 19286 13628
rect 19286 13572 19290 13628
rect 19226 13568 19290 13572
rect 19306 13628 19370 13632
rect 19306 13572 19310 13628
rect 19310 13572 19366 13628
rect 19366 13572 19370 13628
rect 19306 13568 19370 13572
rect 19386 13628 19450 13632
rect 19386 13572 19390 13628
rect 19390 13572 19446 13628
rect 19446 13572 19450 13628
rect 19386 13568 19450 13572
rect 5146 13084 5210 13088
rect 5146 13028 5150 13084
rect 5150 13028 5206 13084
rect 5206 13028 5210 13084
rect 5146 13024 5210 13028
rect 5226 13084 5290 13088
rect 5226 13028 5230 13084
rect 5230 13028 5286 13084
rect 5286 13028 5290 13084
rect 5226 13024 5290 13028
rect 5306 13084 5370 13088
rect 5306 13028 5310 13084
rect 5310 13028 5366 13084
rect 5366 13028 5370 13084
rect 5306 13024 5370 13028
rect 5386 13084 5450 13088
rect 5386 13028 5390 13084
rect 5390 13028 5446 13084
rect 5446 13028 5450 13084
rect 5386 13024 5450 13028
rect 14480 13084 14544 13088
rect 14480 13028 14484 13084
rect 14484 13028 14540 13084
rect 14540 13028 14544 13084
rect 14480 13024 14544 13028
rect 14560 13084 14624 13088
rect 14560 13028 14564 13084
rect 14564 13028 14620 13084
rect 14620 13028 14624 13084
rect 14560 13024 14624 13028
rect 14640 13084 14704 13088
rect 14640 13028 14644 13084
rect 14644 13028 14700 13084
rect 14700 13028 14704 13084
rect 14640 13024 14704 13028
rect 14720 13084 14784 13088
rect 14720 13028 14724 13084
rect 14724 13028 14780 13084
rect 14780 13028 14784 13084
rect 14720 13024 14784 13028
rect 23813 13084 23877 13088
rect 23813 13028 23817 13084
rect 23817 13028 23873 13084
rect 23873 13028 23877 13084
rect 23813 13024 23877 13028
rect 23893 13084 23957 13088
rect 23893 13028 23897 13084
rect 23897 13028 23953 13084
rect 23953 13028 23957 13084
rect 23893 13024 23957 13028
rect 23973 13084 24037 13088
rect 23973 13028 23977 13084
rect 23977 13028 24033 13084
rect 24033 13028 24037 13084
rect 23973 13024 24037 13028
rect 24053 13084 24117 13088
rect 24053 13028 24057 13084
rect 24057 13028 24113 13084
rect 24113 13028 24117 13084
rect 24053 13024 24117 13028
rect 9813 12540 9877 12544
rect 9813 12484 9817 12540
rect 9817 12484 9873 12540
rect 9873 12484 9877 12540
rect 9813 12480 9877 12484
rect 9893 12540 9957 12544
rect 9893 12484 9897 12540
rect 9897 12484 9953 12540
rect 9953 12484 9957 12540
rect 9893 12480 9957 12484
rect 9973 12540 10037 12544
rect 9973 12484 9977 12540
rect 9977 12484 10033 12540
rect 10033 12484 10037 12540
rect 9973 12480 10037 12484
rect 10053 12540 10117 12544
rect 10053 12484 10057 12540
rect 10057 12484 10113 12540
rect 10113 12484 10117 12540
rect 10053 12480 10117 12484
rect 19146 12540 19210 12544
rect 19146 12484 19150 12540
rect 19150 12484 19206 12540
rect 19206 12484 19210 12540
rect 19146 12480 19210 12484
rect 19226 12540 19290 12544
rect 19226 12484 19230 12540
rect 19230 12484 19286 12540
rect 19286 12484 19290 12540
rect 19226 12480 19290 12484
rect 19306 12540 19370 12544
rect 19306 12484 19310 12540
rect 19310 12484 19366 12540
rect 19366 12484 19370 12540
rect 19306 12480 19370 12484
rect 19386 12540 19450 12544
rect 19386 12484 19390 12540
rect 19390 12484 19446 12540
rect 19446 12484 19450 12540
rect 19386 12480 19450 12484
rect 23324 12200 23388 12204
rect 23324 12144 23374 12200
rect 23374 12144 23388 12200
rect 23324 12140 23388 12144
rect 5146 11996 5210 12000
rect 5146 11940 5150 11996
rect 5150 11940 5206 11996
rect 5206 11940 5210 11996
rect 5146 11936 5210 11940
rect 5226 11996 5290 12000
rect 5226 11940 5230 11996
rect 5230 11940 5286 11996
rect 5286 11940 5290 11996
rect 5226 11936 5290 11940
rect 5306 11996 5370 12000
rect 5306 11940 5310 11996
rect 5310 11940 5366 11996
rect 5366 11940 5370 11996
rect 5306 11936 5370 11940
rect 5386 11996 5450 12000
rect 5386 11940 5390 11996
rect 5390 11940 5446 11996
rect 5446 11940 5450 11996
rect 5386 11936 5450 11940
rect 14480 11996 14544 12000
rect 14480 11940 14484 11996
rect 14484 11940 14540 11996
rect 14540 11940 14544 11996
rect 14480 11936 14544 11940
rect 14560 11996 14624 12000
rect 14560 11940 14564 11996
rect 14564 11940 14620 11996
rect 14620 11940 14624 11996
rect 14560 11936 14624 11940
rect 14640 11996 14704 12000
rect 14640 11940 14644 11996
rect 14644 11940 14700 11996
rect 14700 11940 14704 11996
rect 14640 11936 14704 11940
rect 14720 11996 14784 12000
rect 14720 11940 14724 11996
rect 14724 11940 14780 11996
rect 14780 11940 14784 11996
rect 14720 11936 14784 11940
rect 23813 11996 23877 12000
rect 23813 11940 23817 11996
rect 23817 11940 23873 11996
rect 23873 11940 23877 11996
rect 23813 11936 23877 11940
rect 23893 11996 23957 12000
rect 23893 11940 23897 11996
rect 23897 11940 23953 11996
rect 23953 11940 23957 11996
rect 23893 11936 23957 11940
rect 23973 11996 24037 12000
rect 23973 11940 23977 11996
rect 23977 11940 24033 11996
rect 24033 11940 24037 11996
rect 23973 11936 24037 11940
rect 24053 11996 24117 12000
rect 24053 11940 24057 11996
rect 24057 11940 24113 11996
rect 24113 11940 24117 11996
rect 24053 11936 24117 11940
rect 9813 11452 9877 11456
rect 9813 11396 9817 11452
rect 9817 11396 9873 11452
rect 9873 11396 9877 11452
rect 9813 11392 9877 11396
rect 9893 11452 9957 11456
rect 9893 11396 9897 11452
rect 9897 11396 9953 11452
rect 9953 11396 9957 11452
rect 9893 11392 9957 11396
rect 9973 11452 10037 11456
rect 9973 11396 9977 11452
rect 9977 11396 10033 11452
rect 10033 11396 10037 11452
rect 9973 11392 10037 11396
rect 10053 11452 10117 11456
rect 10053 11396 10057 11452
rect 10057 11396 10113 11452
rect 10113 11396 10117 11452
rect 10053 11392 10117 11396
rect 19146 11452 19210 11456
rect 19146 11396 19150 11452
rect 19150 11396 19206 11452
rect 19206 11396 19210 11452
rect 19146 11392 19210 11396
rect 19226 11452 19290 11456
rect 19226 11396 19230 11452
rect 19230 11396 19286 11452
rect 19286 11396 19290 11452
rect 19226 11392 19290 11396
rect 19306 11452 19370 11456
rect 19306 11396 19310 11452
rect 19310 11396 19366 11452
rect 19366 11396 19370 11452
rect 19306 11392 19370 11396
rect 19386 11452 19450 11456
rect 19386 11396 19390 11452
rect 19390 11396 19446 11452
rect 19446 11396 19450 11452
rect 19386 11392 19450 11396
rect 5146 10908 5210 10912
rect 5146 10852 5150 10908
rect 5150 10852 5206 10908
rect 5206 10852 5210 10908
rect 5146 10848 5210 10852
rect 5226 10908 5290 10912
rect 5226 10852 5230 10908
rect 5230 10852 5286 10908
rect 5286 10852 5290 10908
rect 5226 10848 5290 10852
rect 5306 10908 5370 10912
rect 5306 10852 5310 10908
rect 5310 10852 5366 10908
rect 5366 10852 5370 10908
rect 5306 10848 5370 10852
rect 5386 10908 5450 10912
rect 5386 10852 5390 10908
rect 5390 10852 5446 10908
rect 5446 10852 5450 10908
rect 5386 10848 5450 10852
rect 14480 10908 14544 10912
rect 14480 10852 14484 10908
rect 14484 10852 14540 10908
rect 14540 10852 14544 10908
rect 14480 10848 14544 10852
rect 14560 10908 14624 10912
rect 14560 10852 14564 10908
rect 14564 10852 14620 10908
rect 14620 10852 14624 10908
rect 14560 10848 14624 10852
rect 14640 10908 14704 10912
rect 14640 10852 14644 10908
rect 14644 10852 14700 10908
rect 14700 10852 14704 10908
rect 14640 10848 14704 10852
rect 14720 10908 14784 10912
rect 14720 10852 14724 10908
rect 14724 10852 14780 10908
rect 14780 10852 14784 10908
rect 14720 10848 14784 10852
rect 23813 10908 23877 10912
rect 23813 10852 23817 10908
rect 23817 10852 23873 10908
rect 23873 10852 23877 10908
rect 23813 10848 23877 10852
rect 23893 10908 23957 10912
rect 23893 10852 23897 10908
rect 23897 10852 23953 10908
rect 23953 10852 23957 10908
rect 23893 10848 23957 10852
rect 23973 10908 24037 10912
rect 23973 10852 23977 10908
rect 23977 10852 24033 10908
rect 24033 10852 24037 10908
rect 23973 10848 24037 10852
rect 24053 10908 24117 10912
rect 24053 10852 24057 10908
rect 24057 10852 24113 10908
rect 24113 10852 24117 10908
rect 24053 10848 24117 10852
rect 9813 10364 9877 10368
rect 9813 10308 9817 10364
rect 9817 10308 9873 10364
rect 9873 10308 9877 10364
rect 9813 10304 9877 10308
rect 9893 10364 9957 10368
rect 9893 10308 9897 10364
rect 9897 10308 9953 10364
rect 9953 10308 9957 10364
rect 9893 10304 9957 10308
rect 9973 10364 10037 10368
rect 9973 10308 9977 10364
rect 9977 10308 10033 10364
rect 10033 10308 10037 10364
rect 9973 10304 10037 10308
rect 10053 10364 10117 10368
rect 10053 10308 10057 10364
rect 10057 10308 10113 10364
rect 10113 10308 10117 10364
rect 10053 10304 10117 10308
rect 19146 10364 19210 10368
rect 19146 10308 19150 10364
rect 19150 10308 19206 10364
rect 19206 10308 19210 10364
rect 19146 10304 19210 10308
rect 19226 10364 19290 10368
rect 19226 10308 19230 10364
rect 19230 10308 19286 10364
rect 19286 10308 19290 10364
rect 19226 10304 19290 10308
rect 19306 10364 19370 10368
rect 19306 10308 19310 10364
rect 19310 10308 19366 10364
rect 19366 10308 19370 10364
rect 19306 10304 19370 10308
rect 19386 10364 19450 10368
rect 19386 10308 19390 10364
rect 19390 10308 19446 10364
rect 19446 10308 19450 10364
rect 19386 10304 19450 10308
rect 5146 9820 5210 9824
rect 5146 9764 5150 9820
rect 5150 9764 5206 9820
rect 5206 9764 5210 9820
rect 5146 9760 5210 9764
rect 5226 9820 5290 9824
rect 5226 9764 5230 9820
rect 5230 9764 5286 9820
rect 5286 9764 5290 9820
rect 5226 9760 5290 9764
rect 5306 9820 5370 9824
rect 5306 9764 5310 9820
rect 5310 9764 5366 9820
rect 5366 9764 5370 9820
rect 5306 9760 5370 9764
rect 5386 9820 5450 9824
rect 5386 9764 5390 9820
rect 5390 9764 5446 9820
rect 5446 9764 5450 9820
rect 5386 9760 5450 9764
rect 14480 9820 14544 9824
rect 14480 9764 14484 9820
rect 14484 9764 14540 9820
rect 14540 9764 14544 9820
rect 14480 9760 14544 9764
rect 14560 9820 14624 9824
rect 14560 9764 14564 9820
rect 14564 9764 14620 9820
rect 14620 9764 14624 9820
rect 14560 9760 14624 9764
rect 14640 9820 14704 9824
rect 14640 9764 14644 9820
rect 14644 9764 14700 9820
rect 14700 9764 14704 9820
rect 14640 9760 14704 9764
rect 14720 9820 14784 9824
rect 14720 9764 14724 9820
rect 14724 9764 14780 9820
rect 14780 9764 14784 9820
rect 14720 9760 14784 9764
rect 23813 9820 23877 9824
rect 23813 9764 23817 9820
rect 23817 9764 23873 9820
rect 23873 9764 23877 9820
rect 23813 9760 23877 9764
rect 23893 9820 23957 9824
rect 23893 9764 23897 9820
rect 23897 9764 23953 9820
rect 23953 9764 23957 9820
rect 23893 9760 23957 9764
rect 23973 9820 24037 9824
rect 23973 9764 23977 9820
rect 23977 9764 24033 9820
rect 24033 9764 24037 9820
rect 23973 9760 24037 9764
rect 24053 9820 24117 9824
rect 24053 9764 24057 9820
rect 24057 9764 24113 9820
rect 24113 9764 24117 9820
rect 24053 9760 24117 9764
rect 9813 9276 9877 9280
rect 9813 9220 9817 9276
rect 9817 9220 9873 9276
rect 9873 9220 9877 9276
rect 9813 9216 9877 9220
rect 9893 9276 9957 9280
rect 9893 9220 9897 9276
rect 9897 9220 9953 9276
rect 9953 9220 9957 9276
rect 9893 9216 9957 9220
rect 9973 9276 10037 9280
rect 9973 9220 9977 9276
rect 9977 9220 10033 9276
rect 10033 9220 10037 9276
rect 9973 9216 10037 9220
rect 10053 9276 10117 9280
rect 10053 9220 10057 9276
rect 10057 9220 10113 9276
rect 10113 9220 10117 9276
rect 10053 9216 10117 9220
rect 19146 9276 19210 9280
rect 19146 9220 19150 9276
rect 19150 9220 19206 9276
rect 19206 9220 19210 9276
rect 19146 9216 19210 9220
rect 19226 9276 19290 9280
rect 19226 9220 19230 9276
rect 19230 9220 19286 9276
rect 19286 9220 19290 9276
rect 19226 9216 19290 9220
rect 19306 9276 19370 9280
rect 19306 9220 19310 9276
rect 19310 9220 19366 9276
rect 19366 9220 19370 9276
rect 19306 9216 19370 9220
rect 19386 9276 19450 9280
rect 19386 9220 19390 9276
rect 19390 9220 19446 9276
rect 19446 9220 19450 9276
rect 19386 9216 19450 9220
rect 5146 8732 5210 8736
rect 5146 8676 5150 8732
rect 5150 8676 5206 8732
rect 5206 8676 5210 8732
rect 5146 8672 5210 8676
rect 5226 8732 5290 8736
rect 5226 8676 5230 8732
rect 5230 8676 5286 8732
rect 5286 8676 5290 8732
rect 5226 8672 5290 8676
rect 5306 8732 5370 8736
rect 5306 8676 5310 8732
rect 5310 8676 5366 8732
rect 5366 8676 5370 8732
rect 5306 8672 5370 8676
rect 5386 8732 5450 8736
rect 5386 8676 5390 8732
rect 5390 8676 5446 8732
rect 5446 8676 5450 8732
rect 5386 8672 5450 8676
rect 14480 8732 14544 8736
rect 14480 8676 14484 8732
rect 14484 8676 14540 8732
rect 14540 8676 14544 8732
rect 14480 8672 14544 8676
rect 14560 8732 14624 8736
rect 14560 8676 14564 8732
rect 14564 8676 14620 8732
rect 14620 8676 14624 8732
rect 14560 8672 14624 8676
rect 14640 8732 14704 8736
rect 14640 8676 14644 8732
rect 14644 8676 14700 8732
rect 14700 8676 14704 8732
rect 14640 8672 14704 8676
rect 14720 8732 14784 8736
rect 14720 8676 14724 8732
rect 14724 8676 14780 8732
rect 14780 8676 14784 8732
rect 14720 8672 14784 8676
rect 23813 8732 23877 8736
rect 23813 8676 23817 8732
rect 23817 8676 23873 8732
rect 23873 8676 23877 8732
rect 23813 8672 23877 8676
rect 23893 8732 23957 8736
rect 23893 8676 23897 8732
rect 23897 8676 23953 8732
rect 23953 8676 23957 8732
rect 23893 8672 23957 8676
rect 23973 8732 24037 8736
rect 23973 8676 23977 8732
rect 23977 8676 24033 8732
rect 24033 8676 24037 8732
rect 23973 8672 24037 8676
rect 24053 8732 24117 8736
rect 24053 8676 24057 8732
rect 24057 8676 24113 8732
rect 24113 8676 24117 8732
rect 24053 8672 24117 8676
rect 9813 8188 9877 8192
rect 9813 8132 9817 8188
rect 9817 8132 9873 8188
rect 9873 8132 9877 8188
rect 9813 8128 9877 8132
rect 9893 8188 9957 8192
rect 9893 8132 9897 8188
rect 9897 8132 9953 8188
rect 9953 8132 9957 8188
rect 9893 8128 9957 8132
rect 9973 8188 10037 8192
rect 9973 8132 9977 8188
rect 9977 8132 10033 8188
rect 10033 8132 10037 8188
rect 9973 8128 10037 8132
rect 10053 8188 10117 8192
rect 10053 8132 10057 8188
rect 10057 8132 10113 8188
rect 10113 8132 10117 8188
rect 10053 8128 10117 8132
rect 19146 8188 19210 8192
rect 19146 8132 19150 8188
rect 19150 8132 19206 8188
rect 19206 8132 19210 8188
rect 19146 8128 19210 8132
rect 19226 8188 19290 8192
rect 19226 8132 19230 8188
rect 19230 8132 19286 8188
rect 19286 8132 19290 8188
rect 19226 8128 19290 8132
rect 19306 8188 19370 8192
rect 19306 8132 19310 8188
rect 19310 8132 19366 8188
rect 19366 8132 19370 8188
rect 19306 8128 19370 8132
rect 19386 8188 19450 8192
rect 19386 8132 19390 8188
rect 19390 8132 19446 8188
rect 19446 8132 19450 8188
rect 19386 8128 19450 8132
rect 7684 7848 7748 7852
rect 7684 7792 7734 7848
rect 7734 7792 7748 7848
rect 7684 7788 7748 7792
rect 5146 7644 5210 7648
rect 5146 7588 5150 7644
rect 5150 7588 5206 7644
rect 5206 7588 5210 7644
rect 5146 7584 5210 7588
rect 5226 7644 5290 7648
rect 5226 7588 5230 7644
rect 5230 7588 5286 7644
rect 5286 7588 5290 7644
rect 5226 7584 5290 7588
rect 5306 7644 5370 7648
rect 5306 7588 5310 7644
rect 5310 7588 5366 7644
rect 5366 7588 5370 7644
rect 5306 7584 5370 7588
rect 5386 7644 5450 7648
rect 5386 7588 5390 7644
rect 5390 7588 5446 7644
rect 5446 7588 5450 7644
rect 5386 7584 5450 7588
rect 14480 7644 14544 7648
rect 14480 7588 14484 7644
rect 14484 7588 14540 7644
rect 14540 7588 14544 7644
rect 14480 7584 14544 7588
rect 14560 7644 14624 7648
rect 14560 7588 14564 7644
rect 14564 7588 14620 7644
rect 14620 7588 14624 7644
rect 14560 7584 14624 7588
rect 14640 7644 14704 7648
rect 14640 7588 14644 7644
rect 14644 7588 14700 7644
rect 14700 7588 14704 7644
rect 14640 7584 14704 7588
rect 14720 7644 14784 7648
rect 14720 7588 14724 7644
rect 14724 7588 14780 7644
rect 14780 7588 14784 7644
rect 14720 7584 14784 7588
rect 23813 7644 23877 7648
rect 23813 7588 23817 7644
rect 23817 7588 23873 7644
rect 23873 7588 23877 7644
rect 23813 7584 23877 7588
rect 23893 7644 23957 7648
rect 23893 7588 23897 7644
rect 23897 7588 23953 7644
rect 23953 7588 23957 7644
rect 23893 7584 23957 7588
rect 23973 7644 24037 7648
rect 23973 7588 23977 7644
rect 23977 7588 24033 7644
rect 24033 7588 24037 7644
rect 23973 7584 24037 7588
rect 24053 7644 24117 7648
rect 24053 7588 24057 7644
rect 24057 7588 24113 7644
rect 24113 7588 24117 7644
rect 24053 7584 24117 7588
rect 9813 7100 9877 7104
rect 9813 7044 9817 7100
rect 9817 7044 9873 7100
rect 9873 7044 9877 7100
rect 9813 7040 9877 7044
rect 9893 7100 9957 7104
rect 9893 7044 9897 7100
rect 9897 7044 9953 7100
rect 9953 7044 9957 7100
rect 9893 7040 9957 7044
rect 9973 7100 10037 7104
rect 9973 7044 9977 7100
rect 9977 7044 10033 7100
rect 10033 7044 10037 7100
rect 9973 7040 10037 7044
rect 10053 7100 10117 7104
rect 10053 7044 10057 7100
rect 10057 7044 10113 7100
rect 10113 7044 10117 7100
rect 10053 7040 10117 7044
rect 19146 7100 19210 7104
rect 19146 7044 19150 7100
rect 19150 7044 19206 7100
rect 19206 7044 19210 7100
rect 19146 7040 19210 7044
rect 19226 7100 19290 7104
rect 19226 7044 19230 7100
rect 19230 7044 19286 7100
rect 19286 7044 19290 7100
rect 19226 7040 19290 7044
rect 19306 7100 19370 7104
rect 19306 7044 19310 7100
rect 19310 7044 19366 7100
rect 19366 7044 19370 7100
rect 19306 7040 19370 7044
rect 19386 7100 19450 7104
rect 19386 7044 19390 7100
rect 19390 7044 19446 7100
rect 19446 7044 19450 7100
rect 19386 7040 19450 7044
rect 22956 6836 23020 6900
rect 5146 6556 5210 6560
rect 5146 6500 5150 6556
rect 5150 6500 5206 6556
rect 5206 6500 5210 6556
rect 5146 6496 5210 6500
rect 5226 6556 5290 6560
rect 5226 6500 5230 6556
rect 5230 6500 5286 6556
rect 5286 6500 5290 6556
rect 5226 6496 5290 6500
rect 5306 6556 5370 6560
rect 5306 6500 5310 6556
rect 5310 6500 5366 6556
rect 5366 6500 5370 6556
rect 5306 6496 5370 6500
rect 5386 6556 5450 6560
rect 5386 6500 5390 6556
rect 5390 6500 5446 6556
rect 5446 6500 5450 6556
rect 5386 6496 5450 6500
rect 14480 6556 14544 6560
rect 14480 6500 14484 6556
rect 14484 6500 14540 6556
rect 14540 6500 14544 6556
rect 14480 6496 14544 6500
rect 14560 6556 14624 6560
rect 14560 6500 14564 6556
rect 14564 6500 14620 6556
rect 14620 6500 14624 6556
rect 14560 6496 14624 6500
rect 14640 6556 14704 6560
rect 14640 6500 14644 6556
rect 14644 6500 14700 6556
rect 14700 6500 14704 6556
rect 14640 6496 14704 6500
rect 14720 6556 14784 6560
rect 14720 6500 14724 6556
rect 14724 6500 14780 6556
rect 14780 6500 14784 6556
rect 14720 6496 14784 6500
rect 23813 6556 23877 6560
rect 23813 6500 23817 6556
rect 23817 6500 23873 6556
rect 23873 6500 23877 6556
rect 23813 6496 23877 6500
rect 23893 6556 23957 6560
rect 23893 6500 23897 6556
rect 23897 6500 23953 6556
rect 23953 6500 23957 6556
rect 23893 6496 23957 6500
rect 23973 6556 24037 6560
rect 23973 6500 23977 6556
rect 23977 6500 24033 6556
rect 24033 6500 24037 6556
rect 23973 6496 24037 6500
rect 24053 6556 24117 6560
rect 24053 6500 24057 6556
rect 24057 6500 24113 6556
rect 24113 6500 24117 6556
rect 24053 6496 24117 6500
rect 4188 6428 4252 6492
rect 24428 6428 24492 6492
rect 10260 6292 10324 6356
rect 9813 6012 9877 6016
rect 9813 5956 9817 6012
rect 9817 5956 9873 6012
rect 9873 5956 9877 6012
rect 9813 5952 9877 5956
rect 9893 6012 9957 6016
rect 9893 5956 9897 6012
rect 9897 5956 9953 6012
rect 9953 5956 9957 6012
rect 9893 5952 9957 5956
rect 9973 6012 10037 6016
rect 9973 5956 9977 6012
rect 9977 5956 10033 6012
rect 10033 5956 10037 6012
rect 9973 5952 10037 5956
rect 10053 6012 10117 6016
rect 10053 5956 10057 6012
rect 10057 5956 10113 6012
rect 10113 5956 10117 6012
rect 10053 5952 10117 5956
rect 19146 6012 19210 6016
rect 19146 5956 19150 6012
rect 19150 5956 19206 6012
rect 19206 5956 19210 6012
rect 19146 5952 19210 5956
rect 19226 6012 19290 6016
rect 19226 5956 19230 6012
rect 19230 5956 19286 6012
rect 19286 5956 19290 6012
rect 19226 5952 19290 5956
rect 19306 6012 19370 6016
rect 19306 5956 19310 6012
rect 19310 5956 19366 6012
rect 19366 5956 19370 6012
rect 19306 5952 19370 5956
rect 19386 6012 19450 6016
rect 19386 5956 19390 6012
rect 19390 5956 19446 6012
rect 19446 5956 19450 6012
rect 19386 5952 19450 5956
rect 5146 5468 5210 5472
rect 5146 5412 5150 5468
rect 5150 5412 5206 5468
rect 5206 5412 5210 5468
rect 5146 5408 5210 5412
rect 5226 5468 5290 5472
rect 5226 5412 5230 5468
rect 5230 5412 5286 5468
rect 5286 5412 5290 5468
rect 5226 5408 5290 5412
rect 5306 5468 5370 5472
rect 5306 5412 5310 5468
rect 5310 5412 5366 5468
rect 5366 5412 5370 5468
rect 5306 5408 5370 5412
rect 5386 5468 5450 5472
rect 5386 5412 5390 5468
rect 5390 5412 5446 5468
rect 5446 5412 5450 5468
rect 5386 5408 5450 5412
rect 14480 5468 14544 5472
rect 14480 5412 14484 5468
rect 14484 5412 14540 5468
rect 14540 5412 14544 5468
rect 14480 5408 14544 5412
rect 14560 5468 14624 5472
rect 14560 5412 14564 5468
rect 14564 5412 14620 5468
rect 14620 5412 14624 5468
rect 14560 5408 14624 5412
rect 14640 5468 14704 5472
rect 14640 5412 14644 5468
rect 14644 5412 14700 5468
rect 14700 5412 14704 5468
rect 14640 5408 14704 5412
rect 14720 5468 14784 5472
rect 14720 5412 14724 5468
rect 14724 5412 14780 5468
rect 14780 5412 14784 5468
rect 14720 5408 14784 5412
rect 23813 5468 23877 5472
rect 23813 5412 23817 5468
rect 23817 5412 23873 5468
rect 23873 5412 23877 5468
rect 23813 5408 23877 5412
rect 23893 5468 23957 5472
rect 23893 5412 23897 5468
rect 23897 5412 23953 5468
rect 23953 5412 23957 5468
rect 23893 5408 23957 5412
rect 23973 5468 24037 5472
rect 23973 5412 23977 5468
rect 23977 5412 24033 5468
rect 24033 5412 24037 5468
rect 23973 5408 24037 5412
rect 24053 5468 24117 5472
rect 24053 5412 24057 5468
rect 24057 5412 24113 5468
rect 24113 5412 24117 5468
rect 24053 5408 24117 5412
rect 22036 5068 22100 5132
rect 9813 4924 9877 4928
rect 9813 4868 9817 4924
rect 9817 4868 9873 4924
rect 9873 4868 9877 4924
rect 9813 4864 9877 4868
rect 9893 4924 9957 4928
rect 9893 4868 9897 4924
rect 9897 4868 9953 4924
rect 9953 4868 9957 4924
rect 9893 4864 9957 4868
rect 9973 4924 10037 4928
rect 9973 4868 9977 4924
rect 9977 4868 10033 4924
rect 10033 4868 10037 4924
rect 9973 4864 10037 4868
rect 10053 4924 10117 4928
rect 10053 4868 10057 4924
rect 10057 4868 10113 4924
rect 10113 4868 10117 4924
rect 10053 4864 10117 4868
rect 19146 4924 19210 4928
rect 19146 4868 19150 4924
rect 19150 4868 19206 4924
rect 19206 4868 19210 4924
rect 19146 4864 19210 4868
rect 19226 4924 19290 4928
rect 19226 4868 19230 4924
rect 19230 4868 19286 4924
rect 19286 4868 19290 4924
rect 19226 4864 19290 4868
rect 19306 4924 19370 4928
rect 19306 4868 19310 4924
rect 19310 4868 19366 4924
rect 19366 4868 19370 4924
rect 19306 4864 19370 4868
rect 19386 4924 19450 4928
rect 19386 4868 19390 4924
rect 19390 4868 19446 4924
rect 19446 4868 19450 4924
rect 19386 4864 19450 4868
rect 10260 4796 10324 4860
rect 5146 4380 5210 4384
rect 5146 4324 5150 4380
rect 5150 4324 5206 4380
rect 5206 4324 5210 4380
rect 5146 4320 5210 4324
rect 5226 4380 5290 4384
rect 5226 4324 5230 4380
rect 5230 4324 5286 4380
rect 5286 4324 5290 4380
rect 5226 4320 5290 4324
rect 5306 4380 5370 4384
rect 5306 4324 5310 4380
rect 5310 4324 5366 4380
rect 5366 4324 5370 4380
rect 5306 4320 5370 4324
rect 5386 4380 5450 4384
rect 5386 4324 5390 4380
rect 5390 4324 5446 4380
rect 5446 4324 5450 4380
rect 5386 4320 5450 4324
rect 14480 4380 14544 4384
rect 14480 4324 14484 4380
rect 14484 4324 14540 4380
rect 14540 4324 14544 4380
rect 14480 4320 14544 4324
rect 14560 4380 14624 4384
rect 14560 4324 14564 4380
rect 14564 4324 14620 4380
rect 14620 4324 14624 4380
rect 14560 4320 14624 4324
rect 14640 4380 14704 4384
rect 14640 4324 14644 4380
rect 14644 4324 14700 4380
rect 14700 4324 14704 4380
rect 14640 4320 14704 4324
rect 14720 4380 14784 4384
rect 14720 4324 14724 4380
rect 14724 4324 14780 4380
rect 14780 4324 14784 4380
rect 14720 4320 14784 4324
rect 23813 4380 23877 4384
rect 23813 4324 23817 4380
rect 23817 4324 23873 4380
rect 23873 4324 23877 4380
rect 23813 4320 23877 4324
rect 23893 4380 23957 4384
rect 23893 4324 23897 4380
rect 23897 4324 23953 4380
rect 23953 4324 23957 4380
rect 23893 4320 23957 4324
rect 23973 4380 24037 4384
rect 23973 4324 23977 4380
rect 23977 4324 24033 4380
rect 24033 4324 24037 4380
rect 23973 4320 24037 4324
rect 24053 4380 24117 4384
rect 24053 4324 24057 4380
rect 24057 4324 24113 4380
rect 24113 4324 24117 4380
rect 24053 4320 24117 4324
rect 9813 3836 9877 3840
rect 9813 3780 9817 3836
rect 9817 3780 9873 3836
rect 9873 3780 9877 3836
rect 9813 3776 9877 3780
rect 9893 3836 9957 3840
rect 9893 3780 9897 3836
rect 9897 3780 9953 3836
rect 9953 3780 9957 3836
rect 9893 3776 9957 3780
rect 9973 3836 10037 3840
rect 9973 3780 9977 3836
rect 9977 3780 10033 3836
rect 10033 3780 10037 3836
rect 9973 3776 10037 3780
rect 10053 3836 10117 3840
rect 10053 3780 10057 3836
rect 10057 3780 10113 3836
rect 10113 3780 10117 3836
rect 10053 3776 10117 3780
rect 6212 3708 6276 3772
rect 19146 3836 19210 3840
rect 19146 3780 19150 3836
rect 19150 3780 19206 3836
rect 19206 3780 19210 3836
rect 19146 3776 19210 3780
rect 19226 3836 19290 3840
rect 19226 3780 19230 3836
rect 19230 3780 19286 3836
rect 19286 3780 19290 3836
rect 19226 3776 19290 3780
rect 19306 3836 19370 3840
rect 19306 3780 19310 3836
rect 19310 3780 19366 3836
rect 19366 3780 19370 3836
rect 19306 3776 19370 3780
rect 19386 3836 19450 3840
rect 19386 3780 19390 3836
rect 19390 3780 19446 3836
rect 19446 3780 19450 3836
rect 19386 3776 19450 3780
rect 5146 3292 5210 3296
rect 5146 3236 5150 3292
rect 5150 3236 5206 3292
rect 5206 3236 5210 3292
rect 5146 3232 5210 3236
rect 5226 3292 5290 3296
rect 5226 3236 5230 3292
rect 5230 3236 5286 3292
rect 5286 3236 5290 3292
rect 5226 3232 5290 3236
rect 5306 3292 5370 3296
rect 5306 3236 5310 3292
rect 5310 3236 5366 3292
rect 5366 3236 5370 3292
rect 5306 3232 5370 3236
rect 5386 3292 5450 3296
rect 5386 3236 5390 3292
rect 5390 3236 5446 3292
rect 5446 3236 5450 3292
rect 5386 3232 5450 3236
rect 14480 3292 14544 3296
rect 14480 3236 14484 3292
rect 14484 3236 14540 3292
rect 14540 3236 14544 3292
rect 14480 3232 14544 3236
rect 14560 3292 14624 3296
rect 14560 3236 14564 3292
rect 14564 3236 14620 3292
rect 14620 3236 14624 3292
rect 14560 3232 14624 3236
rect 14640 3292 14704 3296
rect 14640 3236 14644 3292
rect 14644 3236 14700 3292
rect 14700 3236 14704 3292
rect 14640 3232 14704 3236
rect 14720 3292 14784 3296
rect 14720 3236 14724 3292
rect 14724 3236 14780 3292
rect 14780 3236 14784 3292
rect 14720 3232 14784 3236
rect 23813 3292 23877 3296
rect 23813 3236 23817 3292
rect 23817 3236 23873 3292
rect 23873 3236 23877 3292
rect 23813 3232 23877 3236
rect 23893 3292 23957 3296
rect 23893 3236 23897 3292
rect 23897 3236 23953 3292
rect 23953 3236 23957 3292
rect 23893 3232 23957 3236
rect 23973 3292 24037 3296
rect 23973 3236 23977 3292
rect 23977 3236 24033 3292
rect 24033 3236 24037 3292
rect 23973 3232 24037 3236
rect 24053 3292 24117 3296
rect 24053 3236 24057 3292
rect 24057 3236 24113 3292
rect 24113 3236 24117 3292
rect 24053 3232 24117 3236
rect 7684 3028 7748 3092
rect 9813 2748 9877 2752
rect 9813 2692 9817 2748
rect 9817 2692 9873 2748
rect 9873 2692 9877 2748
rect 9813 2688 9877 2692
rect 9893 2748 9957 2752
rect 9893 2692 9897 2748
rect 9897 2692 9953 2748
rect 9953 2692 9957 2748
rect 9893 2688 9957 2692
rect 9973 2748 10037 2752
rect 9973 2692 9977 2748
rect 9977 2692 10033 2748
rect 10033 2692 10037 2748
rect 9973 2688 10037 2692
rect 10053 2748 10117 2752
rect 10053 2692 10057 2748
rect 10057 2692 10113 2748
rect 10113 2692 10117 2748
rect 10053 2688 10117 2692
rect 19146 2748 19210 2752
rect 19146 2692 19150 2748
rect 19150 2692 19206 2748
rect 19206 2692 19210 2748
rect 19146 2688 19210 2692
rect 19226 2748 19290 2752
rect 19226 2692 19230 2748
rect 19230 2692 19286 2748
rect 19286 2692 19290 2748
rect 19226 2688 19290 2692
rect 19306 2748 19370 2752
rect 19306 2692 19310 2748
rect 19310 2692 19366 2748
rect 19366 2692 19370 2748
rect 19306 2688 19370 2692
rect 19386 2748 19450 2752
rect 19386 2692 19390 2748
rect 19390 2692 19446 2748
rect 19446 2692 19450 2748
rect 19386 2688 19450 2692
rect 22220 2408 22284 2412
rect 22220 2352 22270 2408
rect 22270 2352 22284 2408
rect 22220 2348 22284 2352
rect 5146 2204 5210 2208
rect 5146 2148 5150 2204
rect 5150 2148 5206 2204
rect 5206 2148 5210 2204
rect 5146 2144 5210 2148
rect 5226 2204 5290 2208
rect 5226 2148 5230 2204
rect 5230 2148 5286 2204
rect 5286 2148 5290 2204
rect 5226 2144 5290 2148
rect 5306 2204 5370 2208
rect 5306 2148 5310 2204
rect 5310 2148 5366 2204
rect 5366 2148 5370 2204
rect 5306 2144 5370 2148
rect 5386 2204 5450 2208
rect 5386 2148 5390 2204
rect 5390 2148 5446 2204
rect 5446 2148 5450 2204
rect 5386 2144 5450 2148
rect 14480 2204 14544 2208
rect 14480 2148 14484 2204
rect 14484 2148 14540 2204
rect 14540 2148 14544 2204
rect 14480 2144 14544 2148
rect 14560 2204 14624 2208
rect 14560 2148 14564 2204
rect 14564 2148 14620 2204
rect 14620 2148 14624 2204
rect 14560 2144 14624 2148
rect 14640 2204 14704 2208
rect 14640 2148 14644 2204
rect 14644 2148 14700 2204
rect 14700 2148 14704 2204
rect 14640 2144 14704 2148
rect 14720 2204 14784 2208
rect 14720 2148 14724 2204
rect 14724 2148 14780 2204
rect 14780 2148 14784 2204
rect 14720 2144 14784 2148
rect 23813 2204 23877 2208
rect 23813 2148 23817 2204
rect 23817 2148 23873 2204
rect 23873 2148 23877 2204
rect 23813 2144 23877 2148
rect 23893 2204 23957 2208
rect 23893 2148 23897 2204
rect 23897 2148 23953 2204
rect 23953 2148 23957 2204
rect 23893 2144 23957 2148
rect 23973 2204 24037 2208
rect 23973 2148 23977 2204
rect 23977 2148 24033 2204
rect 24033 2148 24037 2204
rect 23973 2144 24037 2148
rect 24053 2204 24117 2208
rect 24053 2148 24057 2204
rect 24057 2148 24113 2204
rect 24113 2148 24117 2204
rect 24053 2144 24117 2148
rect 2164 1728 2228 1732
rect 2164 1672 2178 1728
rect 2178 1672 2228 1728
rect 2164 1668 2228 1672
rect 26820 1728 26884 1732
rect 26820 1672 26870 1728
rect 26870 1672 26884 1728
rect 26820 1668 26884 1672
<< metal4 >>
rect 5138 25056 5459 25616
rect 5138 24992 5146 25056
rect 5210 24992 5226 25056
rect 5290 24992 5306 25056
rect 5370 24992 5386 25056
rect 5450 24992 5459 25056
rect 5138 23968 5459 24992
rect 5138 23904 5146 23968
rect 5210 23904 5226 23968
rect 5290 23904 5306 23968
rect 5370 23904 5386 23968
rect 5450 23904 5459 23968
rect 5138 22880 5459 23904
rect 5138 22816 5146 22880
rect 5210 22816 5226 22880
rect 5290 22816 5306 22880
rect 5370 22816 5386 22880
rect 5450 22816 5459 22880
rect 5138 21792 5459 22816
rect 5138 21728 5146 21792
rect 5210 21728 5226 21792
rect 5290 21728 5306 21792
rect 5370 21728 5386 21792
rect 5450 21728 5459 21792
rect 5138 20704 5459 21728
rect 5138 20640 5146 20704
rect 5210 20640 5226 20704
rect 5290 20640 5306 20704
rect 5370 20640 5386 20704
rect 5450 20640 5459 20704
rect 5138 19616 5459 20640
rect 5138 19552 5146 19616
rect 5210 19552 5226 19616
rect 5290 19552 5306 19616
rect 5370 19552 5386 19616
rect 5450 19552 5459 19616
rect 5138 18528 5459 19552
rect 5138 18464 5146 18528
rect 5210 18464 5226 18528
rect 5290 18464 5306 18528
rect 5370 18464 5386 18528
rect 5450 18464 5459 18528
rect 5138 17440 5459 18464
rect 5138 17376 5146 17440
rect 5210 17376 5226 17440
rect 5290 17376 5306 17440
rect 5370 17376 5386 17440
rect 5450 17376 5459 17440
rect 5138 16352 5459 17376
rect 5138 16288 5146 16352
rect 5210 16288 5226 16352
rect 5290 16288 5306 16352
rect 5370 16288 5386 16352
rect 5450 16288 5459 16352
rect 5138 15264 5459 16288
rect 5138 15200 5146 15264
rect 5210 15200 5226 15264
rect 5290 15200 5306 15264
rect 5370 15200 5386 15264
rect 5450 15200 5459 15264
rect 5138 14176 5459 15200
rect 5138 14112 5146 14176
rect 5210 14112 5226 14176
rect 5290 14112 5306 14176
rect 5370 14112 5386 14176
rect 5450 14112 5459 14176
rect 5138 13088 5459 14112
rect 5138 13024 5146 13088
rect 5210 13024 5226 13088
rect 5290 13024 5306 13088
rect 5370 13024 5386 13088
rect 5450 13024 5459 13088
rect 5138 12000 5459 13024
rect 5138 11936 5146 12000
rect 5210 11936 5226 12000
rect 5290 11936 5306 12000
rect 5370 11936 5386 12000
rect 5450 11936 5459 12000
rect 5138 10912 5459 11936
rect 5138 10848 5146 10912
rect 5210 10848 5226 10912
rect 5290 10848 5306 10912
rect 5370 10848 5386 10912
rect 5450 10848 5459 10912
rect 5138 9824 5459 10848
rect 5138 9760 5146 9824
rect 5210 9760 5226 9824
rect 5290 9760 5306 9824
rect 5370 9760 5386 9824
rect 5450 9760 5459 9824
rect 5138 8736 5459 9760
rect 5138 8672 5146 8736
rect 5210 8672 5226 8736
rect 5290 8672 5306 8736
rect 5370 8672 5386 8736
rect 5450 8672 5459 8736
rect 5138 7648 5459 8672
rect 9805 25600 10125 25616
rect 9805 25536 9813 25600
rect 9877 25536 9893 25600
rect 9957 25536 9973 25600
rect 10037 25536 10053 25600
rect 10117 25536 10125 25600
rect 9805 24512 10125 25536
rect 9805 24448 9813 24512
rect 9877 24448 9893 24512
rect 9957 24448 9973 24512
rect 10037 24448 10053 24512
rect 10117 24448 10125 24512
rect 9805 23424 10125 24448
rect 9805 23360 9813 23424
rect 9877 23360 9893 23424
rect 9957 23360 9973 23424
rect 10037 23360 10053 23424
rect 10117 23360 10125 23424
rect 9805 22336 10125 23360
rect 9805 22272 9813 22336
rect 9877 22272 9893 22336
rect 9957 22272 9973 22336
rect 10037 22272 10053 22336
rect 10117 22272 10125 22336
rect 9805 21248 10125 22272
rect 9805 21184 9813 21248
rect 9877 21184 9893 21248
rect 9957 21184 9973 21248
rect 10037 21184 10053 21248
rect 10117 21184 10125 21248
rect 9805 20160 10125 21184
rect 9805 20096 9813 20160
rect 9877 20096 9893 20160
rect 9957 20096 9973 20160
rect 10037 20096 10053 20160
rect 10117 20096 10125 20160
rect 9805 19072 10125 20096
rect 9805 19008 9813 19072
rect 9877 19008 9893 19072
rect 9957 19008 9973 19072
rect 10037 19008 10053 19072
rect 10117 19008 10125 19072
rect 9805 17984 10125 19008
rect 9805 17920 9813 17984
rect 9877 17920 9893 17984
rect 9957 17920 9973 17984
rect 10037 17920 10053 17984
rect 10117 17920 10125 17984
rect 9805 16896 10125 17920
rect 9805 16832 9813 16896
rect 9877 16832 9893 16896
rect 9957 16832 9973 16896
rect 10037 16832 10053 16896
rect 10117 16832 10125 16896
rect 9805 15808 10125 16832
rect 9805 15744 9813 15808
rect 9877 15744 9893 15808
rect 9957 15744 9973 15808
rect 10037 15744 10053 15808
rect 10117 15744 10125 15808
rect 9805 14720 10125 15744
rect 9805 14656 9813 14720
rect 9877 14656 9893 14720
rect 9957 14656 9973 14720
rect 10037 14656 10053 14720
rect 10117 14656 10125 14720
rect 9805 13632 10125 14656
rect 9805 13568 9813 13632
rect 9877 13568 9893 13632
rect 9957 13568 9973 13632
rect 10037 13568 10053 13632
rect 10117 13568 10125 13632
rect 9805 12544 10125 13568
rect 9805 12480 9813 12544
rect 9877 12480 9893 12544
rect 9957 12480 9973 12544
rect 10037 12480 10053 12544
rect 10117 12480 10125 12544
rect 9805 11456 10125 12480
rect 9805 11392 9813 11456
rect 9877 11392 9893 11456
rect 9957 11392 9973 11456
rect 10037 11392 10053 11456
rect 10117 11392 10125 11456
rect 9805 10368 10125 11392
rect 9805 10304 9813 10368
rect 9877 10304 9893 10368
rect 9957 10304 9973 10368
rect 10037 10304 10053 10368
rect 10117 10304 10125 10368
rect 9805 9280 10125 10304
rect 9805 9216 9813 9280
rect 9877 9216 9893 9280
rect 9957 9216 9973 9280
rect 10037 9216 10053 9280
rect 10117 9216 10125 9280
rect 9805 8192 10125 9216
rect 9805 8128 9813 8192
rect 9877 8128 9893 8192
rect 9957 8128 9973 8192
rect 10037 8128 10053 8192
rect 10117 8128 10125 8192
rect 5138 7584 5146 7648
rect 5210 7584 5226 7648
rect 5290 7584 5306 7648
rect 5370 7584 5386 7648
rect 5450 7584 5459 7648
rect 5138 6560 5459 7584
rect 5138 6496 5146 6560
rect 5210 6496 5226 6560
rect 5290 6496 5306 6560
rect 5370 6496 5386 6560
rect 5450 6496 5459 6560
rect 5138 5472 5459 6496
rect 5138 5408 5146 5472
rect 5210 5408 5226 5472
rect 5290 5408 5306 5472
rect 5370 5408 5386 5472
rect 5450 5408 5459 5472
rect 5138 4384 5459 5408
rect 9805 7104 10125 8128
rect 9805 7040 9813 7104
rect 9877 7040 9893 7104
rect 9957 7040 9973 7104
rect 10037 7040 10053 7104
rect 10117 7040 10125 7104
rect 9805 6016 10125 7040
rect 14472 25056 14792 25616
rect 14472 24992 14480 25056
rect 14544 24992 14560 25056
rect 14624 24992 14640 25056
rect 14704 24992 14720 25056
rect 14784 24992 14792 25056
rect 14472 23968 14792 24992
rect 14472 23904 14480 23968
rect 14544 23904 14560 23968
rect 14624 23904 14640 23968
rect 14704 23904 14720 23968
rect 14784 23904 14792 23968
rect 14472 22880 14792 23904
rect 14472 22816 14480 22880
rect 14544 22816 14560 22880
rect 14624 22816 14640 22880
rect 14704 22816 14720 22880
rect 14784 22816 14792 22880
rect 14472 21792 14792 22816
rect 14472 21728 14480 21792
rect 14544 21728 14560 21792
rect 14624 21728 14640 21792
rect 14704 21728 14720 21792
rect 14784 21728 14792 21792
rect 14472 20704 14792 21728
rect 14472 20640 14480 20704
rect 14544 20640 14560 20704
rect 14624 20640 14640 20704
rect 14704 20640 14720 20704
rect 14784 20640 14792 20704
rect 14472 19616 14792 20640
rect 14472 19552 14480 19616
rect 14544 19552 14560 19616
rect 14624 19552 14640 19616
rect 14704 19552 14720 19616
rect 14784 19552 14792 19616
rect 14472 18528 14792 19552
rect 14472 18464 14480 18528
rect 14544 18464 14560 18528
rect 14624 18464 14640 18528
rect 14704 18464 14720 18528
rect 14784 18464 14792 18528
rect 14472 17440 14792 18464
rect 14472 17376 14480 17440
rect 14544 17376 14560 17440
rect 14624 17376 14640 17440
rect 14704 17376 14720 17440
rect 14784 17376 14792 17440
rect 14472 16352 14792 17376
rect 14472 16288 14480 16352
rect 14544 16288 14560 16352
rect 14624 16288 14640 16352
rect 14704 16288 14720 16352
rect 14784 16288 14792 16352
rect 14472 15264 14792 16288
rect 14472 15200 14480 15264
rect 14544 15200 14560 15264
rect 14624 15200 14640 15264
rect 14704 15200 14720 15264
rect 14784 15200 14792 15264
rect 14472 14176 14792 15200
rect 14472 14112 14480 14176
rect 14544 14112 14560 14176
rect 14624 14112 14640 14176
rect 14704 14112 14720 14176
rect 14784 14112 14792 14176
rect 14472 13088 14792 14112
rect 14472 13024 14480 13088
rect 14544 13024 14560 13088
rect 14624 13024 14640 13088
rect 14704 13024 14720 13088
rect 14784 13024 14792 13088
rect 14472 12000 14792 13024
rect 14472 11936 14480 12000
rect 14544 11936 14560 12000
rect 14624 11936 14640 12000
rect 14704 11936 14720 12000
rect 14784 11936 14792 12000
rect 14472 10912 14792 11936
rect 14472 10848 14480 10912
rect 14544 10848 14560 10912
rect 14624 10848 14640 10912
rect 14704 10848 14720 10912
rect 14784 10848 14792 10912
rect 14472 9824 14792 10848
rect 14472 9760 14480 9824
rect 14544 9760 14560 9824
rect 14624 9760 14640 9824
rect 14704 9760 14720 9824
rect 14784 9760 14792 9824
rect 14472 8736 14792 9760
rect 14472 8672 14480 8736
rect 14544 8672 14560 8736
rect 14624 8672 14640 8736
rect 14704 8672 14720 8736
rect 14784 8672 14792 8736
rect 14472 7648 14792 8672
rect 14472 7584 14480 7648
rect 14544 7584 14560 7648
rect 14624 7584 14640 7648
rect 14704 7584 14720 7648
rect 14784 7584 14792 7648
rect 14472 6560 14792 7584
rect 14472 6496 14480 6560
rect 14544 6496 14560 6560
rect 14624 6496 14640 6560
rect 14704 6496 14720 6560
rect 14784 6496 14792 6560
rect 10259 6356 10325 6357
rect 10259 6292 10260 6356
rect 10324 6292 10325 6356
rect 10259 6291 10325 6292
rect 9805 5952 9813 6016
rect 9877 5952 9893 6016
rect 9957 5952 9973 6016
rect 10037 5952 10053 6016
rect 10117 5952 10125 6016
rect 5138 4320 5146 4384
rect 5210 4320 5226 4384
rect 5290 4320 5306 4384
rect 5370 4320 5386 4384
rect 5450 4320 5459 4384
rect 5138 3296 5459 4320
rect 6214 3773 6274 4982
rect 9805 4928 10125 5952
rect 9805 4864 9813 4928
rect 9877 4864 9893 4928
rect 9957 4864 9973 4928
rect 10037 4864 10053 4928
rect 10117 4864 10125 4928
rect 9805 3840 10125 4864
rect 10262 4861 10322 6291
rect 14472 5472 14792 6496
rect 14472 5408 14480 5472
rect 14544 5408 14560 5472
rect 14624 5408 14640 5472
rect 14704 5408 14720 5472
rect 14784 5408 14792 5472
rect 10259 4860 10325 4861
rect 10259 4796 10260 4860
rect 10324 4796 10325 4860
rect 10259 4795 10325 4796
rect 9805 3776 9813 3840
rect 9877 3776 9893 3840
rect 9957 3776 9973 3840
rect 10037 3776 10053 3840
rect 10117 3776 10125 3840
rect 6211 3772 6277 3773
rect 6211 3708 6212 3772
rect 6276 3708 6277 3772
rect 6211 3707 6277 3708
rect 5138 3232 5146 3296
rect 5210 3232 5226 3296
rect 5290 3232 5306 3296
rect 5370 3232 5386 3296
rect 5450 3232 5459 3296
rect 5138 2208 5459 3232
rect 7683 3092 7749 3093
rect 7683 3028 7684 3092
rect 7748 3028 7749 3092
rect 7683 3027 7749 3028
rect 7686 2498 7746 3027
rect 9805 2752 10125 3776
rect 9805 2688 9813 2752
rect 9877 2688 9893 2752
rect 9957 2688 9973 2752
rect 10037 2688 10053 2752
rect 10117 2688 10125 2752
rect 5138 2144 5146 2208
rect 5210 2144 5226 2208
rect 5290 2144 5306 2208
rect 5370 2144 5386 2208
rect 5450 2144 5459 2208
rect 5138 2128 5459 2144
rect 9805 2128 10125 2688
rect 14472 4384 14792 5408
rect 14472 4320 14480 4384
rect 14544 4320 14560 4384
rect 14624 4320 14640 4384
rect 14704 4320 14720 4384
rect 14784 4320 14792 4384
rect 14472 3296 14792 4320
rect 14472 3232 14480 3296
rect 14544 3232 14560 3296
rect 14624 3232 14640 3296
rect 14704 3232 14720 3296
rect 14784 3232 14792 3296
rect 14472 2208 14792 3232
rect 14472 2144 14480 2208
rect 14544 2144 14560 2208
rect 14624 2144 14640 2208
rect 14704 2144 14720 2208
rect 14784 2144 14792 2208
rect 14472 2128 14792 2144
rect 19138 25600 19458 25616
rect 19138 25536 19146 25600
rect 19210 25536 19226 25600
rect 19290 25536 19306 25600
rect 19370 25536 19386 25600
rect 19450 25536 19458 25600
rect 19138 24512 19458 25536
rect 19138 24448 19146 24512
rect 19210 24448 19226 24512
rect 19290 24448 19306 24512
rect 19370 24448 19386 24512
rect 19450 24448 19458 24512
rect 19138 23424 19458 24448
rect 19138 23360 19146 23424
rect 19210 23360 19226 23424
rect 19290 23360 19306 23424
rect 19370 23360 19386 23424
rect 19450 23360 19458 23424
rect 19138 22336 19458 23360
rect 19138 22272 19146 22336
rect 19210 22272 19226 22336
rect 19290 22272 19306 22336
rect 19370 22272 19386 22336
rect 19450 22272 19458 22336
rect 19138 21248 19458 22272
rect 19138 21184 19146 21248
rect 19210 21184 19226 21248
rect 19290 21184 19306 21248
rect 19370 21184 19386 21248
rect 19450 21184 19458 21248
rect 19138 20160 19458 21184
rect 19138 20096 19146 20160
rect 19210 20096 19226 20160
rect 19290 20096 19306 20160
rect 19370 20096 19386 20160
rect 19450 20096 19458 20160
rect 19138 19072 19458 20096
rect 19138 19008 19146 19072
rect 19210 19008 19226 19072
rect 19290 19008 19306 19072
rect 19370 19008 19386 19072
rect 19450 19008 19458 19072
rect 19138 17984 19458 19008
rect 19138 17920 19146 17984
rect 19210 17920 19226 17984
rect 19290 17920 19306 17984
rect 19370 17920 19386 17984
rect 19450 17920 19458 17984
rect 19138 16896 19458 17920
rect 19138 16832 19146 16896
rect 19210 16832 19226 16896
rect 19290 16832 19306 16896
rect 19370 16832 19386 16896
rect 19450 16832 19458 16896
rect 19138 15808 19458 16832
rect 23805 25056 24125 25616
rect 23805 24992 23813 25056
rect 23877 24992 23893 25056
rect 23957 24992 23973 25056
rect 24037 24992 24053 25056
rect 24117 24992 24125 25056
rect 23805 23968 24125 24992
rect 23805 23904 23813 23968
rect 23877 23904 23893 23968
rect 23957 23904 23973 23968
rect 24037 23904 24053 23968
rect 24117 23904 24125 23968
rect 23805 22880 24125 23904
rect 23805 22816 23813 22880
rect 23877 22816 23893 22880
rect 23957 22816 23973 22880
rect 24037 22816 24053 22880
rect 24117 22816 24125 22880
rect 23805 21792 24125 22816
rect 23805 21728 23813 21792
rect 23877 21728 23893 21792
rect 23957 21728 23973 21792
rect 24037 21728 24053 21792
rect 24117 21728 24125 21792
rect 23805 20704 24125 21728
rect 23805 20640 23813 20704
rect 23877 20640 23893 20704
rect 23957 20640 23973 20704
rect 24037 20640 24053 20704
rect 24117 20640 24125 20704
rect 23805 19616 24125 20640
rect 23805 19552 23813 19616
rect 23877 19552 23893 19616
rect 23957 19552 23973 19616
rect 24037 19552 24053 19616
rect 24117 19552 24125 19616
rect 23805 18528 24125 19552
rect 23805 18464 23813 18528
rect 23877 18464 23893 18528
rect 23957 18464 23973 18528
rect 24037 18464 24053 18528
rect 24117 18464 24125 18528
rect 23805 17440 24125 18464
rect 23805 17376 23813 17440
rect 23877 17376 23893 17440
rect 23957 17376 23973 17440
rect 24037 17376 24053 17440
rect 24117 17376 24125 17440
rect 23805 16352 24125 17376
rect 23805 16288 23813 16352
rect 23877 16288 23893 16352
rect 23957 16288 23973 16352
rect 24037 16288 24053 16352
rect 24117 16288 24125 16352
rect 23323 16012 23389 16013
rect 23323 15948 23324 16012
rect 23388 15948 23389 16012
rect 23323 15947 23389 15948
rect 19138 15744 19146 15808
rect 19210 15744 19226 15808
rect 19290 15744 19306 15808
rect 19370 15744 19386 15808
rect 19450 15744 19458 15808
rect 19138 14720 19458 15744
rect 19138 14656 19146 14720
rect 19210 14656 19226 14720
rect 19290 14656 19306 14720
rect 19370 14656 19386 14720
rect 19450 14656 19458 14720
rect 19138 13632 19458 14656
rect 19138 13568 19146 13632
rect 19210 13568 19226 13632
rect 19290 13568 19306 13632
rect 19370 13568 19386 13632
rect 19450 13568 19458 13632
rect 19138 12544 19458 13568
rect 19138 12480 19146 12544
rect 19210 12480 19226 12544
rect 19290 12480 19306 12544
rect 19370 12480 19386 12544
rect 19450 12480 19458 12544
rect 19138 11456 19458 12480
rect 23326 12205 23386 15947
rect 23805 15264 24125 16288
rect 23805 15200 23813 15264
rect 23877 15200 23893 15264
rect 23957 15200 23973 15264
rect 24037 15200 24053 15264
rect 24117 15200 24125 15264
rect 23805 14176 24125 15200
rect 23805 14112 23813 14176
rect 23877 14112 23893 14176
rect 23957 14112 23973 14176
rect 24037 14112 24053 14176
rect 24117 14112 24125 14176
rect 23805 13088 24125 14112
rect 23805 13024 23813 13088
rect 23877 13024 23893 13088
rect 23957 13024 23973 13088
rect 24037 13024 24053 13088
rect 24117 13024 24125 13088
rect 23323 12204 23389 12205
rect 23323 12140 23324 12204
rect 23388 12140 23389 12204
rect 23323 12139 23389 12140
rect 19138 11392 19146 11456
rect 19210 11392 19226 11456
rect 19290 11392 19306 11456
rect 19370 11392 19386 11456
rect 19450 11392 19458 11456
rect 19138 10368 19458 11392
rect 19138 10304 19146 10368
rect 19210 10304 19226 10368
rect 19290 10304 19306 10368
rect 19370 10304 19386 10368
rect 19450 10304 19458 10368
rect 19138 9280 19458 10304
rect 19138 9216 19146 9280
rect 19210 9216 19226 9280
rect 19290 9216 19306 9280
rect 19370 9216 19386 9280
rect 19450 9216 19458 9280
rect 19138 8192 19458 9216
rect 19138 8128 19146 8192
rect 19210 8128 19226 8192
rect 19290 8128 19306 8192
rect 19370 8128 19386 8192
rect 19450 8128 19458 8192
rect 19138 7104 19458 8128
rect 23805 12000 24125 13024
rect 23805 11936 23813 12000
rect 23877 11936 23893 12000
rect 23957 11936 23973 12000
rect 24037 11936 24053 12000
rect 24117 11936 24125 12000
rect 23805 10912 24125 11936
rect 23805 10848 23813 10912
rect 23877 10848 23893 10912
rect 23957 10848 23973 10912
rect 24037 10848 24053 10912
rect 24117 10848 24125 10912
rect 23805 9824 24125 10848
rect 23805 9760 23813 9824
rect 23877 9760 23893 9824
rect 23957 9760 23973 9824
rect 24037 9760 24053 9824
rect 24117 9760 24125 9824
rect 23805 8736 24125 9760
rect 23805 8672 23813 8736
rect 23877 8672 23893 8736
rect 23957 8672 23973 8736
rect 24037 8672 24053 8736
rect 24117 8672 24125 8736
rect 19138 7040 19146 7104
rect 19210 7040 19226 7104
rect 19290 7040 19306 7104
rect 19370 7040 19386 7104
rect 19450 7040 19458 7104
rect 19138 6016 19458 7040
rect 22958 6901 23018 7702
rect 23805 7648 24125 8672
rect 23805 7584 23813 7648
rect 23877 7584 23893 7648
rect 23957 7584 23973 7648
rect 24037 7584 24053 7648
rect 24117 7584 24125 7648
rect 22955 6900 23021 6901
rect 22955 6836 22956 6900
rect 23020 6836 23021 6900
rect 22955 6835 23021 6836
rect 19138 5952 19146 6016
rect 19210 5952 19226 6016
rect 19290 5952 19306 6016
rect 19370 5952 19386 6016
rect 19450 5952 19458 6016
rect 19138 4928 19458 5952
rect 23805 6560 24125 7584
rect 23805 6496 23813 6560
rect 23877 6496 23893 6560
rect 23957 6496 23973 6560
rect 24037 6496 24053 6560
rect 24117 6496 24125 6560
rect 23805 5472 24125 6496
rect 23805 5408 23813 5472
rect 23877 5408 23893 5472
rect 23957 5408 23973 5472
rect 24037 5408 24053 5472
rect 24117 5408 24125 5472
rect 19138 4864 19146 4928
rect 19210 4864 19226 4928
rect 19290 4864 19306 4928
rect 19370 4864 19386 4928
rect 19450 4864 19458 4928
rect 19138 3840 19458 4864
rect 19138 3776 19146 3840
rect 19210 3776 19226 3840
rect 19290 3776 19306 3840
rect 19370 3776 19386 3840
rect 19450 3776 19458 3840
rect 19138 2752 19458 3776
rect 19138 2688 19146 2752
rect 19210 2688 19226 2752
rect 19290 2688 19306 2752
rect 19370 2688 19386 2752
rect 19450 2688 19458 2752
rect 19138 2128 19458 2688
rect 23805 4384 24125 5408
rect 23805 4320 23813 4384
rect 23877 4320 23893 4384
rect 23957 4320 23973 4384
rect 24037 4320 24053 4384
rect 24117 4320 24125 4384
rect 23805 3296 24125 4320
rect 23805 3232 23813 3296
rect 23877 3232 23893 3296
rect 23957 3232 23973 3296
rect 24037 3232 24053 3296
rect 24117 3232 24125 3296
rect 23805 2208 24125 3232
rect 23805 2144 23813 2208
rect 23877 2144 23893 2208
rect 23957 2144 23973 2208
rect 24037 2144 24053 2208
rect 24117 2144 24125 2208
rect 23805 2128 24125 2144
<< via4 >>
rect 7598 7852 7834 7938
rect 7598 7788 7684 7852
rect 7684 7788 7748 7852
rect 7748 7788 7834 7852
rect 7598 7702 7834 7788
rect 4102 6492 4338 6578
rect 4102 6428 4188 6492
rect 4188 6428 4252 6492
rect 4252 6428 4338 6492
rect 4102 6342 4338 6428
rect 6126 4982 6362 5218
rect 7598 2262 7834 2498
rect 22870 7702 23106 7938
rect 24342 6492 24578 6578
rect 24342 6428 24428 6492
rect 24428 6428 24492 6492
rect 24492 6428 24578 6492
rect 24342 6342 24578 6428
rect 21950 5132 22186 5218
rect 21950 5068 22036 5132
rect 22036 5068 22100 5132
rect 22100 5068 22186 5132
rect 21950 4982 22186 5068
rect 22134 2412 22370 2498
rect 22134 2348 22220 2412
rect 22220 2348 22284 2412
rect 22284 2348 22370 2412
rect 22134 2262 22370 2348
rect 2078 1732 2314 1818
rect 2078 1668 2164 1732
rect 2164 1668 2228 1732
rect 2228 1668 2314 1732
rect 2078 1582 2314 1668
rect 26734 1732 26970 1818
rect 26734 1668 26820 1732
rect 26820 1668 26884 1732
rect 26884 1668 26970 1732
rect 26734 1582 26970 1668
<< metal5 >>
rect 7556 7938 23148 7980
rect 7556 7702 7598 7938
rect 7834 7702 22870 7938
rect 23106 7702 23148 7938
rect 7556 7660 23148 7702
rect 4060 6578 24620 6620
rect 4060 6342 4102 6578
rect 4338 6342 24342 6578
rect 24578 6342 24620 6578
rect 4060 6300 24620 6342
rect 6084 5218 22228 5260
rect 6084 4982 6126 5218
rect 6362 4982 21950 5218
rect 22186 4982 22228 5218
rect 6084 4940 22228 4982
rect 7556 2498 22412 2540
rect 7556 2262 7598 2498
rect 7834 2262 22134 2498
rect 22370 2262 22412 2498
rect 7556 2220 22412 2262
rect 2036 1818 27012 1860
rect 2036 1582 2078 1818
rect 2314 1582 26734 1818
rect 26970 1582 27012 1818
rect 2036 1540 27012 1582
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1460 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 632 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 632 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 908 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_12 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1736 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 908 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_15
timestamp 1586364061
transform 1 0 2012 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_16 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2104 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1920 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2196 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_20
timestamp 1586364061
transform 1 0 2472 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 2748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2656 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2472 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_24
timestamp 1586364061
transform 1 0 2840 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_27
timestamp 1586364061
transform 1 0 3116 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2932 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3208 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4220 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4312 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3484 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3668 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4036 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3576 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_31
timestamp 1586364061
transform 1 0 3484 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_35
timestamp 1586364061
transform 1 0 3852 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_46
timestamp 1586364061
transform 1 0 4864 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_42
timestamp 1586364061
transform 1 0 4496 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_47
timestamp 1586364061
transform 1 0 4956 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_43
timestamp 1586364061
transform 1 0 4588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5048 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4680 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5508 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5692 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5232 0 1 2720
box -38 -48 314 592
use scs8hd_conb_1  _215_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5324 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_54
timestamp 1586364061
transform 1 0 5600 0 -1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6336 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6244 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6060 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_63
timestamp 1586364061
transform 1 0 6428 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 5876 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_62
timestamp 1586364061
transform 1 0 6336 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_74
timestamp 1586364061
transform 1 0 7440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7072 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7256 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7164 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_75
timestamp 1586364061
transform 1 0 7532 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_78
timestamp 1586364061
transform 1 0 7808 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7624 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_81
timestamp 1586364061
transform 1 0 8084 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7900 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8176 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8268 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_86
timestamp 1586364061
transform 1 0 8544 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8452 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_90
timestamp 1586364061
transform 1 0 8912 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 8820 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8728 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8636 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_94
timestamp 1586364061
transform 1 0 9280 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 9004 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9096 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9188 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9280 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9464 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 9924 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 9556 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_99
timestamp 1586364061
transform 1 0 9740 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10108 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9740 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10292 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10292 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _197_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10476 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11120 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11304 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11304 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11488 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 11672 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11672 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11488 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11856 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 11856 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12040 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11948 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12132 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 13144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 12960 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_138
timestamp 1586364061
transform 1 0 13328 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_132
timestamp 1586364061
transform 1 0 12776 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13328 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _240_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13788 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13696 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13512 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 14340 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_142 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13696 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14156 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14524 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_151
timestamp 1586364061
transform 1 0 14524 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_156
timestamp 1586364061
transform 1 0 14984 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 14708 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14800 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 14892 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_162
timestamp 1586364061
transform 1 0 15536 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 15812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 15352 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15720 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 14984 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 15904 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 16640 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16916 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15996 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_169
timestamp 1586364061
transform 1 0 16180 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_173
timestamp 1586364061
transform 1 0 16548 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17008 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 16732 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17100 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17376 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17560 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 17192 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17284 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17468 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 17744 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_193
timestamp 1586364061
transform 1 0 18388 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_187
timestamp 1586364061
transform 1 0 17836 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18204 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17560 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18388 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19216 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19032 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18664 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 19400 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_202
timestamp 1586364061
transform 1 0 19216 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_206
timestamp 1586364061
transform 1 0 19584 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_198
timestamp 1586364061
transform 1 0 18848 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_211
timestamp 1586364061
transform 1 0 20044 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20228 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_210
timestamp 1586364061
transform 1 0 19952 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20044 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_215
timestamp 1586364061
transform 1 0 20412 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 20412 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20596 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20596 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20780 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 20688 0 -1 2720
box -38 -48 866 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 22252 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21976 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_227
timestamp 1586364061
transform 1 0 21516 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_228
timestamp 1586364061
transform 1 0 21608 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_234
timestamp 1586364061
transform 1 0 22160 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_238
timestamp 1586364061
transform 1 0 22528 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_239
timestamp 1586364061
transform 1 0 22620 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 22804 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 22896 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22344 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_243
timestamp 1586364061
transform 1 0 22988 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 23264 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23080 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23448 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 23540 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 23172 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 24736 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24184 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24552 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_258
timestamp 1586364061
transform 1 0 24368 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_254
timestamp 1586364061
transform 1 0 24000 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_258
timestamp 1586364061
transform 1 0 24368 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25104 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25564 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 25288 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_269
timestamp 1586364061
transform 1 0 25380 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 25748 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_266
timestamp 1586364061
transform 1 0 25104 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_270
timestamp 1586364061
transform 1 0 25472 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_276
timestamp 1586364061
transform 1 0 26024 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26392 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26392 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 632 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 908 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2012 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3116 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3852 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3484 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_32
timestamp 1586364061
transform 1 0 3576 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_38
timestamp 1586364061
transform 1 0 4128 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4864 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_49
timestamp 1586364061
transform 1 0 5140 0 -1 3808
box -38 -48 774 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 6888 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5876 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_60
timestamp 1586364061
transform 1 0 6152 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7900 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_71
timestamp 1586364061
transform 1 0 7164 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_82
timestamp 1586364061
transform 1 0 8176 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9096 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9464 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_90
timestamp 1586364061
transform 1 0 8912 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_93
timestamp 1586364061
transform 1 0 9188 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9648 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10660 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_107
timestamp 1586364061
transform 1 0 10476 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11212 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11028 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_111
timestamp 1586364061
transform 1 0 10844 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_124
timestamp 1586364061
transform 1 0 12040 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 13144 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12316 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12684 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_129
timestamp 1586364061
transform 1 0 12500 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_133
timestamp 1586364061
transform 1 0 12868 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14156 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 13972 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_149
timestamp 1586364061
transform 1 0 14340 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15812 0 -1 3808
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14800 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 14708 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 15260 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_157
timestamp 1586364061
transform 1 0 15076 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_161
timestamp 1586364061
transform 1 0 15444 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16824 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_174
timestamp 1586364061
transform 1 0 16640 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_178
timestamp 1586364061
transform 1 0 17008 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17376 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17192 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18388 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_191
timestamp 1586364061
transform 1 0 18204 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 18940 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19492 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_195
timestamp 1586364061
transform 1 0 18572 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_203
timestamp 1586364061
transform 1 0 19308 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_207
timestamp 1586364061
transform 1 0 19676 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20412 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20320 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20136 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_211
timestamp 1586364061
transform 1 0 20044 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21976 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21424 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_224
timestamp 1586364061
transform 1 0 21240 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_228
timestamp 1586364061
transform 1 0 21608 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23540 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23172 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_241
timestamp 1586364061
transform 1 0 22804 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_247
timestamp 1586364061
transform 1 0 23356 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_258
timestamp 1586364061
transform 1 0 24368 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 25932 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_270
timestamp 1586364061
transform 1 0 25472 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 25840 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26024 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26392 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 632 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 908 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2012 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_3_27
timestamp 1586364061
transform 1 0 3116 0 1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3208 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4220 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3668 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_31
timestamp 1586364061
transform 1 0 3484 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_35
timestamp 1586364061
transform 1 0 3852 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5232 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4680 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5048 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5692 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_42
timestamp 1586364061
transform 1 0 4496 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_46
timestamp 1586364061
transform 1 0 4864 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5508 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 6704 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6244 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6060 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 5876 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_62
timestamp 1586364061
transform 1 0 6336 0 1 3808
box -38 -48 406 592
use scs8hd_decap_6  FILLER_3_69
timestamp 1586364061
transform 1 0 6980 0 1 3808
box -38 -48 590 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 7716 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 7532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_80
timestamp 1586364061
transform 1 0 7992 0 1 3808
box -38 -48 590 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 8728 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 8544 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10292 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10108 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_97
timestamp 1586364061
transform 1 0 9556 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 11856 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11304 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11120 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_118
timestamp 1586364061
transform 1 0 11488 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 11948 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12316 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12132 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13328 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13144 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13880 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13696 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_140
timestamp 1586364061
transform 1 0 13512 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 15628 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 15444 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14892 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_153
timestamp 1586364061
transform 1 0 14708 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_157
timestamp 1586364061
transform 1 0 15076 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16640 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_172
timestamp 1586364061
transform 1 0 16456 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_176
timestamp 1586364061
transform 1 0 16824 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17560 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17468 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17284 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_180
timestamp 1586364061
transform 1 0 17192 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18388 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19492 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18572 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19308 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18940 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 18756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_201
timestamp 1586364061
transform 1 0 19124 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20504 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20872 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_214
timestamp 1586364061
transform 1 0 20320 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_218
timestamp 1586364061
transform 1 0 20688 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21424 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21240 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_222
timestamp 1586364061
transform 1 0 21056 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_235
timestamp 1586364061
transform 1 0 22252 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23172 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23080 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22528 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 22712 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 24736 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24184 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_254
timestamp 1586364061
transform 1 0 24000 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_258
timestamp 1586364061
transform 1 0 24368 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 25288 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_266
timestamp 1586364061
transform 1 0 25104 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_270
timestamp 1586364061
transform 1 0 25472 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_276
timestamp 1586364061
transform 1 0 26024 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26392 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 632 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 908 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2012 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3116 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3484 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_32
timestamp 1586364061
transform 1 0 3576 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_40
timestamp 1586364061
transform 1 0 4312 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4496 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5508 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_45
timestamp 1586364061
transform 1 0 4772 0 -1 4896
box -38 -48 774 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 6520 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_56
timestamp 1586364061
transform 1 0 5784 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_8  FILLER_4_67
timestamp 1586364061
transform 1 0 6796 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 7532 0 -1 4896
box -38 -48 866 592
use scs8hd_conb_1  _222_
timestamp 1586364061
transform 1 0 9464 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9096 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_84
timestamp 1586364061
transform 1 0 8360 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_93
timestamp 1586364061
transform 1 0 9188 0 -1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10476 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10292 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_99
timestamp 1586364061
transform 1 0 9740 0 -1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11672 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_118
timestamp 1586364061
transform 1 0 11488 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_122
timestamp 1586364061
transform 1 0 11856 0 -1 4896
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13144 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12500 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12868 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_128
timestamp 1586364061
transform 1 0 12408 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_131
timestamp 1586364061
transform 1 0 12684 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_135
timestamp 1586364061
transform 1 0 13052 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_145
timestamp 1586364061
transform 1 0 13972 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 15076 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 14708 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_154
timestamp 1586364061
transform 1 0 14800 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_161
timestamp 1586364061
transform 1 0 15444 0 -1 4896
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16180 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 18112 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17560 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_180
timestamp 1586364061
transform 1 0 17192 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_186
timestamp 1586364061
transform 1 0 17744 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_4_192
timestamp 1586364061
transform 1 0 18296 0 -1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18572 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_4_206
timestamp 1586364061
transform 1 0 19584 0 -1 4896
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20412 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20320 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 22160 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21976 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_226
timestamp 1586364061
transform 1 0 21424 0 -1 4896
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23448 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 22712 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23264 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_238
timestamp 1586364061
transform 1 0 22528 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_242
timestamp 1586364061
transform 1 0 22896 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_257
timestamp 1586364061
transform 1 0 24276 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 25932 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_269
timestamp 1586364061
transform 1 0 25380 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26024 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26392 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 632 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 908 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2012 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3116 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4220 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5324 0 1 4896
box -38 -48 774 592
use scs8hd_conb_1  _223_
timestamp 1586364061
transform 1 0 6428 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6244 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 6888 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6060 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_62
timestamp 1586364061
transform 1 0 6336 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 6704 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 7440 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 7256 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_70
timestamp 1586364061
transform 1 0 7072 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_83
timestamp 1586364061
transform 1 0 8268 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9004 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8820 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8452 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_87
timestamp 1586364061
transform 1 0 8636 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10016 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10384 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_100
timestamp 1586364061
transform 1 0 9832 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_104
timestamp 1586364061
transform 1 0 10200 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_108
timestamp 1586364061
transform 1 0 10568 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10844 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 11856 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11304 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11672 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11120 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11488 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_123
timestamp 1586364061
transform 1 0 11948 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12500 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12316 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _207_
timestamp 1586364061
transform 1 0 14616 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13696 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 14432 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14064 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_140
timestamp 1586364061
transform 1 0 13512 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_144
timestamp 1586364061
transform 1 0 13880 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_148
timestamp 1586364061
transform 1 0 14248 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15628 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_161
timestamp 1586364061
transform 1 0 15444 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_165
timestamp 1586364061
transform 1 0 15812 0 1 4896
box -38 -48 406 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 16364 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16916 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 16180 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 16732 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17100 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18296 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17468 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18112 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 17744 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17284 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_184
timestamp 1586364061
transform 1 0 17560 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_188
timestamp 1586364061
transform 1 0 17928 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 19676 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_203
timestamp 1586364061
transform 1 0 19308 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20596 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20412 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 20044 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_209
timestamp 1586364061
transform 1 0 19860 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_213
timestamp 1586364061
transform 1 0 20228 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21976 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_228
timestamp 1586364061
transform 1 0 21608 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_234
timestamp 1586364061
transform 1 0 22160 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23448 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23080 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22344 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_238
timestamp 1586364061
transform 1 0 22528 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_5_245
timestamp 1586364061
transform 1 0 23172 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24460 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_257
timestamp 1586364061
transform 1 0 24276 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_261
timestamp 1586364061
transform 1 0 24644 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 25012 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 25564 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24828 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_269
timestamp 1586364061
transform 1 0 25380 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_273
timestamp 1586364061
transform 1 0 25748 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26392 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 632 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 632 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 908 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 908 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2012 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3116 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2012 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3116 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3484 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 3576 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4220 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 4680 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5324 0 1 5984
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6520 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6336 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6244 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6796 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_56
timestamp 1586364061
transform 1 0 5784 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_6_67
timestamp 1586364061
transform 1 0 6796 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6060 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_65
timestamp 1586364061
transform 1 0 6612 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_69
timestamp 1586364061
transform 1 0 6980 0 1 5984
box -38 -48 590 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 7532 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7532 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7992 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_78
timestamp 1586364061
transform 1 0 7808 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_82
timestamp 1586364061
transform 1 0 8176 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 8544 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9464 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9096 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 8360 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8360 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_93
timestamp 1586364061
transform 1 0 9188 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9372 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10108 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9556 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10476 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_105
timestamp 1586364061
transform 1 0 10292 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_109
timestamp 1586364061
transform 1 0 10660 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_99
timestamp 1586364061
transform 1 0 9740 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11948 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11028 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 11856 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11672 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 11304 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10844 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_124
timestamp 1586364061
transform 1 0 12040 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11120 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11488 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12868 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 12224 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12592 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_128
timestamp 1586364061
transform 1 0 12408 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_132
timestamp 1586364061
transform 1 0 12776 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 12960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13328 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14156 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13972 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14156 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13512 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_142
timestamp 1586364061
transform 1 0 13696 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_146
timestamp 1586364061
transform 1 0 14064 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_149
timestamp 1586364061
transform 1 0 14340 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_142
timestamp 1586364061
transform 1 0 13696 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14800 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15904 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 14708 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15720 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 15352 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_165
timestamp 1586364061
transform 1 0 15812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_158
timestamp 1586364061
transform 1 0 15168 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_162
timestamp 1586364061
transform 1 0 15536 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16548 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15996 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_169
timestamp 1586364061
transform 1 0 16180 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_7_175
timestamp 1586364061
transform 1 0 16732 0 1 5984
box -38 -48 590 592
use scs8hd_nor2_4  _105_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18112 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17560 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17468 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17284 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17560 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17928 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_182
timestamp 1586364061
transform 1 0 17376 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_186
timestamp 1586364061
transform 1 0 17744 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 19584 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19124 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_199
timestamp 1586364061
transform 1 0 18940 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_203
timestamp 1586364061
transform 1 0 19308 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_207
timestamp 1586364061
transform 1 0 19676 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_197
timestamp 1586364061
transform 1 0 18756 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_205
timestamp 1586364061
transform 1 0 19492 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 20412 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 19768 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20320 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 19768 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20780 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20136 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_210
timestamp 1586364061
transform 1 0 19952 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_217
timestamp 1586364061
transform 1 0 20596 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_221
timestamp 1586364061
transform 1 0 20964 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21332 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21976 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21148 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21424 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21792 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_224
timestamp 1586364061
transform 1 0 21240 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_228
timestamp 1586364061
transform 1 0 21608 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 22712 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22344 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 22528 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_247
timestamp 1586364061
transform 1 0 23356 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_243
timestamp 1586364061
transform 1 0 22988 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23540 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 23172 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23080 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 23172 0 1 5984
box -38 -48 866 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 24736 0 1 5984
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23724 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 24552 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_260
timestamp 1586364061
transform 1 0 24552 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_254
timestamp 1586364061
transform 1 0 24000 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 25932 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 25288 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 25656 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26024 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_266
timestamp 1586364061
transform 1 0 25104 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_270
timestamp 1586364061
transform 1 0 25472 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_276
timestamp 1586364061
transform 1 0 26024 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26392 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26392 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 632 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 908 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2012 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3116 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3484 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 3576 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 4680 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 5784 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 6888 0 -1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 8084 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_80
timestamp 1586364061
transform 1 0 7992 0 -1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9096 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 8728 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_84
timestamp 1586364061
transform 1 0 8360 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_90
timestamp 1586364061
transform 1 0 8912 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_93
timestamp 1586364061
transform 1 0 9188 0 -1 7072
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9832 0 -1 7072
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_8_99
timestamp 1586364061
transform 1 0 9740 0 -1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 11580 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 11028 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_111
timestamp 1586364061
transform 1 0 10844 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_115
timestamp 1586364061
transform 1 0 11212 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13144 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12592 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_128
timestamp 1586364061
transform 1 0 12408 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_132
timestamp 1586364061
transform 1 0 12776 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 14156 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 13972 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_149
timestamp 1586364061
transform 1 0 14340 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 15812 0 -1 7072
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14800 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 14708 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15260 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15628 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_157
timestamp 1586364061
transform 1 0 15076 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_161
timestamp 1586364061
transform 1 0 15444 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_174
timestamp 1586364061
transform 1 0 16640 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17928 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_8_186
timestamp 1586364061
transform 1 0 17744 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 19584 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 18940 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_197
timestamp 1586364061
transform 1 0 18756 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_201
timestamp 1586364061
transform 1 0 19124 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_205
timestamp 1586364061
transform 1 0 19492 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20412 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20320 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20872 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_208
timestamp 1586364061
transform 1 0 19768 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_8_218
timestamp 1586364061
transform 1 0 20688 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21424 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21240 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_222
timestamp 1586364061
transform 1 0 21056 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_235
timestamp 1586364061
transform 1 0 22252 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23172 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22436 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_239
timestamp 1586364061
transform 1 0 22620 0 -1 7072
box -38 -48 590 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 24736 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_254
timestamp 1586364061
transform 1 0 24000 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 25932 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_266
timestamp 1586364061
transform 1 0 25104 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 25840 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26024 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26392 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 632 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 908 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2012 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3116 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4220 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5324 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6244 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6060 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6336 0 1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 7716 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 7532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_74
timestamp 1586364061
transform 1 0 7440 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_80
timestamp 1586364061
transform 1 0 7992 0 1 7072
box -38 -48 590 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 8728 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 8544 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 10292 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 10108 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 9740 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_97
timestamp 1586364061
transform 1 0 9556 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 9924 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 11948 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 11856 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 11672 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 11304 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11120 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11488 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 13328 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 12960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 12776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13144 0 1 7072
box -38 -48 222 592
use scs8hd_nor3_4  _170_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13880 0 1 7072
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 13696 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_140
timestamp 1586364061
transform 1 0 13512 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 15812 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15260 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 15628 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_157
timestamp 1586364061
transform 1 0 15076 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_161
timestamp 1586364061
transform 1 0 15444 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16824 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_174
timestamp 1586364061
transform 1 0 16640 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_178
timestamp 1586364061
transform 1 0 17008 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18020 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17468 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17836 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17192 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17376 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_184
timestamp 1586364061
transform 1 0 17560 0 1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 19584 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 19400 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 19032 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_198
timestamp 1586364061
transform 1 0 18848 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_202
timestamp 1586364061
transform 1 0 19216 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20964 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20596 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_215
timestamp 1586364061
transform 1 0 20412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_219
timestamp 1586364061
transform 1 0 20780 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21148 0 1 7072
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_9_234
timestamp 1586364061
transform 1 0 22160 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23172 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23080 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22344 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_238
timestamp 1586364061
transform 1 0 22528 0 1 7072
box -38 -48 406 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 24736 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 24184 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24000 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_258
timestamp 1586364061
transform 1 0 24368 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 25288 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_266
timestamp 1586364061
transform 1 0 25104 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_270
timestamp 1586364061
transform 1 0 25472 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_276
timestamp 1586364061
transform 1 0 26024 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26392 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 632 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 908 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2012 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3116 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3484 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 3576 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 4680 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 5784 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_10_68
timestamp 1586364061
transform 1 0 6888 0 -1 8160
box -38 -48 590 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 7532 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_1  FILLER_10_74
timestamp 1586364061
transform 1 0 7440 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 9280 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9096 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8360 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_93
timestamp 1586364061
transform 1 0 9188 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 10292 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 9924 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_97
timestamp 1586364061
transform 1 0 9556 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_103
timestamp 1586364061
transform 1 0 10108 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 11948 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11304 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_114
timestamp 1586364061
transform 1 0 11120 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_118
timestamp 1586364061
transform 1 0 11488 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_122
timestamp 1586364061
transform 1 0 11856 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 13144 0 -1 8160
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12132 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12868 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_128
timestamp 1586364061
transform 1 0 12408 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_132
timestamp 1586364061
transform 1 0 12776 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_135
timestamp 1586364061
transform 1 0 13052 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 14524 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 14156 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 13972 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14340 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14800 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 14708 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_165
timestamp 1586364061
transform 1 0 15812 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16824 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 15996 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16364 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_169
timestamp 1586364061
transform 1 0 16180 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_173
timestamp 1586364061
transform 1 0 16548 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18020 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 18388 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_187
timestamp 1586364061
transform 1 0 17836 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_191
timestamp 1586364061
transform 1 0 18204 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 18756 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_10_195
timestamp 1586364061
transform 1 0 18572 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_206
timestamp 1586364061
transform 1 0 19584 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20412 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20320 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19768 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_210
timestamp 1586364061
transform 1 0 19952 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22160 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21608 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_226
timestamp 1586364061
transform 1 0 21424 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_230
timestamp 1586364061
transform 1 0 21792 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23172 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23540 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_243
timestamp 1586364061
transform 1 0 22988 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_247
timestamp 1586364061
transform 1 0 23356 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 23724 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_260
timestamp 1586364061
transform 1 0 24552 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 25932 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_272
timestamp 1586364061
transform 1 0 25656 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26024 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26392 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 632 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 908 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2012 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3116 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4220 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5324 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6244 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6060 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6336 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7440 0 1 8160
box -38 -48 1142 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 8912 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 9372 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_86
timestamp 1586364061
transform 1 0 8544 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_93
timestamp 1586364061
transform 1 0 9188 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 9924 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 9740 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_97
timestamp 1586364061
transform 1 0 9556 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_110
timestamp 1586364061
transform 1 0 10752 0 1 8160
box -38 -48 406 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 11948 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 11856 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11120 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 11672 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_116
timestamp 1586364061
transform 1 0 11304 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 13328 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 12776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13144 0 1 8160
box -38 -48 222 592
use scs8hd_nor3_4  _171_
timestamp 1586364061
transform 1 0 13512 0 1 8160
box -38 -48 1234 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15444 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15260 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 14892 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_153
timestamp 1586364061
transform 1 0 14708 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_157
timestamp 1586364061
transform 1 0 15076 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16916 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_172
timestamp 1586364061
transform 1 0 16456 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_176
timestamp 1586364061
transform 1 0 16824 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17100 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 17560 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17468 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17284 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_193
timestamp 1586364061
transform 1 0 18388 0 1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 19308 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 19124 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 18756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_199
timestamp 1586364061
transform 1 0 18940 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 20872 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 20688 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_212
timestamp 1586364061
transform 1 0 20136 0 1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21884 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_229
timestamp 1586364061
transform 1 0 21700 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_233
timestamp 1586364061
transform 1 0 22068 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23172 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23080 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22528 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_237
timestamp 1586364061
transform 1 0 22436 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 22712 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 24736 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 24368 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_254
timestamp 1586364061
transform 1 0 24000 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_260
timestamp 1586364061
transform 1 0 24552 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 25288 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_266
timestamp 1586364061
transform 1 0 25104 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_270
timestamp 1586364061
transform 1 0 25472 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_276
timestamp 1586364061
transform 1 0 26024 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26392 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 632 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 908 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2012 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3116 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3484 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 3576 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 4680 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 5784 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 6888 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 7992 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9096 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_93
timestamp 1586364061
transform 1 0 9188 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 9556 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10568 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_106
timestamp 1586364061
transform 1 0 10384 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_110
timestamp 1586364061
transform 1 0 10752 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11120 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10936 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12868 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12316 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12684 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_125
timestamp 1586364061
transform 1 0 12132 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_129
timestamp 1586364061
transform 1 0 12500 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 14524 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 13880 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_142
timestamp 1586364061
transform 1 0 13696 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_146
timestamp 1586364061
transform 1 0 14064 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_150
timestamp 1586364061
transform 1 0 14432 0 -1 9248
box -38 -48 130 592
use scs8hd_nor3_4  _168_
timestamp 1586364061
transform 1 0 14800 0 -1 9248
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 14708 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16364 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16732 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_167
timestamp 1586364061
transform 1 0 15996 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_173
timestamp 1586364061
transform 1 0 16548 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_177
timestamp 1586364061
transform 1 0 16916 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17468 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17284 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_192
timestamp 1586364061
transform 1 0 18296 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19308 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 19124 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 18480 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_196
timestamp 1586364061
transform 1 0 18664 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_200
timestamp 1586364061
transform 1 0 19032 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 19584 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20320 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 19768 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 20872 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_210
timestamp 1586364061
transform 1 0 19952 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_12_215
timestamp 1586364061
transform 1 0 20412 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_219
timestamp 1586364061
transform 1 0 20780 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21240 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_12_222
timestamp 1586364061
transform 1 0 21056 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_233
timestamp 1586364061
transform 1 0 22068 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22804 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22620 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 24368 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24000 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_250
timestamp 1586364061
transform 1 0 23632 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_256
timestamp 1586364061
transform 1 0 24184 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 25932 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_267
timestamp 1586364061
transform 1 0 25196 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26024 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26392 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 632 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 632 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 908 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 908 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2012 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3116 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2012 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3116 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3484 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4220 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 3576 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5324 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 4680 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6244 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6060 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6336 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 5784 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 6888 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7440 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 7992 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_1  _152_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9280 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9096 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9096 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 8912 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_86
timestamp 1586364061
transform 1 0 8544 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9372 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_93
timestamp 1586364061
transform 1 0 9188 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10292 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10292 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 10108 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 9740 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_99
timestamp 1586364061
transform 1 0 9740 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_97
timestamp 1586364061
transform 1 0 9556 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_101
timestamp 1586364061
transform 1 0 9924 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_116
timestamp 1586364061
transform 1 0 11304 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11120 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11304 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_120
timestamp 1586364061
transform 1 0 11672 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11488 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11672 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 11856 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 11488 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 11856 0 1 9248
box -38 -48 130 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 11948 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12040 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 13236 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 12868 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 12500 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13052 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_126
timestamp 1586364061
transform 1 0 12224 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_131
timestamp 1586364061
transform 1 0 12684 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_135
timestamp 1586364061
transform 1 0 13052 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_133
timestamp 1586364061
transform 1 0 12868 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_137
timestamp 1586364061
transform 1 0 13236 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 13604 0 -1 10336
box -38 -48 314 592
use scs8hd_nor3_4  _169_
timestamp 1586364061
transform 1 0 13420 0 1 9248
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 14524 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 14064 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 13420 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_152
timestamp 1586364061
transform 1 0 14616 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 13880 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_148
timestamp 1586364061
transform 1 0 14248 0 -1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 14800 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15352 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 14708 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 14800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 15168 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15812 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_156
timestamp 1586364061
transform 1 0 14984 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_163
timestamp 1586364061
transform 1 0 15628 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16364 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16364 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 16180 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16916 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_169
timestamp 1586364061
transform 1 0 16180 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_173
timestamp 1586364061
transform 1 0 16548 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17100 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_167
timestamp 1586364061
transform 1 0 15996 0 -1 10336
box -38 -48 222 592
use scs8hd_or4_4  _104_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18112 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17560 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17468 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 17284 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 17928 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 17560 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18388 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_182
timestamp 1586364061
transform 1 0 17376 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_186
timestamp 1586364061
transform 1 0 17744 0 -1 10336
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 19124 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 19124 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 18940 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 18572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 19492 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 18756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_199
timestamp 1586364061
transform 1 0 18940 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_203
timestamp 1586364061
transform 1 0 19308 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_207
timestamp 1586364061
transform 1 0 19676 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_211
timestamp 1586364061
transform 1 0 20044 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_214
timestamp 1586364061
transform 1 0 20320 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_210
timestamp 1586364061
transform 1 0 19952 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 19860 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 20136 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20320 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_219
timestamp 1586364061
transform 1 0 20780 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_215
timestamp 1586364061
transform 1 0 20412 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_220
timestamp 1586364061
transform 1 0 20872 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 20596 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20688 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20964 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21240 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21056 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_235
timestamp 1586364061
transform 1 0 22252 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_232
timestamp 1586364061
transform 1 0 21976 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_239
timestamp 1586364061
transform 1 0 22620 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_236
timestamp 1586364061
transform 1 0 22344 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_239
timestamp 1586364061
transform 1 0 22620 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22436 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22804 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22436 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_249
timestamp 1586364061
transform 1 0 23540 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_245
timestamp 1586364061
transform 1 0 23172 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 22988 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23356 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23080 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22988 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_246
timestamp 1586364061
transform 1 0 23264 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24000 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24092 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23908 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 25932 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25104 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25472 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_264
timestamp 1586364061
transform 1 0 24920 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_268
timestamp 1586364061
transform 1 0 25288 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_272
timestamp 1586364061
transform 1 0 25656 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26024 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 24828 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26024 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26392 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26392 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 632 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 908 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2012 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3116 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4220 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5324 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6244 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6060 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6336 0 1 10336
box -38 -48 1142 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 8268 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 8084 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_74
timestamp 1586364061
transform 1 0 7440 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_80
timestamp 1586364061
transform 1 0 7992 0 1 10336
box -38 -48 130 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 9280 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 9096 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 8728 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_86
timestamp 1586364061
transform 1 0 8544 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_90
timestamp 1586364061
transform 1 0 8912 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 10292 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 9832 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_97
timestamp 1586364061
transform 1 0 9556 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_102
timestamp 1586364061
transform 1 0 10016 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11948 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 11856 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 11304 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 11672 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11120 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11488 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 12960 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 12776 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_136
timestamp 1586364061
transform 1 0 13144 0 1 10336
box -38 -48 314 592
use scs8hd_or4_4  _143_
timestamp 1586364061
transform 1 0 13972 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 13788 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 13420 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_141
timestamp 1586364061
transform 1 0 13604 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 15536 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 15352 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 14984 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_154
timestamp 1586364061
transform 1 0 14800 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_158
timestamp 1586364061
transform 1 0 15168 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 16548 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 16916 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_171
timestamp 1586364061
transform 1 0 16364 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 16732 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17100 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 17560 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17468 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 17284 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_193
timestamp 1586364061
transform 1 0 18388 0 1 10336
box -38 -48 314 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 19124 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 18664 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_198
timestamp 1586364061
transform 1 0 18848 0 1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 20688 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 20504 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 20136 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_210
timestamp 1586364061
transform 1 0 19952 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_214
timestamp 1586364061
transform 1 0 20320 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 21700 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22160 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_227
timestamp 1586364061
transform 1 0 21516 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_231
timestamp 1586364061
transform 1 0 21884 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23172 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23080 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 22896 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22528 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22344 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 22712 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 24368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 24736 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_256
timestamp 1586364061
transform 1 0 24184 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_260
timestamp 1586364061
transform 1 0 24552 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 24920 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 25472 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_268
timestamp 1586364061
transform 1 0 25288 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_272
timestamp 1586364061
transform 1 0 25656 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26024 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26392 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 632 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 908 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2012 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3116 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3484 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 3576 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 4680 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 5784 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 6888 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 8084 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_80
timestamp 1586364061
transform 1 0 7992 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9096 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_84
timestamp 1586364061
transform 1 0 8360 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_4  FILLER_16_93
timestamp 1586364061
transform 1 0 9188 0 -1 11424
box -38 -48 406 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 9832 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 10476 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 9648 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_97
timestamp 1586364061
transform 1 0 9556 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_103
timestamp 1586364061
transform 1 0 10108 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_109
timestamp 1586364061
transform 1 0 10660 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 11028 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 10844 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 12040 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_122
timestamp 1586364061
transform 1 0 11856 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 12592 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 12408 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_126
timestamp 1586364061
transform 1 0 12224 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 13972 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 13604 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 14340 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_139
timestamp 1586364061
transform 1 0 13420 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_143
timestamp 1586364061
transform 1 0 13788 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_147
timestamp 1586364061
transform 1 0 14156 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14524 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 14800 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 14708 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_163
timestamp 1586364061
transform 1 0 15628 0 -1 11424
box -38 -48 590 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 16364 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16180 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 18112 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 17744 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 17376 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_180
timestamp 1586364061
transform 1 0 17192 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_184
timestamp 1586364061
transform 1 0 17560 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_188
timestamp 1586364061
transform 1 0 17928 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_192
timestamp 1586364061
transform 1 0 18296 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 18664 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 18480 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 19676 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_205
timestamp 1586364061
transform 1 0 19492 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 20412 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20320 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_209
timestamp 1586364061
transform 1 0 19860 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20228 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 21424 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21792 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22160 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_224
timestamp 1586364061
transform 1 0 21240 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_228
timestamp 1586364061
transform 1 0 21608 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_232
timestamp 1586364061
transform 1 0 21976 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22436 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23448 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_236
timestamp 1586364061
transform 1 0 22344 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_246
timestamp 1586364061
transform 1 0 23264 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 24000 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_4  FILLER_16_250
timestamp 1586364061
transform 1 0 23632 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 25932 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 24828 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26024 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26392 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 632 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 908 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2012 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3116 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4220 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5324 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6244 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6060 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_62
timestamp 1586364061
transform 1 0 6336 0 1 11424
box -38 -48 774 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 7164 0 1 11424
box -38 -48 314 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 8176 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 7624 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_70
timestamp 1586364061
transform 1 0 7072 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_74
timestamp 1586364061
transform 1 0 7440 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_78
timestamp 1586364061
transform 1 0 7808 0 1 11424
box -38 -48 406 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 9188 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 8636 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 9004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_85
timestamp 1586364061
transform 1 0 8452 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_89
timestamp 1586364061
transform 1 0 8820 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_96
timestamp 1586364061
transform 1 0 9464 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 10200 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 9648 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 10016 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_100
timestamp 1586364061
transform 1 0 9832 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 11948 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 11856 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 11212 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 11672 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_113
timestamp 1586364061
transform 1 0 11028 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_117
timestamp 1586364061
transform 1 0 11396 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 13144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_132
timestamp 1586364061
transform 1 0 12776 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_17_138
timestamp 1586364061
transform 1 0 13328 0 1 11424
box -38 -48 314 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 13788 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 13604 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_152
timestamp 1586364061
transform 1 0 14616 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 15352 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 14800 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 15168 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_156
timestamp 1586364061
transform 1 0 14984 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16364 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16732 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_169
timestamp 1586364061
transform 1 0 16180 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_173
timestamp 1586364061
transform 1 0 16548 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_177
timestamp 1586364061
transform 1 0 16916 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17652 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17468 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 18112 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 17284 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_184
timestamp 1586364061
transform 1 0 17560 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_188
timestamp 1586364061
transform 1 0 17928 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_192
timestamp 1586364061
transform 1 0 18296 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 18664 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 18480 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 19676 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_205
timestamp 1586364061
transform 1 0 19492 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20320 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20780 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20136 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_209
timestamp 1586364061
transform 1 0 19860 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_217
timestamp 1586364061
transform 1 0 20596 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_221
timestamp 1586364061
transform 1 0 20964 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21332 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21148 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23264 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23080 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22528 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22344 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 22712 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_245
timestamp 1586364061
transform 1 0 23172 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24276 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24644 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_255
timestamp 1586364061
transform 1 0 24092 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_259
timestamp 1586364061
transform 1 0 24460 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 24828 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 25380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_267
timestamp 1586364061
transform 1 0 25196 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_271
timestamp 1586364061
transform 1 0 25564 0 1 11424
box -38 -48 590 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26392 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 632 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 908 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2012 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3116 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3484 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 3576 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 4680 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 5784 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 6888 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 8084 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_80
timestamp 1586364061
transform 1 0 7992 0 -1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9096 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_84
timestamp 1586364061
transform 1 0 8360 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_6  FILLER_18_93
timestamp 1586364061
transform 1 0 9188 0 -1 12512
box -38 -48 590 592
use scs8hd_buf_1  _139_
timestamp 1586364061
transform 1 0 10016 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 10476 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 9832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_99
timestamp 1586364061
transform 1 0 9740 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_105
timestamp 1586364061
transform 1 0 10292 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_109
timestamp 1586364061
transform 1 0 10660 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _157_
timestamp 1586364061
transform 1 0 11028 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 12040 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 10844 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_122
timestamp 1586364061
transform 1 0 11856 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 13144 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 12960 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 12408 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_126
timestamp 1586364061
transform 1 0 12224 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_130
timestamp 1586364061
transform 1 0 12592 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 14156 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 14524 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 13972 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14340 0 -1 12512
box -38 -48 222 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 15260 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 14708 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 15720 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_154
timestamp 1586364061
transform 1 0 14800 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_158
timestamp 1586364061
transform 1 0 15168 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_162
timestamp 1586364061
transform 1 0 15536 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_166
timestamp 1586364061
transform 1 0 15904 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16272 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16088 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_179
timestamp 1586364061
transform 1 0 17100 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 18296 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 18112 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 17744 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17284 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_183
timestamp 1586364061
transform 1 0 17468 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_188
timestamp 1586364061
transform 1 0 17928 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 19308 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 19676 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_201
timestamp 1586364061
transform 1 0 19124 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_205
timestamp 1586364061
transform 1 0 19492 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20320 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 20688 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20136 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_209
timestamp 1586364061
transform 1 0 19860 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_215
timestamp 1586364061
transform 1 0 20412 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_220
timestamp 1586364061
transform 1 0 20872 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21332 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 21056 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_224
timestamp 1586364061
transform 1 0 21240 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23264 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22528 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_236
timestamp 1586364061
transform 1 0 22344 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_240
timestamp 1586364061
transform 1 0 22712 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_8  FILLER_18_255
timestamp 1586364061
transform 1 0 24092 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24828 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 25932 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_266
timestamp 1586364061
transform 1 0 25104 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_274
timestamp 1586364061
transform 1 0 25840 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26024 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26392 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 632 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 632 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 908 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 908 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2012 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3116 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2012 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3116 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3484 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4220 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 3576 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5324 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 4680 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6244 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6060 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6336 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 5784 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 6888 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7440 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 7992 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 9280 0 1 12512
box -38 -48 314 592
use scs8hd_nand2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9372 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9096 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 9096 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_86
timestamp 1586364061
transform 1 0 8544 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9188 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 10292 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 9740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 10108 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 10384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 10752 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_97
timestamp 1586364061
transform 1 0 9556 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_101
timestamp 1586364061
transform 1 0 9924 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_104
timestamp 1586364061
transform 1 0 10200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_108
timestamp 1586364061
transform 1 0 10568 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 11948 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 11212 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 11856 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 11672 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 11304 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11120 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11488 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_112
timestamp 1586364061
transform 1 0 10936 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_124
timestamp 1586364061
transform 1 0 12040 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 12776 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 12960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 12316 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 12776 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_136
timestamp 1586364061
transform 1 0 13144 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_129
timestamp 1586364061
transform 1 0 12500 0 -1 13600
box -38 -48 314 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 13788 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 13604 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 13788 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 14156 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_140
timestamp 1586364061
transform 1 0 13512 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_152
timestamp 1586364061
transform 1 0 14616 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_141
timestamp 1586364061
transform 1 0 13604 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 13972 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_149
timestamp 1586364061
transform 1 0 14340 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_158
timestamp 1586364061
transform 1 0 15168 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 14800 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_156
timestamp 1586364061
transform 1 0 14984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14984 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 14800 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15168 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 14708 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_160
timestamp 1586364061
transform 1 0 15352 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15352 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15536 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15720 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15536 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16916 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17100 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 16732 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17100 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_173
timestamp 1586364061
transform 1 0 16548 0 -1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17284 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17560 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17468 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17284 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_193
timestamp 1586364061
transform 1 0 18388 0 1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_20_190
timestamp 1586364061
transform 1 0 18112 0 -1 13600
box -38 -48 590 592
use scs8hd_or2_4  _099_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18848 0 -1 13600
box -38 -48 682 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 19124 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 18848 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 19676 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 18664 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_197
timestamp 1586364061
transform 1 0 18756 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_200
timestamp 1586364061
transform 1 0 19032 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_205
timestamp 1586364061
transform 1 0 19492 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 20688 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20412 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20320 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20412 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_210
timestamp 1586364061
transform 1 0 19952 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_214
timestamp 1586364061
transform 1 0 20320 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_217
timestamp 1586364061
transform 1 0 20596 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_209
timestamp 1586364061
transform 1 0 19860 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_213
timestamp 1586364061
transform 1 0 20228 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 21700 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 21424 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22160 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_227
timestamp 1586364061
transform 1 0 21516 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_231
timestamp 1586364061
transform 1 0 21884 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_235
timestamp 1586364061
transform 1 0 22252 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_224
timestamp 1586364061
transform 1 0 21240 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_228
timestamp 1586364061
transform 1 0 21608 0 -1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23172 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22344 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23080 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22344 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22896 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23356 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_238
timestamp 1586364061
transform 1 0 22528 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_245
timestamp 1586364061
transform 1 0 23172 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_249
timestamp 1586364061
transform 1 0 23540 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 23908 0 -1 13600
box -38 -48 866 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 24736 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 24184 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_254
timestamp 1586364061
transform 1 0 24000 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_258
timestamp 1586364061
transform 1 0 24368 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_262
timestamp 1586364061
transform 1 0 24736 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 25932 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 25288 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_266
timestamp 1586364061
transform 1 0 25104 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_270
timestamp 1586364061
transform 1 0 25472 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_276
timestamp 1586364061
transform 1 0 26024 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 25840 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26024 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26392 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26392 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 632 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 908 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2012 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3116 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4220 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5324 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6244 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6060 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6336 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7440 0 1 13600
box -38 -48 1142 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 9096 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 8912 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_86
timestamp 1586364061
transform 1 0 8544 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 10108 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 10476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_101
timestamp 1586364061
transform 1 0 9924 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_105
timestamp 1586364061
transform 1 0 10292 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_109
timestamp 1586364061
transform 1 0 10660 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 10844 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 11856 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 11304 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 11672 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11120 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11488 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 11948 0 1 13600
box -38 -48 222 592
use scs8hd_nand2_4  _138_
timestamp 1586364061
transform 1 0 12316 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 12132 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 13328 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_136
timestamp 1586364061
transform 1 0 13144 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 14616 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 14432 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 14064 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 13696 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_140
timestamp 1586364061
transform 1 0 13512 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_144
timestamp 1586364061
transform 1 0 13880 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_148
timestamp 1586364061
transform 1 0 14248 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15628 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_161
timestamp 1586364061
transform 1 0 15444 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_165
timestamp 1586364061
transform 1 0 15812 0 1 13600
box -38 -48 406 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 16456 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 16916 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 16272 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_169
timestamp 1586364061
transform 1 0 16180 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 16732 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17100 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17560 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17468 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17284 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_193
timestamp 1586364061
transform 1 0 18388 0 1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19308 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19124 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 18756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_199
timestamp 1586364061
transform 1 0 18940 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20504 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20872 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_214
timestamp 1586364061
transform 1 0 20320 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_218
timestamp 1586364061
transform 1 0 20688 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21516 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21332 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_222
timestamp 1586364061
transform 1 0 21056 0 1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 23172 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23080 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22528 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 22896 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22344 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 22712 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 24736 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 24184 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_254
timestamp 1586364061
transform 1 0 24000 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_258
timestamp 1586364061
transform 1 0 24368 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 25288 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_266
timestamp 1586364061
transform 1 0 25104 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_270
timestamp 1586364061
transform 1 0 25472 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_276
timestamp 1586364061
transform 1 0 26024 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26392 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 632 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 908 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2012 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3116 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3484 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 3576 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 4680 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 5784 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 6888 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 7992 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9096 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_93
timestamp 1586364061
transform 1 0 9188 0 -1 14688
box -38 -48 406 592
use scs8hd_or2_4  _102_
timestamp 1586364061
transform 1 0 9648 0 -1 14688
box -38 -48 682 592
use scs8hd_fill_1  FILLER_22_97
timestamp 1586364061
transform 1 0 9556 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10292 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 11764 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_117
timestamp 1586364061
transform 1 0 11396 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_124
timestamp 1586364061
transform 1 0 12040 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 13144 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 12868 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_132
timestamp 1586364061
transform 1 0 12776 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_135
timestamp 1586364061
transform 1 0 13052 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_145
timestamp 1586364061
transform 1 0 13972 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14800 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 14708 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_163
timestamp 1586364061
transform 1 0 15628 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 16364 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17376 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17744 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_180
timestamp 1586364061
transform 1 0 17192 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_184
timestamp 1586364061
transform 1 0 17560 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_188
timestamp 1586364061
transform 1 0 17928 0 -1 14688
box -38 -48 590 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 18756 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 18480 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_196
timestamp 1586364061
transform 1 0 18664 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_206
timestamp 1586364061
transform 1 0 19584 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20412 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20320 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19768 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20136 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_210
timestamp 1586364061
transform 1 0 19952 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22160 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21608 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_226
timestamp 1586364061
transform 1 0 21424 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_230
timestamp 1586364061
transform 1 0 21792 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 23172 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_243
timestamp 1586364061
transform 1 0 22988 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_247
timestamp 1586364061
transform 1 0 23356 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 23724 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_260
timestamp 1586364061
transform 1 0 24552 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 25932 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_272
timestamp 1586364061
transform 1 0 25656 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26024 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26392 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 632 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 908 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2012 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3116 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4220 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5324 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6244 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6060 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6336 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7440 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 8544 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 9648 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 10752 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 11856 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 11948 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 13144 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 12868 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 12500 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 12132 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_127
timestamp 1586364061
transform 1 0 12316 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_131
timestamp 1586364061
transform 1 0 12684 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_135
timestamp 1586364061
transform 1 0 13052 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14524 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 14156 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_145
timestamp 1586364061
transform 1 0 13972 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_149
timestamp 1586364061
transform 1 0 14340 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14708 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15904 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_164
timestamp 1586364061
transform 1 0 15720 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 16456 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17008 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16272 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_168
timestamp 1586364061
transform 1 0 16088 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_175
timestamp 1586364061
transform 1 0 16732 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17468 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 18296 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 17928 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_180
timestamp 1586364061
transform 1 0 17192 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_184
timestamp 1586364061
transform 1 0 17560 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_190
timestamp 1586364061
transform 1 0 18112 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 18480 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 19492 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_203
timestamp 1586364061
transform 1 0 19308 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_207
timestamp 1586364061
transform 1 0 19676 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20688 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20412 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20044 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_213
timestamp 1586364061
transform 1 0 20228 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_217
timestamp 1586364061
transform 1 0 20596 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22160 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21700 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_227
timestamp 1586364061
transform 1 0 21516 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_231
timestamp 1586364061
transform 1 0 21884 0 1 14688
box -38 -48 314 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 23172 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23080 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22528 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 22896 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_236
timestamp 1586364061
transform 1 0 22344 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_240
timestamp 1586364061
transform 1 0 22712 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24736 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 24184 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_254
timestamp 1586364061
transform 1 0 24000 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_258
timestamp 1586364061
transform 1 0 24368 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25196 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_265
timestamp 1586364061
transform 1 0 25012 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25380 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26392 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 632 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 908 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2012 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3116 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3484 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 3576 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 4680 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 5784 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 6888 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 7992 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9096 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9188 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10292 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11396 0 -1 15776
box -38 -48 1142 592
use scs8hd_or4_4  _166_
timestamp 1586364061
transform 1 0 12868 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_4  FILLER_24_129
timestamp 1586364061
transform 1 0 12500 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 13880 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_142
timestamp 1586364061
transform 1 0 13696 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_146
timestamp 1586364061
transform 1 0 14064 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 14616 0 -1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15260 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 14708 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14984 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_154
timestamp 1586364061
transform 1 0 14800 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_158
timestamp 1586364061
transform 1 0 15168 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17008 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_170
timestamp 1586364061
transform 1 0 16272 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_8  FILLER_24_187
timestamp 1586364061
transform 1 0 17836 0 -1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 18756 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_24_195
timestamp 1586364061
transform 1 0 18572 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_206
timestamp 1586364061
transform 1 0 19584 0 -1 15776
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20412 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20320 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20136 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22160 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21608 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_226
timestamp 1586364061
transform 1 0 21424 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_230
timestamp 1586364061
transform 1 0 21792 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_243
timestamp 1586364061
transform 1 0 22988 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 23724 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_260
timestamp 1586364061
transform 1 0 24552 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 25932 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_272
timestamp 1586364061
transform 1 0 25656 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26024 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26392 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 632 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 908 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2012 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3116 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4220 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5324 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6244 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6060 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6336 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7440 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 8544 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 9648 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 10752 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 11856 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 11948 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13052 0 1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 14524 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_147
timestamp 1586364061
transform 1 0 14156 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15536 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15352 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 14984 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_154
timestamp 1586364061
transform 1 0 14800 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15168 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16548 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16916 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_171
timestamp 1586364061
transform 1 0 16364 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 16732 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17100 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 17560 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17468 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 17284 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18388 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19492 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19308 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 18572 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_197
timestamp 1586364061
transform 1 0 18756 0 1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20688 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_216
timestamp 1586364061
transform 1 0 20504 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_220
timestamp 1586364061
transform 1 0 20872 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21516 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21332 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_224
timestamp 1586364061
transform 1 0 21240 0 1 15776
box -38 -48 130 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 23172 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23080 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 22528 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 22896 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22344 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 22712 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 24736 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24184 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_254
timestamp 1586364061
transform 1 0 24000 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_258
timestamp 1586364061
transform 1 0 24368 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25196 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_265
timestamp 1586364061
transform 1 0 25012 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25380 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26392 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 632 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 632 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 908 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 908 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2012 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3116 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2012 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3116 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3484 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 3576 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4220 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 4680 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5324 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6244 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 5784 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 6888 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6060 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6336 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 7992 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7440 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9096 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9188 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 8544 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10292 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 9648 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 10752 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 11856 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11396 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 11948 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12500 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13052 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 13604 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14156 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 15812 0 1 16864
box -38 -48 866 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 14892 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 14708 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 15628 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15904 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_154
timestamp 1586364061
transform 1 0 14800 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_164
timestamp 1586364061
transform 1 0 15720 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_159
timestamp 1586364061
transform 1 0 15260 0 1 16864
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16456 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_26_168
timestamp 1586364061
transform 1 0 16088 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_27_174
timestamp 1586364061
transform 1 0 16640 0 1 16864
box -38 -48 774 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 18204 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17468 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_181
timestamp 1586364061
transform 1 0 17284 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_189
timestamp 1586364061
transform 1 0 18020 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_182
timestamp 1586364061
transform 1 0 17376 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 17560 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 19584 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19492 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 19400 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_194
timestamp 1586364061
transform 1 0 18480 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_202
timestamp 1586364061
transform 1 0 19216 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_26_207
timestamp 1586364061
transform 1 0 19676 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_8  FILLER_27_196
timestamp 1586364061
transform 1 0 18664 0 1 16864
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20596 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20320 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20964 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 20596 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20228 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_215
timestamp 1586364061
transform 1 0 20412 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_215
timestamp 1586364061
transform 1 0 20412 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_219
timestamp 1586364061
transform 1 0 20780 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 22160 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21148 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 22160 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_226
timestamp 1586364061
transform 1 0 21424 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_232
timestamp 1586364061
transform 1 0 21976 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23080 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_243
timestamp 1586364061
transform 1 0 22988 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_27_236
timestamp 1586364061
transform 1 0 22344 0 1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_245
timestamp 1586364061
transform 1 0 23172 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_249
timestamp 1586364061
transform 1 0 23540 0 1 16864
box -38 -48 130 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 23632 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24644 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24736 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23724 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24092 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_254
timestamp 1586364061
transform 1 0 24000 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_253
timestamp 1586364061
transform 1 0 23908 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_257
timestamp 1586364061
transform 1 0 24276 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 25932 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25104 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_265
timestamp 1586364061
transform 1 0 25012 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_273
timestamp 1586364061
transform 1 0 25748 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26024 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_264
timestamp 1586364061
transform 1 0 24920 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_268
timestamp 1586364061
transform 1 0 25288 0 1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26024 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26392 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26392 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 632 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 908 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2012 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3116 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3484 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 3576 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 4680 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 5784 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 6888 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 7992 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9096 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9188 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10292 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11396 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12500 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 13604 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 14708 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 14800 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 15904 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17008 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18112 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19216 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 20412 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20320 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 21976 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21424 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_224
timestamp 1586364061
transform 1 0 21240 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_228
timestamp 1586364061
transform 1 0 21608 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_241
timestamp 1586364061
transform 1 0 22804 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_253
timestamp 1586364061
transform 1 0 23908 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_258
timestamp 1586364061
transform 1 0 24368 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 25932 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_270
timestamp 1586364061
transform 1 0 25472 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_274
timestamp 1586364061
transform 1 0 25840 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26024 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26392 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 632 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 908 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2012 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3116 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4220 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5324 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6244 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6060 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6336 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7440 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 8544 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 9648 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 10752 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 11856 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 11948 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13052 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14156 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15260 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16364 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17468 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 17560 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 18664 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20412 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_208
timestamp 1586364061
transform 1 0 19768 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_214
timestamp 1586364061
transform 1 0 20320 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_217
timestamp 1586364061
transform 1 0 20596 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22068 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_229
timestamp 1586364061
transform 1 0 21700 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23080 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23356 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22528 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_236
timestamp 1586364061
transform 1 0 22344 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_240
timestamp 1586364061
transform 1 0 22712 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_245
timestamp 1586364061
transform 1 0 23172 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_249
timestamp 1586364061
transform 1 0 23540 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24552 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_258
timestamp 1586364061
transform 1 0 24368 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_262
timestamp 1586364061
transform 1 0 24736 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25564 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24920 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_269
timestamp 1586364061
transform 1 0 25380 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_273
timestamp 1586364061
transform 1 0 25748 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26392 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 632 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 908 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2012 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3116 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3484 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 3576 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 4680 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 5784 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 6888 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 7992 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9096 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9188 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10292 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11396 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12500 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 13604 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 14708 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 14800 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 15904 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17008 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18112 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19216 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20412 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20320 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_218
timestamp 1586364061
transform 1 0 20688 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_230
timestamp 1586364061
transform 1 0 21792 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23080 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_242
timestamp 1586364061
transform 1 0 22896 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_247
timestamp 1586364061
transform 1 0 23356 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_258
timestamp 1586364061
transform 1 0 24368 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 25932 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_270
timestamp 1586364061
transform 1 0 25472 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_274
timestamp 1586364061
transform 1 0 25840 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26024 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26392 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 632 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 908 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2012 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3116 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4220 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5324 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6244 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6060 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6336 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7440 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 8544 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 9648 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 10752 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 11856 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 11948 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13052 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14156 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15260 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16364 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17468 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 17560 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 18664 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 19768 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 20872 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 21976 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23080 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23172 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24552 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 23908 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_258
timestamp 1586364061
transform 1 0 24368 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_262
timestamp 1586364061
transform 1 0 24736 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24920 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_266
timestamp 1586364061
transform 1 0 25104 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_274
timestamp 1586364061
transform 1 0 25840 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26392 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 632 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 908 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2012 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3116 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3484 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 3576 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 4680 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 5784 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 6888 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 7992 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9096 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9188 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10292 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11396 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12500 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 13604 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 14708 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 14800 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 15904 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17008 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18112 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19216 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20320 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20412 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21516 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 22620 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_251
timestamp 1586364061
transform 1 0 23724 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_258
timestamp 1586364061
transform 1 0 24368 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 25932 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_270
timestamp 1586364061
transform 1 0 25472 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_274
timestamp 1586364061
transform 1 0 25840 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26024 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26392 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 632 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 632 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 908 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 908 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2012 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3116 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2012 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3116 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3484 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4220 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 3576 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5324 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 4680 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6244 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6060 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6336 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 5784 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 6888 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7440 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 7992 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9096 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 8544 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9188 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 9648 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 10752 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10292 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 11856 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 11948 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11396 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13052 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12500 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14156 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 13604 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 14708 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15260 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 14800 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 15904 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16364 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17008 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17468 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 17560 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18112 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 18664 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19216 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20320 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 19768 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 20872 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20412 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 21976 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21516 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23080 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23172 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 22620 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24092 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 23908 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24276 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_251
timestamp 1586364061
transform 1 0 23724 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_258
timestamp 1586364061
transform 1 0 24368 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 25932 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25380 0 1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_270
timestamp 1586364061
transform 1 0 25472 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 25840 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26024 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26392 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26392 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 632 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 908 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2012 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3116 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4220 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5324 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6244 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6060 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6336 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7440 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 8544 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 9648 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 10752 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 11856 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 11948 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13052 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14156 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15260 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16364 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17468 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 17560 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 18664 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 19768 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 20872 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 21976 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23080 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23172 0 1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24552 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_253
timestamp 1586364061
transform 1 0 23908 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_258
timestamp 1586364061
transform 1 0 24368 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_262
timestamp 1586364061
transform 1 0 24736 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_35_274
timestamp 1586364061
transform 1 0 25840 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26392 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 632 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 908 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2012 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3116 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3484 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 3576 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 4680 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 5784 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 6888 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 7992 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9096 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9188 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10292 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11396 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12500 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 13604 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 14708 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 14800 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 15904 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17008 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18112 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19216 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20320 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20412 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21516 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 22620 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 23724 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 25932 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 24828 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26024 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26392 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 632 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 908 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2012 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3116 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4220 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5324 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6244 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6060 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6336 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7440 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 8544 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 9648 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 10752 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 11856 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 11948 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13052 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14156 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15260 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16364 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17468 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 17560 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 18664 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 19768 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 20872 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 21976 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23080 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23172 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24276 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25380 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26392 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 632 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 908 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2012 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3116 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3484 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 3576 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 4680 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 5784 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 6888 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 7992 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9096 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9188 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10292 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11396 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12500 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 13604 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 14708 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 14800 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 15904 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17008 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18112 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19216 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20320 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20412 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21516 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 22620 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 23724 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 25932 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 24828 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26024 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26392 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 632 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 632 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 908 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 908 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2012 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3116 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2012 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3116 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3484 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4220 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 3576 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5324 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 4680 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6244 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6060 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6336 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 5784 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 6888 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7440 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 7992 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9096 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 8544 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9188 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 9648 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 10752 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10292 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 11856 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 11948 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11396 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13052 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12500 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14156 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 13604 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 14708 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15260 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 14800 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 15904 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16364 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17008 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17468 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 17560 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18112 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 18664 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19216 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20320 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 19768 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_39_220
timestamp 1586364061
transform 1 0 20872 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20412 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21148 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21608 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_226
timestamp 1586364061
transform 1 0 21424 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_230
timestamp 1586364061
transform 1 0 21792 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21516 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23080 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_242
timestamp 1586364061
transform 1 0 22896 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23172 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 22620 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24092 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24552 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 23908 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_258
timestamp 1586364061
transform 1 0 24368 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_262
timestamp 1586364061
transform 1 0 24736 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 23724 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 25932 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_274
timestamp 1586364061
transform 1 0 25840 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 24828 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26024 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26392 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26392 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 632 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 908 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2012 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3116 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4220 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5324 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6244 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6060 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6336 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7440 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 8544 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 9648 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 10752 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 11856 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 11948 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13052 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14156 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15260 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16364 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17468 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 17560 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 18664 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 19768 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 20872 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 21976 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23080 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23172 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24276 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25380 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26392 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 632 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 908 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3116 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3484 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 3576 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 4680 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6336 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 5784 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6428 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 7532 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9188 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 8636 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9280 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10384 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12040 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11488 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12132 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13236 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14340 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 14892 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 14984 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16088 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 17744 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17192 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 17836 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 18940 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 20596 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20044 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 20688 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 21792 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23448 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 22896 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 23540 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 24644 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 25748 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26392 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 4790 27520 4846 28000 6 address[0]
port 0 nsew default input
rlabel metal2 s 8286 27520 8342 28000 6 address[1]
port 1 nsew default input
rlabel metal2 s 11782 27520 11838 28000 6 address[2]
port 2 nsew default input
rlabel metal2 s 15278 27520 15334 28000 6 address[3]
port 3 nsew default input
rlabel metal2 s 18774 27520 18830 28000 6 address[4]
port 4 nsew default input
rlabel metal2 s 22270 27520 22326 28000 6 address[5]
port 5 nsew default input
rlabel metal2 s 5158 0 5214 480 6 bottom_left_grid_pin_11_
port 6 nsew default input
rlabel metal2 s 6170 0 6226 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 7182 0 7238 480 6 bottom_left_grid_pin_15_
port 8 nsew default input
rlabel metal2 s 6 0 62 480 6 bottom_left_grid_pin_1_
port 9 nsew default input
rlabel metal2 s 1018 0 1074 480 6 bottom_left_grid_pin_3_
port 10 nsew default input
rlabel metal2 s 2030 0 2086 480 6 bottom_left_grid_pin_5_
port 11 nsew default input
rlabel metal2 s 3042 0 3098 480 6 bottom_left_grid_pin_7_
port 12 nsew default input
rlabel metal2 s 4146 0 4202 480 6 bottom_left_grid_pin_9_
port 13 nsew default input
rlabel metal2 s 26870 0 26926 480 6 bottom_right_grid_pin_11_
port 14 nsew default input
rlabel metal3 s 27048 10752 27528 10872 6 chanx_right_in[0]
port 15 nsew default input
rlabel metal3 s 27048 11704 27528 11824 6 chanx_right_in[1]
port 16 nsew default input
rlabel metal3 s 27048 12792 27528 12912 6 chanx_right_in[2]
port 17 nsew default input
rlabel metal3 s 27048 13880 27528 14000 6 chanx_right_in[3]
port 18 nsew default input
rlabel metal3 s 27048 14832 27528 14952 6 chanx_right_in[4]
port 19 nsew default input
rlabel metal3 s 27048 15920 27528 16040 6 chanx_right_in[5]
port 20 nsew default input
rlabel metal3 s 27048 17008 27528 17128 6 chanx_right_in[6]
port 21 nsew default input
rlabel metal3 s 27048 17960 27528 18080 6 chanx_right_in[7]
port 22 nsew default input
rlabel metal3 s 27048 19048 27528 19168 6 chanx_right_in[8]
port 23 nsew default input
rlabel metal3 s 27048 1368 27528 1488 6 chanx_right_out[0]
port 24 nsew default tristate
rlabel metal3 s 27048 2456 27528 2576 6 chanx_right_out[1]
port 25 nsew default tristate
rlabel metal3 s 27048 3408 27528 3528 6 chanx_right_out[2]
port 26 nsew default tristate
rlabel metal3 s 27048 4496 27528 4616 6 chanx_right_out[3]
port 27 nsew default tristate
rlabel metal3 s 27048 5584 27528 5704 6 chanx_right_out[4]
port 28 nsew default tristate
rlabel metal3 s 27048 6536 27528 6656 6 chanx_right_out[5]
port 29 nsew default tristate
rlabel metal3 s 27048 7624 27528 7744 6 chanx_right_out[6]
port 30 nsew default tristate
rlabel metal3 s 27048 8712 27528 8832 6 chanx_right_out[7]
port 31 nsew default tristate
rlabel metal3 s 27048 9664 27528 9784 6 chanx_right_out[8]
port 32 nsew default tristate
rlabel metal2 s 8286 0 8342 480 6 chany_bottom_in[0]
port 33 nsew default input
rlabel metal2 s 9298 0 9354 480 6 chany_bottom_in[1]
port 34 nsew default input
rlabel metal2 s 10310 0 10366 480 6 chany_bottom_in[2]
port 35 nsew default input
rlabel metal2 s 11322 0 11378 480 6 chany_bottom_in[3]
port 36 nsew default input
rlabel metal2 s 12426 0 12482 480 6 chany_bottom_in[4]
port 37 nsew default input
rlabel metal2 s 13438 0 13494 480 6 chany_bottom_in[5]
port 38 nsew default input
rlabel metal2 s 14450 0 14506 480 6 chany_bottom_in[6]
port 39 nsew default input
rlabel metal2 s 15462 0 15518 480 6 chany_bottom_in[7]
port 40 nsew default input
rlabel metal2 s 16566 0 16622 480 6 chany_bottom_in[8]
port 41 nsew default input
rlabel metal2 s 17578 0 17634 480 6 chany_bottom_out[0]
port 42 nsew default tristate
rlabel metal2 s 18590 0 18646 480 6 chany_bottom_out[1]
port 43 nsew default tristate
rlabel metal2 s 19602 0 19658 480 6 chany_bottom_out[2]
port 44 nsew default tristate
rlabel metal2 s 20706 0 20762 480 6 chany_bottom_out[3]
port 45 nsew default tristate
rlabel metal2 s 21718 0 21774 480 6 chany_bottom_out[4]
port 46 nsew default tristate
rlabel metal2 s 22730 0 22786 480 6 chany_bottom_out[5]
port 47 nsew default tristate
rlabel metal2 s 23742 0 23798 480 6 chany_bottom_out[6]
port 48 nsew default tristate
rlabel metal2 s 24846 0 24902 480 6 chany_bottom_out[7]
port 49 nsew default tristate
rlabel metal2 s 25858 0 25914 480 6 chany_bottom_out[8]
port 50 nsew default tristate
rlabel metal2 s 25766 27520 25822 28000 6 data_in
port 51 nsew default input
rlabel metal2 s 1294 27520 1350 28000 6 enable
port 52 nsew default input
rlabel metal3 s 27048 416 27528 536 6 right_bottom_grid_pin_12_
port 53 nsew default input
rlabel metal3 s 27048 25304 27528 25424 6 right_top_grid_pin_11_
port 54 nsew default input
rlabel metal3 s 27048 26256 27528 26376 6 right_top_grid_pin_13_
port 55 nsew default input
rlabel metal3 s 27048 27344 27528 27464 6 right_top_grid_pin_15_
port 56 nsew default input
rlabel metal3 s 27048 20000 27528 20120 6 right_top_grid_pin_1_
port 57 nsew default input
rlabel metal3 s 27048 21088 27528 21208 6 right_top_grid_pin_3_
port 58 nsew default input
rlabel metal3 s 27048 22176 27528 22296 6 right_top_grid_pin_5_
port 59 nsew default input
rlabel metal3 s 27048 23128 27528 23248 6 right_top_grid_pin_7_
port 60 nsew default input
rlabel metal3 s 27048 24216 27528 24336 6 right_top_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 5139 2128 5459 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 9805 2128 10125 25616 6 vgnd
port 63 nsew default input
<< properties >>
string FIXED_BBOX 1 0 27528 28000
<< end >>
