VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__0_
  CLASS BLOCK ;
  FOREIGN sb_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 2.400 36.000 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.400 41.440 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 2.400 44.840 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 2.400 47.560 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 2.400 50.280 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 2.400 53.000 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 2.400 55.720 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 2.400 10.160 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 2.400 16.280 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.400 19.000 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 2.400 24.440 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 2.400 27.160 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 2.400 30.560 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 2.400 61.840 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.400 90.400 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.400 93.120 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 2.400 98.560 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 2.400 101.960 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 2.400 104.680 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 2.400 107.400 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 2.400 110.120 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 2.400 112.840 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.400 116.240 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 2.400 67.280 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 2.400 76.120 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.400 78.840 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 2.400 81.560 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 2.400 84.280 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 2.400 87.680 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 4.120 140.000 4.720 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 32.680 140.000 33.280 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 35.400 140.000 36.000 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 38.120 140.000 38.720 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 40.840 140.000 41.440 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.240 140.000 44.840 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 46.960 140.000 47.560 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 49.680 140.000 50.280 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 52.400 140.000 53.000 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 55.120 140.000 55.720 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 58.520 140.000 59.120 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 6.840 140.000 7.440 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 9.560 140.000 10.160 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 12.280 140.000 12.880 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 15.680 140.000 16.280 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 18.400 140.000 19.000 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 21.120 140.000 21.720 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 23.840 140.000 24.440 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 26.560 140.000 27.160 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 29.960 140.000 30.560 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 61.240 140.000 61.840 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 89.800 140.000 90.400 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 92.520 140.000 93.120 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 95.240 140.000 95.840 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 97.960 140.000 98.560 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 101.360 140.000 101.960 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 104.080 140.000 104.680 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 106.800 140.000 107.400 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 109.520 140.000 110.120 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 112.240 140.000 112.840 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 115.640 140.000 116.240 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 63.960 140.000 64.560 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 66.680 140.000 67.280 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 72.800 140.000 73.400 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 75.520 140.000 76.120 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 78.240 140.000 78.840 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 80.960 140.000 81.560 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 83.680 140.000 84.280 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 87.080 140.000 87.680 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.470 137.600 24.750 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.910 137.600 54.190 140.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 137.600 56.950 140.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 137.600 59.710 140.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 137.600 62.930 140.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 137.600 65.690 140.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 137.600 68.450 140.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.390 137.600 71.670 140.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.150 137.600 74.430 140.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 137.600 77.190 140.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 137.600 80.410 140.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.690 137.600 27.970 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 137.600 30.730 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 137.600 33.490 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 137.600 36.710 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.190 137.600 39.470 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 137.600 42.230 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 137.600 45.450 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.930 137.600 48.210 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 137.600 50.970 140.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 137.600 83.170 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.870 137.600 112.150 140.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.090 137.600 115.370 140.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.850 137.600 118.130 140.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 137.600 120.890 140.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.830 137.600 124.110 140.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.590 137.600 126.870 140.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.350 137.600 129.630 140.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 137.600 132.850 140.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 137.600 135.610 140.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.090 137.600 138.370 140.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.650 137.600 85.930 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.870 137.600 89.150 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.630 137.600 91.910 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.390 137.600 94.670 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.610 137.600 97.890 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 137.600 100.650 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.130 137.600 103.410 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.350 137.600 106.630 140.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.110 137.600 109.390 140.000 ;
    END
  END chany_top_out[9]
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 2.400 2.000 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_top_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 2.400 118.960 ;
    END
  END left_top_grid_pin_42_
  PIN left_top_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 2.400 121.680 ;
    END
  END left_top_grid_pin_43_
  PIN left_top_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 2.400 124.400 ;
    END
  END left_top_grid_pin_44_
  PIN left_top_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.400 127.120 ;
    END
  END left_top_grid_pin_45_
  PIN left_top_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 2.400 130.520 ;
    END
  END left_top_grid_pin_46_
  PIN left_top_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 2.400 133.240 ;
    END
  END left_top_grid_pin_47_
  PIN left_top_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 2.400 135.960 ;
    END
  END left_top_grid_pin_48_
  PIN left_top_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 2.400 138.680 ;
    END
  END left_top_grid_pin_49_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 2.400 ;
    END
  END prog_clk
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 1.400 140.000 2.000 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_top_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 118.360 140.000 118.960 ;
    END
  END right_top_grid_pin_42_
  PIN right_top_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 121.080 140.000 121.680 ;
    END
  END right_top_grid_pin_43_
  PIN right_top_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 123.800 140.000 124.400 ;
    END
  END right_top_grid_pin_44_
  PIN right_top_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 126.520 140.000 127.120 ;
    END
  END right_top_grid_pin_45_
  PIN right_top_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 129.920 140.000 130.520 ;
    END
  END right_top_grid_pin_46_
  PIN right_top_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 132.640 140.000 133.240 ;
    END
  END right_top_grid_pin_47_
  PIN right_top_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 135.360 140.000 135.960 ;
    END
  END right_top_grid_pin_48_
  PIN right_top_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 138.080 140.000 138.680 ;
    END
  END right_top_grid_pin_49_
  PIN top_left_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 137.600 1.750 140.000 ;
    END
  END top_left_grid_pin_34_
  PIN top_left_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 137.600 4.510 140.000 ;
    END
  END top_left_grid_pin_35_
  PIN top_left_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 137.600 7.270 140.000 ;
    END
  END top_left_grid_pin_36_
  PIN top_left_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 137.600 10.490 140.000 ;
    END
  END top_left_grid_pin_37_
  PIN top_left_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 137.600 13.250 140.000 ;
    END
  END top_left_grid_pin_38_
  PIN top_left_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 137.600 16.010 140.000 ;
    END
  END top_left_grid_pin_39_
  PIN top_left_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 137.600 19.230 140.000 ;
    END
  END top_left_grid_pin_40_
  PIN top_left_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 137.600 21.990 140.000 ;
    END
  END top_left_grid_pin_41_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 1.450 10.640 134.320 130.180 ;
      LAYER met2 ;
        RECT 2.030 137.320 3.950 138.565 ;
        RECT 4.790 137.320 6.710 138.565 ;
        RECT 7.550 137.320 9.930 138.565 ;
        RECT 10.770 137.320 12.690 138.565 ;
        RECT 13.530 137.320 15.450 138.565 ;
        RECT 16.290 137.320 18.670 138.565 ;
        RECT 19.510 137.320 21.430 138.565 ;
        RECT 22.270 137.320 24.190 138.565 ;
        RECT 25.030 137.320 27.410 138.565 ;
        RECT 28.250 137.320 30.170 138.565 ;
        RECT 31.010 137.320 32.930 138.565 ;
        RECT 33.770 137.320 36.150 138.565 ;
        RECT 36.990 137.320 38.910 138.565 ;
        RECT 39.750 137.320 41.670 138.565 ;
        RECT 42.510 137.320 44.890 138.565 ;
        RECT 45.730 137.320 47.650 138.565 ;
        RECT 48.490 137.320 50.410 138.565 ;
        RECT 51.250 137.320 53.630 138.565 ;
        RECT 54.470 137.320 56.390 138.565 ;
        RECT 57.230 137.320 59.150 138.565 ;
        RECT 59.990 137.320 62.370 138.565 ;
        RECT 63.210 137.320 65.130 138.565 ;
        RECT 65.970 137.320 67.890 138.565 ;
        RECT 68.730 137.320 71.110 138.565 ;
        RECT 71.950 137.320 73.870 138.565 ;
        RECT 74.710 137.320 76.630 138.565 ;
        RECT 77.470 137.320 79.850 138.565 ;
        RECT 80.690 137.320 82.610 138.565 ;
        RECT 83.450 137.320 85.370 138.565 ;
        RECT 86.210 137.320 88.590 138.565 ;
        RECT 89.430 137.320 91.350 138.565 ;
        RECT 92.190 137.320 94.110 138.565 ;
        RECT 94.950 137.320 97.330 138.565 ;
        RECT 98.170 137.320 100.090 138.565 ;
        RECT 100.930 137.320 102.850 138.565 ;
        RECT 103.690 137.320 106.070 138.565 ;
        RECT 106.910 137.320 108.830 138.565 ;
        RECT 109.670 137.320 111.590 138.565 ;
        RECT 112.430 137.320 114.810 138.565 ;
        RECT 115.650 137.320 117.570 138.565 ;
        RECT 118.410 137.320 120.330 138.565 ;
        RECT 121.170 137.320 123.550 138.565 ;
        RECT 124.390 137.320 126.310 138.565 ;
        RECT 127.150 137.320 129.070 138.565 ;
        RECT 129.910 137.320 132.290 138.565 ;
        RECT 133.130 137.320 135.050 138.565 ;
        RECT 135.890 137.320 137.810 138.565 ;
        RECT 1.480 2.680 138.370 137.320 ;
        RECT 1.480 1.515 22.810 2.680 ;
        RECT 23.650 1.515 69.270 2.680 ;
        RECT 70.110 1.515 115.730 2.680 ;
        RECT 116.570 1.515 138.370 2.680 ;
      LAYER met3 ;
        RECT 2.800 137.680 137.200 138.545 ;
        RECT 2.400 136.360 138.395 137.680 ;
        RECT 2.800 134.960 137.200 136.360 ;
        RECT 2.400 133.640 138.395 134.960 ;
        RECT 2.800 132.240 137.200 133.640 ;
        RECT 2.400 130.920 138.395 132.240 ;
        RECT 2.800 129.520 137.200 130.920 ;
        RECT 2.400 127.520 138.395 129.520 ;
        RECT 2.800 126.120 137.200 127.520 ;
        RECT 2.400 124.800 138.395 126.120 ;
        RECT 2.800 123.400 137.200 124.800 ;
        RECT 2.400 122.080 138.395 123.400 ;
        RECT 2.800 120.680 137.200 122.080 ;
        RECT 2.400 119.360 138.395 120.680 ;
        RECT 2.800 117.960 137.200 119.360 ;
        RECT 2.400 116.640 138.395 117.960 ;
        RECT 2.800 115.240 137.200 116.640 ;
        RECT 2.400 113.240 138.395 115.240 ;
        RECT 2.800 111.840 137.200 113.240 ;
        RECT 2.400 110.520 138.395 111.840 ;
        RECT 2.800 109.120 137.200 110.520 ;
        RECT 2.400 107.800 138.395 109.120 ;
        RECT 2.800 106.400 137.200 107.800 ;
        RECT 2.400 105.080 138.395 106.400 ;
        RECT 2.800 103.680 137.200 105.080 ;
        RECT 2.400 102.360 138.395 103.680 ;
        RECT 2.800 100.960 137.200 102.360 ;
        RECT 2.400 98.960 138.395 100.960 ;
        RECT 2.800 97.560 137.200 98.960 ;
        RECT 2.400 96.240 138.395 97.560 ;
        RECT 2.800 94.840 137.200 96.240 ;
        RECT 2.400 93.520 138.395 94.840 ;
        RECT 2.800 92.120 137.200 93.520 ;
        RECT 2.400 90.800 138.395 92.120 ;
        RECT 2.800 89.400 137.200 90.800 ;
        RECT 2.400 88.080 138.395 89.400 ;
        RECT 2.800 86.680 137.200 88.080 ;
        RECT 2.400 84.680 138.395 86.680 ;
        RECT 2.800 83.280 137.200 84.680 ;
        RECT 2.400 81.960 138.395 83.280 ;
        RECT 2.800 80.560 137.200 81.960 ;
        RECT 2.400 79.240 138.395 80.560 ;
        RECT 2.800 77.840 137.200 79.240 ;
        RECT 2.400 76.520 138.395 77.840 ;
        RECT 2.800 75.120 137.200 76.520 ;
        RECT 2.400 73.800 138.395 75.120 ;
        RECT 2.800 72.400 137.200 73.800 ;
        RECT 2.400 70.400 138.395 72.400 ;
        RECT 2.800 69.000 137.200 70.400 ;
        RECT 2.400 67.680 138.395 69.000 ;
        RECT 2.800 66.280 137.200 67.680 ;
        RECT 2.400 64.960 138.395 66.280 ;
        RECT 2.800 63.560 137.200 64.960 ;
        RECT 2.400 62.240 138.395 63.560 ;
        RECT 2.800 60.840 137.200 62.240 ;
        RECT 2.400 59.520 138.395 60.840 ;
        RECT 2.800 58.120 137.200 59.520 ;
        RECT 2.400 56.120 138.395 58.120 ;
        RECT 2.800 54.720 137.200 56.120 ;
        RECT 2.400 53.400 138.395 54.720 ;
        RECT 2.800 52.000 137.200 53.400 ;
        RECT 2.400 50.680 138.395 52.000 ;
        RECT 2.800 49.280 137.200 50.680 ;
        RECT 2.400 47.960 138.395 49.280 ;
        RECT 2.800 46.560 137.200 47.960 ;
        RECT 2.400 45.240 138.395 46.560 ;
        RECT 2.800 43.840 137.200 45.240 ;
        RECT 2.400 41.840 138.395 43.840 ;
        RECT 2.800 40.440 137.200 41.840 ;
        RECT 2.400 39.120 138.395 40.440 ;
        RECT 2.800 37.720 137.200 39.120 ;
        RECT 2.400 36.400 138.395 37.720 ;
        RECT 2.800 35.000 137.200 36.400 ;
        RECT 2.400 33.680 138.395 35.000 ;
        RECT 2.800 32.280 137.200 33.680 ;
        RECT 2.400 30.960 138.395 32.280 ;
        RECT 2.800 29.560 137.200 30.960 ;
        RECT 2.400 27.560 138.395 29.560 ;
        RECT 2.800 26.160 137.200 27.560 ;
        RECT 2.400 24.840 138.395 26.160 ;
        RECT 2.800 23.440 137.200 24.840 ;
        RECT 2.400 22.120 138.395 23.440 ;
        RECT 2.800 20.720 137.200 22.120 ;
        RECT 2.400 19.400 138.395 20.720 ;
        RECT 2.800 18.000 137.200 19.400 ;
        RECT 2.400 16.680 138.395 18.000 ;
        RECT 2.800 15.280 137.200 16.680 ;
        RECT 2.400 13.280 138.395 15.280 ;
        RECT 2.800 11.880 137.200 13.280 ;
        RECT 2.400 10.560 138.395 11.880 ;
        RECT 2.800 9.160 137.200 10.560 ;
        RECT 2.400 7.840 138.395 9.160 ;
        RECT 2.800 6.440 137.200 7.840 ;
        RECT 2.400 5.120 138.395 6.440 ;
        RECT 2.800 3.720 137.200 5.120 ;
        RECT 2.400 2.400 138.395 3.720 ;
        RECT 2.800 1.535 137.200 2.400 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 123.905 128.080 ;
  END
END sb_1__0_
END LIBRARY

