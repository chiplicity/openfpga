magic
tech sky130A
magscale 1 2
timestamp 1606227617
<< locali >>
rect 4629 12631 4663 12801
rect 8861 12087 8895 12257
rect 11529 12087 11563 12189
rect 10333 10455 10367 10557
rect 17049 10455 17083 10557
rect 18429 10455 18463 10557
rect 6837 9367 6871 9537
rect 11345 9503 11379 9605
rect 4905 8891 4939 9061
rect 4445 8279 4479 8585
rect 5549 8279 5583 8449
rect 18981 8279 19015 8517
rect 5491 8245 5583 8279
rect 18521 7871 18555 8041
rect 15669 7191 15703 7497
rect 17601 5559 17635 5729
rect 11069 5151 11103 5253
rect 16037 4675 16071 4777
rect 15117 3587 15151 3689
rect 12541 3383 12575 3485
rect 15945 2975 15979 3145
rect 11161 2295 11195 2397
rect 13277 2295 13311 2465
<< viali >>
rect 1961 19465 1995 19499
rect 18705 19465 18739 19499
rect 20729 19465 20763 19499
rect 1777 19261 1811 19295
rect 2329 19261 2363 19295
rect 18521 19261 18555 19295
rect 20545 19261 20579 19295
rect 2513 19125 2547 19159
rect 1961 18921 1995 18955
rect 17877 18853 17911 18887
rect 1777 18785 1811 18819
rect 17601 18785 17635 18819
rect 1961 18377 1995 18411
rect 20729 18377 20763 18411
rect 1777 18173 1811 18207
rect 20545 18173 20579 18207
rect 2421 17765 2455 17799
rect 19901 17765 19935 17799
rect 1593 17697 1627 17731
rect 2145 17697 2179 17731
rect 19625 17697 19659 17731
rect 1777 17561 1811 17595
rect 1961 17289 1995 17323
rect 20177 17289 20211 17323
rect 20729 17289 20763 17323
rect 1777 17085 1811 17119
rect 19993 17085 20027 17119
rect 20545 17085 20579 17119
rect 1961 16745 1995 16779
rect 20453 16745 20487 16779
rect 1777 16609 1811 16643
rect 20269 16609 20303 16643
rect 1961 16201 1995 16235
rect 3709 16201 3743 16235
rect 14565 16201 14599 16235
rect 20729 16201 20763 16235
rect 1777 15997 1811 16031
rect 3525 15997 3559 16031
rect 14381 15997 14415 16031
rect 20545 15997 20579 16031
rect 1961 15657 1995 15691
rect 2513 15657 2547 15691
rect 19901 15657 19935 15691
rect 20453 15657 20487 15691
rect 4353 15589 4387 15623
rect 13737 15589 13771 15623
rect 1777 15521 1811 15555
rect 2329 15521 2363 15555
rect 4077 15521 4111 15555
rect 13461 15521 13495 15555
rect 19717 15521 19751 15555
rect 20269 15521 20303 15555
rect 2513 15113 2547 15147
rect 3065 15113 3099 15147
rect 3617 15113 3651 15147
rect 6193 15113 6227 15147
rect 20729 15113 20763 15147
rect 1961 15045 1995 15079
rect 11805 15045 11839 15079
rect 14289 14977 14323 15011
rect 1777 14909 1811 14943
rect 2329 14909 2363 14943
rect 2881 14909 2915 14943
rect 3433 14909 3467 14943
rect 6009 14909 6043 14943
rect 11621 14909 11655 14943
rect 14105 14909 14139 14943
rect 19441 14909 19475 14943
rect 19993 14909 20027 14943
rect 20545 14909 20579 14943
rect 13645 14773 13679 14807
rect 14013 14773 14047 14807
rect 16957 14773 16991 14807
rect 19625 14773 19659 14807
rect 20177 14773 20211 14807
rect 9137 14569 9171 14603
rect 17509 14569 17543 14603
rect 19901 14569 19935 14603
rect 20453 14569 20487 14603
rect 2145 14501 2179 14535
rect 2973 14501 3007 14535
rect 6653 14501 6687 14535
rect 8002 14501 8036 14535
rect 11590 14501 11624 14535
rect 18030 14501 18064 14535
rect 1869 14433 1903 14467
rect 6377 14433 6411 14467
rect 10701 14433 10735 14467
rect 11345 14433 11379 14467
rect 13001 14433 13035 14467
rect 13268 14433 13302 14467
rect 16396 14433 16430 14467
rect 19717 14433 19751 14467
rect 20269 14433 20303 14467
rect 3065 14365 3099 14399
rect 3157 14365 3191 14399
rect 7757 14365 7791 14399
rect 10793 14365 10827 14399
rect 10885 14365 10919 14399
rect 16129 14365 16163 14399
rect 17785 14365 17819 14399
rect 12725 14297 12759 14331
rect 2605 14229 2639 14263
rect 10333 14229 10367 14263
rect 14381 14229 14415 14263
rect 19165 14229 19199 14263
rect 2605 14025 2639 14059
rect 7021 14025 7055 14059
rect 16681 14025 16715 14059
rect 10333 13957 10367 13991
rect 16957 13957 16991 13991
rect 1869 13889 1903 13923
rect 5181 13889 5215 13923
rect 7665 13889 7699 13923
rect 10977 13889 11011 13923
rect 11621 13889 11655 13923
rect 14473 13889 14507 13923
rect 17601 13889 17635 13923
rect 19717 13889 19751 13923
rect 20453 13889 20487 13923
rect 1685 13821 1719 13855
rect 2421 13821 2455 13855
rect 2973 13821 3007 13855
rect 10701 13821 10735 13855
rect 10793 13821 10827 13855
rect 11345 13821 11379 13855
rect 12817 13821 12851 13855
rect 13084 13821 13118 13855
rect 15301 13821 15335 13855
rect 15568 13821 15602 13855
rect 18061 13821 18095 13855
rect 18337 13821 18371 13855
rect 18981 13821 19015 13855
rect 19533 13821 19567 13855
rect 20269 13821 20303 13855
rect 3240 13753 3274 13787
rect 4997 13753 5031 13787
rect 8033 13753 8067 13787
rect 4353 13685 4387 13719
rect 4629 13685 4663 13719
rect 5089 13685 5123 13719
rect 7389 13685 7423 13719
rect 7481 13685 7515 13719
rect 14197 13685 14231 13719
rect 17325 13685 17359 13719
rect 17417 13685 17451 13719
rect 19165 13685 19199 13719
rect 1593 13481 1627 13515
rect 2973 13481 3007 13515
rect 3433 13481 3467 13515
rect 6653 13481 6687 13515
rect 7021 13481 7055 13515
rect 7665 13481 7699 13515
rect 11161 13481 11195 13515
rect 11437 13481 11471 13515
rect 12909 13481 12943 13515
rect 15577 13481 15611 13515
rect 16589 13481 16623 13515
rect 16957 13481 16991 13515
rect 17049 13481 17083 13515
rect 20269 13481 20303 13515
rect 2329 13413 2363 13447
rect 4414 13413 4448 13447
rect 8125 13413 8159 13447
rect 13001 13413 13035 13447
rect 13820 13413 13854 13447
rect 18144 13413 18178 13447
rect 1409 13345 1443 13379
rect 3341 13345 3375 13379
rect 8033 13345 8067 13379
rect 10048 13345 10082 13379
rect 11805 13345 11839 13379
rect 11897 13345 11931 13379
rect 13553 13345 13587 13379
rect 15945 13345 15979 13379
rect 16037 13345 16071 13379
rect 20177 13345 20211 13379
rect 2421 13277 2455 13311
rect 2605 13277 2639 13311
rect 3617 13277 3651 13311
rect 4169 13277 4203 13311
rect 7113 13277 7147 13311
rect 7297 13277 7331 13311
rect 8217 13277 8251 13311
rect 9781 13277 9815 13311
rect 11989 13277 12023 13311
rect 13185 13277 13219 13311
rect 16221 13277 16255 13311
rect 17141 13277 17175 13311
rect 17877 13277 17911 13311
rect 20361 13277 20395 13311
rect 1961 13141 1995 13175
rect 5549 13141 5583 13175
rect 12541 13141 12575 13175
rect 14933 13141 14967 13175
rect 19257 13141 19291 13175
rect 19809 13141 19843 13175
rect 1777 12937 1811 12971
rect 4169 12937 4203 12971
rect 4721 12937 4755 12971
rect 5733 12937 5767 12971
rect 8217 12937 8251 12971
rect 10057 12937 10091 12971
rect 13921 12937 13955 12971
rect 20269 12937 20303 12971
rect 12909 12869 12943 12903
rect 16957 12869 16991 12903
rect 2237 12801 2271 12835
rect 2421 12801 2455 12835
rect 4629 12801 4663 12835
rect 5365 12801 5399 12835
rect 6377 12801 6411 12835
rect 8677 12801 8711 12835
rect 10701 12801 10735 12835
rect 13461 12801 13495 12835
rect 14381 12801 14415 12835
rect 14565 12801 14599 12835
rect 17509 12801 17543 12835
rect 20729 12801 20763 12835
rect 2145 12733 2179 12767
rect 2789 12733 2823 12767
rect 3056 12665 3090 12699
rect 5089 12733 5123 12767
rect 6101 12733 6135 12767
rect 6837 12733 6871 12767
rect 10968 12733 11002 12767
rect 13277 12733 13311 12767
rect 14289 12733 14323 12767
rect 15301 12733 15335 12767
rect 15557 12733 15591 12767
rect 18061 12733 18095 12767
rect 18889 12733 18923 12767
rect 19156 12733 19190 12767
rect 20545 12733 20579 12767
rect 7104 12665 7138 12699
rect 8944 12665 8978 12699
rect 18337 12665 18371 12699
rect 4629 12597 4663 12631
rect 5181 12597 5215 12631
rect 6193 12597 6227 12631
rect 12081 12597 12115 12631
rect 13369 12597 13403 12631
rect 16681 12597 16715 12631
rect 17325 12597 17359 12631
rect 17417 12597 17451 12631
rect 1685 12393 1719 12427
rect 2421 12393 2455 12427
rect 4077 12393 4111 12427
rect 4445 12393 4479 12427
rect 6469 12393 6503 12427
rect 6745 12393 6779 12427
rect 7941 12393 7975 12427
rect 10057 12393 10091 12427
rect 10701 12393 10735 12427
rect 14197 12393 14231 12427
rect 14565 12393 14599 12427
rect 17877 12393 17911 12427
rect 2513 12325 2547 12359
rect 3341 12325 3375 12359
rect 7205 12325 7239 12359
rect 8309 12325 8343 12359
rect 17325 12325 17359 12359
rect 1501 12257 1535 12291
rect 3065 12257 3099 12291
rect 5345 12257 5379 12291
rect 7113 12257 7147 12291
rect 8401 12257 8435 12291
rect 8861 12257 8895 12291
rect 9137 12257 9171 12291
rect 10149 12257 10183 12291
rect 11069 12257 11103 12291
rect 12449 12257 12483 12291
rect 12909 12257 12943 12291
rect 13553 12257 13587 12291
rect 15669 12257 15703 12291
rect 17233 12257 17267 12291
rect 18245 12257 18279 12291
rect 19993 12257 20027 12291
rect 2697 12189 2731 12223
rect 4537 12189 4571 12223
rect 4721 12189 4755 12223
rect 5089 12189 5123 12223
rect 7297 12189 7331 12223
rect 8585 12189 8619 12223
rect 10241 12189 10275 12223
rect 11161 12189 11195 12223
rect 11345 12189 11379 12223
rect 11529 12189 11563 12223
rect 11713 12189 11747 12223
rect 13001 12189 13035 12223
rect 13185 12189 13219 12223
rect 14657 12189 14691 12223
rect 14841 12189 14875 12223
rect 15761 12189 15795 12223
rect 15945 12189 15979 12223
rect 17509 12189 17543 12223
rect 18337 12189 18371 12223
rect 18521 12189 18555 12223
rect 18889 12189 18923 12223
rect 20085 12189 20119 12223
rect 20269 12189 20303 12223
rect 9689 12121 9723 12155
rect 16865 12121 16899 12155
rect 2053 12053 2087 12087
rect 8861 12053 8895 12087
rect 8953 12053 8987 12087
rect 11529 12053 11563 12087
rect 12265 12053 12299 12087
rect 12541 12053 12575 12087
rect 15301 12053 15335 12087
rect 19441 12053 19475 12087
rect 19625 12053 19659 12087
rect 1593 11849 1627 11883
rect 4721 11849 4755 11883
rect 8493 11849 8527 11883
rect 8769 11849 8803 11883
rect 10701 11849 10735 11883
rect 12449 11849 12483 11883
rect 13461 11849 13495 11883
rect 15301 11849 15335 11883
rect 17693 11849 17727 11883
rect 18061 11849 18095 11883
rect 21005 11849 21039 11883
rect 1961 11781 1995 11815
rect 2605 11713 2639 11747
rect 5733 11713 5767 11747
rect 7113 11713 7147 11747
rect 9321 11713 9355 11747
rect 11253 11713 11287 11747
rect 12909 11713 12943 11747
rect 13001 11713 13035 11747
rect 14105 11713 14139 11747
rect 15761 11713 15795 11747
rect 15945 11713 15979 11747
rect 18613 11713 18647 11747
rect 1409 11645 1443 11679
rect 3341 11645 3375 11679
rect 9229 11645 9263 11679
rect 11069 11645 11103 11679
rect 16313 11645 16347 11679
rect 18429 11645 18463 11679
rect 19625 11645 19659 11679
rect 19892 11645 19926 11679
rect 2329 11577 2363 11611
rect 3586 11577 3620 11611
rect 5549 11577 5583 11611
rect 5641 11577 5675 11611
rect 7358 11577 7392 11611
rect 9137 11577 9171 11611
rect 11897 11577 11931 11611
rect 12817 11577 12851 11611
rect 13921 11577 13955 11611
rect 16580 11577 16614 11611
rect 18521 11577 18555 11611
rect 2421 11509 2455 11543
rect 5181 11509 5215 11543
rect 11161 11509 11195 11543
rect 13829 11509 13863 11543
rect 15669 11509 15703 11543
rect 2053 11305 2087 11339
rect 5273 11305 5307 11339
rect 6469 11305 6503 11339
rect 7849 11305 7883 11339
rect 8585 11305 8619 11339
rect 10057 11305 10091 11339
rect 12541 11305 12575 11339
rect 13185 11305 13219 11339
rect 13829 11305 13863 11339
rect 14841 11305 14875 11339
rect 15853 11305 15887 11339
rect 18521 11305 18555 11339
rect 19533 11305 19567 11339
rect 20453 11305 20487 11339
rect 20913 11305 20947 11339
rect 3341 11237 3375 11271
rect 9045 11237 9079 11271
rect 11406 11237 11440 11271
rect 14197 11237 14231 11271
rect 2421 11169 2455 11203
rect 2513 11169 2547 11203
rect 3065 11169 3099 11203
rect 5181 11169 5215 11203
rect 6837 11169 6871 11203
rect 7941 11169 7975 11203
rect 8953 11169 8987 11203
rect 15025 11169 15059 11203
rect 15761 11169 15795 11203
rect 16221 11169 16255 11203
rect 17408 11169 17442 11203
rect 20269 11169 20303 11203
rect 2697 11101 2731 11135
rect 5457 11101 5491 11135
rect 6929 11101 6963 11135
rect 7113 11101 7147 11135
rect 8033 11101 8067 11135
rect 9229 11101 9263 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 11161 11101 11195 11135
rect 13277 11101 13311 11135
rect 13461 11101 13495 11135
rect 14289 11101 14323 11135
rect 14381 11101 14415 11135
rect 16313 11101 16347 11135
rect 16497 11101 16531 11135
rect 17141 11101 17175 11135
rect 19625 11101 19659 11135
rect 19809 11101 19843 11135
rect 4813 11033 4847 11067
rect 7481 11033 7515 11067
rect 9689 11033 9723 11067
rect 12817 11033 12851 11067
rect 15577 11033 15611 11067
rect 19165 11033 19199 11067
rect 3249 10761 3283 10795
rect 8217 10761 8251 10795
rect 10241 10761 10275 10795
rect 14105 10761 14139 10795
rect 15117 10761 15151 10795
rect 5825 10693 5859 10727
rect 3525 10625 3559 10659
rect 6837 10625 6871 10659
rect 8861 10625 8895 10659
rect 14657 10625 14691 10659
rect 15577 10625 15611 10659
rect 15761 10625 15795 10659
rect 16681 10625 16715 10659
rect 20637 10625 20671 10659
rect 20729 10625 20763 10659
rect 1869 10557 1903 10591
rect 4169 10557 4203 10591
rect 4436 10557 4470 10591
rect 6009 10557 6043 10591
rect 10333 10557 10367 10591
rect 10517 10557 10551 10591
rect 10773 10557 10807 10591
rect 12449 10557 12483 10591
rect 12716 10557 12750 10591
rect 17049 10557 17083 10591
rect 2136 10489 2170 10523
rect 7104 10489 7138 10523
rect 9128 10489 9162 10523
rect 14473 10489 14507 10523
rect 15485 10489 15519 10523
rect 16497 10489 16531 10523
rect 18429 10557 18463 10591
rect 18521 10557 18555 10591
rect 18788 10557 18822 10591
rect 17141 10489 17175 10523
rect 5549 10421 5583 10455
rect 10333 10421 10367 10455
rect 11897 10421 11931 10455
rect 13829 10421 13863 10455
rect 14565 10421 14599 10455
rect 16129 10421 16163 10455
rect 16589 10421 16623 10455
rect 17049 10421 17083 10455
rect 18429 10421 18463 10455
rect 19901 10421 19935 10455
rect 20177 10421 20211 10455
rect 20545 10421 20579 10455
rect 3065 10217 3099 10251
rect 7389 10217 7423 10251
rect 7665 10217 7699 10251
rect 9689 10217 9723 10251
rect 10609 10217 10643 10251
rect 12081 10217 12115 10251
rect 16865 10217 16899 10251
rect 4620 10149 4654 10183
rect 11069 10149 11103 10183
rect 12900 10149 12934 10183
rect 17386 10149 17420 10183
rect 19432 10149 19466 10183
rect 1952 10081 1986 10115
rect 4353 10081 4387 10115
rect 6265 10081 6299 10115
rect 7849 10081 7883 10115
rect 8208 10081 8242 10115
rect 10977 10081 11011 10115
rect 11989 10081 12023 10115
rect 12633 10081 12667 10115
rect 14289 10081 14323 10115
rect 15741 10081 15775 10115
rect 17141 10081 17175 10115
rect 1685 10013 1719 10047
rect 6009 10013 6043 10047
rect 7941 10013 7975 10047
rect 11253 10013 11287 10047
rect 12265 10013 12299 10047
rect 14565 10013 14599 10047
rect 15485 10013 15519 10047
rect 19165 10013 19199 10047
rect 11621 9945 11655 9979
rect 5733 9877 5767 9911
rect 9321 9877 9355 9911
rect 14013 9877 14047 9911
rect 18521 9877 18555 9911
rect 20545 9877 20579 9911
rect 15393 9673 15427 9707
rect 1869 9605 1903 9639
rect 2881 9605 2915 9639
rect 4445 9605 4479 9639
rect 6929 9605 6963 9639
rect 10149 9605 10183 9639
rect 11345 9605 11379 9639
rect 12817 9605 12851 9639
rect 15669 9605 15703 9639
rect 18521 9605 18555 9639
rect 2513 9537 2547 9571
rect 3433 9537 3467 9571
rect 4905 9537 4939 9571
rect 5089 9537 5123 9571
rect 6009 9537 6043 9571
rect 6837 9537 6871 9571
rect 7389 9537 7423 9571
rect 7481 9537 7515 9571
rect 8769 9537 8803 9571
rect 10977 9537 11011 9571
rect 5917 9469 5951 9503
rect 3249 9401 3283 9435
rect 4813 9401 4847 9435
rect 13461 9537 13495 9571
rect 14013 9537 14047 9571
rect 16221 9537 16255 9571
rect 17233 9537 17267 9571
rect 19119 9537 19153 9571
rect 10793 9469 10827 9503
rect 11345 9469 11379 9503
rect 11437 9469 11471 9503
rect 16037 9469 16071 9503
rect 18981 9469 19015 9503
rect 19533 9469 19567 9503
rect 19800 9469 19834 9503
rect 9036 9401 9070 9435
rect 11713 9401 11747 9435
rect 13185 9401 13219 9435
rect 14258 9401 14292 9435
rect 18889 9401 18923 9435
rect 1409 9333 1443 9367
rect 2237 9333 2271 9367
rect 2329 9333 2363 9367
rect 3341 9333 3375 9367
rect 5457 9333 5491 9367
rect 5825 9333 5859 9367
rect 6837 9333 6871 9367
rect 7297 9333 7331 9367
rect 10425 9333 10459 9367
rect 10885 9333 10919 9367
rect 13277 9333 13311 9367
rect 16129 9333 16163 9367
rect 16681 9333 16715 9367
rect 17049 9333 17083 9367
rect 17141 9333 17175 9367
rect 20913 9333 20947 9367
rect 1961 9129 1995 9163
rect 2973 9129 3007 9163
rect 3341 9129 3375 9163
rect 3433 9129 3467 9163
rect 4077 9129 4111 9163
rect 5089 9129 5123 9163
rect 5457 9129 5491 9163
rect 8125 9129 8159 9163
rect 14105 9129 14139 9163
rect 15301 9129 15335 9163
rect 15669 9129 15703 9163
rect 16681 9129 16715 9163
rect 18797 9129 18831 9163
rect 20269 9129 20303 9163
rect 2329 9061 2363 9095
rect 4905 9061 4939 9095
rect 4445 8993 4479 9027
rect 2421 8925 2455 8959
rect 2513 8925 2547 8959
rect 3525 8925 3559 8959
rect 4537 8925 4571 8959
rect 4721 8925 4755 8959
rect 6469 8993 6503 9027
rect 6736 8993 6770 9027
rect 8493 8993 8527 9027
rect 8585 8993 8619 9027
rect 10609 8993 10643 9027
rect 12716 8993 12750 9027
rect 14289 8993 14323 9027
rect 17684 8993 17718 9027
rect 19073 8993 19107 9027
rect 20177 8993 20211 9027
rect 20913 8993 20947 9027
rect 5549 8925 5583 8959
rect 5641 8925 5675 8959
rect 8677 8925 8711 8959
rect 12449 8925 12483 8959
rect 15761 8925 15795 8959
rect 15853 8925 15887 8959
rect 16773 8925 16807 8959
rect 16865 8925 16899 8959
rect 17417 8925 17451 8959
rect 19349 8925 19383 8959
rect 20453 8925 20487 8959
rect 4905 8857 4939 8891
rect 7849 8857 7883 8891
rect 16313 8857 16347 8891
rect 11897 8789 11931 8823
rect 13829 8789 13863 8823
rect 19809 8789 19843 8823
rect 3157 8585 3191 8619
rect 3617 8585 3651 8619
rect 4445 8585 4479 8619
rect 4629 8585 4663 8619
rect 6837 8585 6871 8619
rect 7849 8585 7883 8619
rect 9965 8585 9999 8619
rect 11345 8585 11379 8619
rect 13829 8585 13863 8619
rect 15485 8585 15519 8619
rect 19349 8585 19383 8619
rect 1777 8449 1811 8483
rect 4169 8449 4203 8483
rect 2044 8313 2078 8347
rect 8861 8517 8895 8551
rect 9137 8517 9171 8551
rect 16405 8517 16439 8551
rect 17601 8517 17635 8551
rect 18981 8517 19015 8551
rect 5089 8449 5123 8483
rect 5273 8449 5307 8483
rect 5549 8449 5583 8483
rect 6193 8449 6227 8483
rect 7481 8449 7515 8483
rect 8493 8449 8527 8483
rect 9689 8449 9723 8483
rect 10425 8449 10459 8483
rect 10609 8449 10643 8483
rect 11805 8449 11839 8483
rect 11989 8449 12023 8483
rect 16865 8449 16899 8483
rect 17049 8449 17083 8483
rect 18705 8449 18739 8483
rect 6009 8381 6043 8415
rect 7297 8381 7331 8415
rect 9045 8381 9079 8415
rect 12449 8381 12483 8415
rect 14105 8381 14139 8415
rect 14361 8381 14395 8415
rect 17417 8381 17451 8415
rect 18613 8381 18647 8415
rect 7205 8313 7239 8347
rect 8217 8313 8251 8347
rect 9505 8313 9539 8347
rect 10793 8313 10827 8347
rect 12716 8313 12750 8347
rect 16773 8313 16807 8347
rect 19165 8381 19199 8415
rect 19717 8381 19751 8415
rect 19984 8381 20018 8415
rect 3985 8245 4019 8279
rect 4077 8245 4111 8279
rect 4445 8245 4479 8279
rect 4997 8245 5031 8279
rect 5457 8245 5491 8279
rect 5641 8245 5675 8279
rect 6101 8245 6135 8279
rect 8309 8245 8343 8279
rect 9597 8245 9631 8279
rect 10333 8245 10367 8279
rect 11713 8245 11747 8279
rect 15761 8245 15795 8279
rect 18153 8245 18187 8279
rect 18521 8245 18555 8279
rect 18981 8245 19015 8279
rect 21097 8245 21131 8279
rect 3525 8041 3559 8075
rect 5089 8041 5123 8075
rect 6561 8041 6595 8075
rect 9321 8041 9355 8075
rect 10057 8041 10091 8075
rect 10149 8041 10183 8075
rect 10701 8041 10735 8075
rect 11069 8041 11103 8075
rect 12541 8041 12575 8075
rect 12633 8041 12667 8075
rect 13185 8041 13219 8075
rect 13645 8041 13679 8075
rect 14197 8041 14231 8075
rect 16681 8041 16715 8075
rect 18521 8041 18555 8075
rect 20453 8041 20487 8075
rect 4445 7973 4479 8007
rect 5457 7973 5491 8007
rect 8208 7973 8242 8007
rect 11161 7973 11195 8007
rect 15568 7973 15602 8007
rect 17224 7973 17258 8007
rect 2421 7905 2455 7939
rect 2513 7905 2547 7939
rect 4537 7905 4571 7939
rect 6101 7905 6135 7939
rect 6929 7905 6963 7939
rect 7941 7905 7975 7939
rect 13553 7905 13587 7939
rect 14565 7905 14599 7939
rect 15301 7905 15335 7939
rect 16957 7905 16991 7939
rect 18869 7905 18903 7939
rect 20269 7905 20303 7939
rect 2697 7837 2731 7871
rect 4721 7837 4755 7871
rect 5549 7837 5583 7871
rect 5641 7837 5675 7871
rect 7021 7837 7055 7871
rect 7205 7837 7239 7871
rect 10241 7837 10275 7871
rect 11253 7837 11287 7871
rect 12817 7837 12851 7871
rect 13737 7837 13771 7871
rect 14657 7837 14691 7871
rect 14841 7837 14875 7871
rect 18521 7837 18555 7871
rect 18613 7837 18647 7871
rect 20913 7837 20947 7871
rect 4077 7769 4111 7803
rect 9689 7769 9723 7803
rect 12173 7769 12207 7803
rect 2053 7701 2087 7735
rect 18337 7701 18371 7735
rect 19993 7701 20027 7735
rect 2237 7497 2271 7531
rect 4445 7497 4479 7531
rect 5549 7497 5583 7531
rect 6837 7497 6871 7531
rect 7849 7497 7883 7531
rect 10701 7497 10735 7531
rect 13461 7497 13495 7531
rect 15669 7497 15703 7531
rect 18153 7497 18187 7531
rect 19165 7497 19199 7531
rect 10425 7429 10459 7463
rect 2881 7361 2915 7395
rect 3801 7361 3835 7395
rect 5089 7361 5123 7395
rect 6101 7361 6135 7395
rect 7389 7361 7423 7395
rect 8401 7361 8435 7395
rect 9045 7361 9079 7395
rect 11253 7361 11287 7395
rect 13093 7361 13127 7395
rect 13921 7361 13955 7395
rect 14105 7361 14139 7395
rect 15485 7361 15519 7395
rect 2605 7293 2639 7327
rect 4905 7293 4939 7327
rect 5917 7293 5951 7327
rect 8217 7293 8251 7327
rect 9312 7293 9346 7327
rect 13829 7293 13863 7327
rect 14657 7293 14691 7327
rect 15209 7293 15243 7327
rect 4813 7225 4847 7259
rect 7205 7225 7239 7259
rect 7297 7225 7331 7259
rect 16405 7361 16439 7395
rect 17325 7361 17359 7395
rect 17509 7361 17543 7395
rect 18705 7361 18739 7395
rect 19717 7361 19751 7395
rect 20729 7361 20763 7395
rect 16221 7293 16255 7327
rect 16313 7225 16347 7259
rect 18613 7225 18647 7259
rect 20545 7225 20579 7259
rect 20637 7225 20671 7259
rect 2697 7157 2731 7191
rect 3249 7157 3283 7191
rect 3617 7157 3651 7191
rect 3709 7157 3743 7191
rect 6009 7157 6043 7191
rect 8309 7157 8343 7191
rect 11069 7157 11103 7191
rect 11161 7157 11195 7191
rect 12449 7157 12483 7191
rect 12817 7157 12851 7191
rect 12909 7157 12943 7191
rect 14473 7157 14507 7191
rect 14841 7157 14875 7191
rect 15301 7157 15335 7191
rect 15669 7157 15703 7191
rect 15853 7157 15887 7191
rect 16865 7157 16899 7191
rect 17233 7157 17267 7191
rect 18521 7157 18555 7191
rect 19533 7157 19567 7191
rect 19625 7157 19659 7191
rect 20177 7157 20211 7191
rect 2053 6953 2087 6987
rect 4077 6953 4111 6987
rect 4537 6953 4571 6987
rect 5641 6953 5675 6987
rect 9689 6953 9723 6987
rect 13185 6953 13219 6987
rect 15301 6953 15335 6987
rect 15669 6953 15703 6987
rect 17325 6953 17359 6987
rect 18153 6953 18187 6987
rect 18797 6953 18831 6987
rect 19809 6953 19843 6987
rect 2421 6885 2455 6919
rect 3065 6885 3099 6919
rect 7113 6885 7147 6919
rect 8125 6885 8159 6919
rect 14289 6885 14323 6919
rect 16681 6885 16715 6919
rect 16773 6885 16807 6919
rect 19165 6885 19199 6919
rect 4445 6817 4479 6851
rect 5733 6817 5767 6851
rect 6653 6817 6687 6851
rect 7205 6817 7239 6851
rect 8217 6817 8251 6851
rect 10057 6817 10091 6851
rect 11796 6817 11830 6851
rect 17509 6817 17543 6851
rect 19257 6817 19291 6851
rect 20177 6817 20211 6851
rect 2513 6749 2547 6783
rect 2605 6749 2639 6783
rect 4629 6749 4663 6783
rect 5917 6749 5951 6783
rect 7389 6749 7423 6783
rect 8401 6749 8435 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 11529 6749 11563 6783
rect 14381 6749 14415 6783
rect 14565 6749 14599 6783
rect 15761 6749 15795 6783
rect 15945 6749 15979 6783
rect 16865 6749 16899 6783
rect 18245 6749 18279 6783
rect 18337 6749 18371 6783
rect 19349 6749 19383 6783
rect 20269 6749 20303 6783
rect 20361 6749 20395 6783
rect 6745 6681 6779 6715
rect 5273 6613 5307 6647
rect 6469 6613 6503 6647
rect 7757 6613 7791 6647
rect 12909 6613 12943 6647
rect 13921 6613 13955 6647
rect 16313 6613 16347 6647
rect 17785 6613 17819 6647
rect 3157 6409 3191 6443
rect 3433 6409 3467 6443
rect 9965 6409 9999 6443
rect 10977 6409 11011 6443
rect 13921 6409 13955 6443
rect 16957 6409 16991 6443
rect 19257 6409 19291 6443
rect 20269 6409 20303 6443
rect 12081 6341 12115 6375
rect 16589 6341 16623 6375
rect 3985 6273 4019 6307
rect 7389 6273 7423 6307
rect 8309 6273 8343 6307
rect 8401 6273 8435 6307
rect 9413 6273 9447 6307
rect 10609 6273 10643 6307
rect 11529 6273 11563 6307
rect 12541 6273 12575 6307
rect 14657 6273 14691 6307
rect 14749 6273 14783 6307
rect 15761 6273 15795 6307
rect 17509 6273 17543 6307
rect 18797 6273 18831 6307
rect 19717 6273 19751 6307
rect 19809 6273 19843 6307
rect 20821 6273 20855 6307
rect 1777 6205 1811 6239
rect 2044 6205 2078 6239
rect 4721 6205 4755 6239
rect 4813 6205 4847 6239
rect 5080 6205 5114 6239
rect 7297 6205 7331 6239
rect 8217 6205 8251 6239
rect 9321 6205 9355 6239
rect 10425 6205 10459 6239
rect 12265 6205 12299 6239
rect 12808 6205 12842 6239
rect 15669 6205 15703 6239
rect 16405 6205 16439 6239
rect 18613 6205 18647 6239
rect 3893 6137 3927 6171
rect 7205 6137 7239 6171
rect 10333 6137 10367 6171
rect 14565 6137 14599 6171
rect 17417 6137 17451 6171
rect 19625 6137 19659 6171
rect 20637 6137 20671 6171
rect 3801 6069 3835 6103
rect 4537 6069 4571 6103
rect 6193 6069 6227 6103
rect 6837 6069 6871 6103
rect 7849 6069 7883 6103
rect 8861 6069 8895 6103
rect 9229 6069 9263 6103
rect 11345 6069 11379 6103
rect 11437 6069 11471 6103
rect 14197 6069 14231 6103
rect 15209 6069 15243 6103
rect 15577 6069 15611 6103
rect 17325 6069 17359 6103
rect 18245 6069 18279 6103
rect 18705 6069 18739 6103
rect 20729 6069 20763 6103
rect 3709 5865 3743 5899
rect 4997 5865 5031 5899
rect 5457 5865 5491 5899
rect 8677 5865 8711 5899
rect 11069 5865 11103 5899
rect 12449 5865 12483 5899
rect 13093 5865 13127 5899
rect 19073 5865 19107 5899
rect 19809 5865 19843 5899
rect 2596 5797 2630 5831
rect 5365 5797 5399 5831
rect 6920 5797 6954 5831
rect 13820 5797 13854 5831
rect 6653 5729 6687 5763
rect 9945 5729 9979 5763
rect 13553 5729 13587 5763
rect 15485 5729 15519 5763
rect 15853 5729 15887 5763
rect 16037 5729 16071 5763
rect 16304 5729 16338 5763
rect 17601 5729 17635 5763
rect 17949 5729 17983 5763
rect 20177 5729 20211 5763
rect 2329 5661 2363 5695
rect 5549 5661 5583 5695
rect 8769 5661 8803 5695
rect 8953 5661 8987 5695
rect 9689 5661 9723 5695
rect 12541 5661 12575 5695
rect 12725 5661 12759 5695
rect 17693 5661 17727 5695
rect 19349 5661 19383 5695
rect 20269 5661 20303 5695
rect 20453 5661 20487 5695
rect 8033 5525 8067 5559
rect 8309 5525 8343 5559
rect 12081 5525 12115 5559
rect 14933 5525 14967 5559
rect 15669 5525 15703 5559
rect 17417 5525 17451 5559
rect 17601 5525 17635 5559
rect 8953 5321 8987 5355
rect 9229 5321 9263 5355
rect 12449 5321 12483 5355
rect 16037 5321 16071 5355
rect 16957 5321 16991 5355
rect 18613 5321 18647 5355
rect 21005 5321 21039 5355
rect 3341 5253 3375 5287
rect 5089 5253 5123 5287
rect 11069 5253 11103 5287
rect 11161 5253 11195 5287
rect 16589 5253 16623 5287
rect 18245 5253 18279 5287
rect 6009 5185 6043 5219
rect 7021 5185 7055 5219
rect 10793 5185 10827 5219
rect 11805 5185 11839 5219
rect 13093 5185 13127 5219
rect 14289 5185 14323 5219
rect 14657 5185 14691 5219
rect 17417 5185 17451 5219
rect 17509 5185 17543 5219
rect 19257 5185 19291 5219
rect 1961 5117 1995 5151
rect 3709 5117 3743 5151
rect 3965 5117 3999 5151
rect 5733 5117 5767 5151
rect 7573 5117 7607 5151
rect 9413 5117 9447 5151
rect 11069 5117 11103 5151
rect 11621 5117 11655 5151
rect 12909 5117 12943 5151
rect 16405 5117 16439 5151
rect 18061 5117 18095 5151
rect 19625 5117 19659 5151
rect 2228 5049 2262 5083
rect 7840 5049 7874 5083
rect 10517 5049 10551 5083
rect 10609 5049 10643 5083
rect 14105 5049 14139 5083
rect 14924 5049 14958 5083
rect 17325 5049 17359 5083
rect 19892 5049 19926 5083
rect 5365 4981 5399 5015
rect 5825 4981 5859 5015
rect 10149 4981 10183 5015
rect 11529 4981 11563 5015
rect 12817 4981 12851 5015
rect 13645 4981 13679 5015
rect 14013 4981 14047 5015
rect 18981 4981 19015 5015
rect 19073 4981 19107 5015
rect 2789 4777 2823 4811
rect 7021 4777 7055 4811
rect 8125 4777 8159 4811
rect 8493 4777 8527 4811
rect 9689 4777 9723 4811
rect 13093 4777 13127 4811
rect 16037 4777 16071 4811
rect 18521 4777 18555 4811
rect 20177 4777 20211 4811
rect 4804 4709 4838 4743
rect 8585 4709 8619 4743
rect 13820 4709 13854 4743
rect 16589 4709 16623 4743
rect 19042 4709 19076 4743
rect 1409 4641 1443 4675
rect 1676 4641 1710 4675
rect 4537 4641 4571 4675
rect 6929 4641 6963 4675
rect 10057 4641 10091 4675
rect 10885 4641 10919 4675
rect 11704 4641 11738 4675
rect 13553 4641 13587 4675
rect 15301 4641 15335 4675
rect 16037 4641 16071 4675
rect 16497 4641 16531 4675
rect 17141 4641 17175 4675
rect 17408 4641 17442 4675
rect 18797 4641 18831 4675
rect 7113 4573 7147 4607
rect 8677 4573 8711 4607
rect 10149 4573 10183 4607
rect 10241 4573 10275 4607
rect 11437 4573 11471 4607
rect 16773 4573 16807 4607
rect 16129 4505 16163 4539
rect 5917 4437 5951 4471
rect 6561 4437 6595 4471
rect 11069 4437 11103 4471
rect 12817 4437 12851 4471
rect 14933 4437 14967 4471
rect 15485 4437 15519 4471
rect 9229 4233 9263 4267
rect 19993 4233 20027 4267
rect 6837 4165 6871 4199
rect 16589 4165 16623 4199
rect 2605 4097 2639 4131
rect 2973 4097 3007 4131
rect 5273 4097 5307 4131
rect 6193 4097 6227 4131
rect 7481 4097 7515 4131
rect 13001 4097 13035 4131
rect 16037 4097 16071 4131
rect 17233 4097 17267 4131
rect 19533 4097 19567 4131
rect 20545 4097 20579 4131
rect 3240 4029 3274 4063
rect 5089 4029 5123 4063
rect 6009 4029 6043 4063
rect 7205 4029 7239 4063
rect 7849 4029 7883 4063
rect 10057 4029 10091 4063
rect 10324 4029 10358 4063
rect 11805 4029 11839 4063
rect 12817 4029 12851 4063
rect 12909 4029 12943 4063
rect 13829 4029 13863 4063
rect 14096 4029 14130 4063
rect 17049 4029 17083 4063
rect 18429 4029 18463 4063
rect 4997 3961 5031 3995
rect 6101 3961 6135 3995
rect 8116 3961 8150 3995
rect 15853 3961 15887 3995
rect 15945 3961 15979 3995
rect 16957 3961 16991 3995
rect 1961 3893 1995 3927
rect 2329 3893 2363 3927
rect 2421 3893 2455 3927
rect 4353 3893 4387 3927
rect 4629 3893 4663 3927
rect 5641 3893 5675 3927
rect 7297 3893 7331 3927
rect 11437 3893 11471 3927
rect 11989 3893 12023 3927
rect 12449 3893 12483 3927
rect 15209 3893 15243 3927
rect 15485 3893 15519 3927
rect 18613 3893 18647 3927
rect 18981 3893 19015 3927
rect 19349 3893 19383 3927
rect 19441 3893 19475 3927
rect 20361 3893 20395 3927
rect 20453 3893 20487 3927
rect 2605 3689 2639 3723
rect 4077 3689 4111 3723
rect 4537 3689 4571 3723
rect 5089 3689 5123 3723
rect 6377 3689 6411 3723
rect 13093 3689 13127 3723
rect 14197 3689 14231 3723
rect 14657 3689 14691 3723
rect 15117 3689 15151 3723
rect 15761 3689 15795 3723
rect 18613 3689 18647 3723
rect 18981 3689 19015 3723
rect 20913 3689 20947 3723
rect 4445 3621 4479 3655
rect 10324 3621 10358 3655
rect 13185 3621 13219 3655
rect 15669 3621 15703 3655
rect 16764 3621 16798 3655
rect 20085 3621 20119 3655
rect 2973 3553 3007 3587
rect 5457 3553 5491 3587
rect 7104 3553 7138 3587
rect 8861 3553 8895 3587
rect 8953 3553 8987 3587
rect 12081 3553 12115 3587
rect 13737 3553 13771 3587
rect 14565 3553 14599 3587
rect 15117 3553 15151 3587
rect 16497 3553 16531 3587
rect 19993 3553 20027 3587
rect 3065 3485 3099 3519
rect 3157 3485 3191 3519
rect 4629 3485 4663 3519
rect 5549 3485 5583 3519
rect 5733 3485 5767 3519
rect 6837 3485 6871 3519
rect 9045 3485 9079 3519
rect 10057 3485 10091 3519
rect 12173 3485 12207 3519
rect 12357 3485 12391 3519
rect 12541 3485 12575 3519
rect 13277 3485 13311 3519
rect 14841 3485 14875 3519
rect 15853 3485 15887 3519
rect 19073 3485 19107 3519
rect 19257 3485 19291 3519
rect 20177 3485 20211 3519
rect 11713 3417 11747 3451
rect 19625 3417 19659 3451
rect 8217 3349 8251 3383
rect 8493 3349 8527 3383
rect 11437 3349 11471 3383
rect 12541 3349 12575 3383
rect 12725 3349 12759 3383
rect 15301 3349 15335 3383
rect 17877 3349 17911 3383
rect 3157 3145 3191 3179
rect 5733 3145 5767 3179
rect 8217 3145 8251 3179
rect 8585 3145 8619 3179
rect 15945 3145 15979 3179
rect 16129 3145 16163 3179
rect 11989 3077 12023 3111
rect 3617 3009 3651 3043
rect 3801 3009 3835 3043
rect 4813 3009 4847 3043
rect 6193 3009 6227 3043
rect 6377 3009 6411 3043
rect 9045 3009 9079 3043
rect 9229 3009 9263 3043
rect 10057 3009 10091 3043
rect 13001 3009 13035 3043
rect 17325 3077 17359 3111
rect 20913 3077 20947 3111
rect 16589 3009 16623 3043
rect 16773 3009 16807 3043
rect 19257 3009 19291 3043
rect 20269 3009 20303 3043
rect 3525 2941 3559 2975
rect 4629 2941 4663 2975
rect 6101 2941 6135 2975
rect 6837 2941 6871 2975
rect 7104 2941 7138 2975
rect 10324 2941 10358 2975
rect 11805 2941 11839 2975
rect 12817 2941 12851 2975
rect 13461 2941 13495 2975
rect 13737 2941 13771 2975
rect 14197 2941 14231 2975
rect 14841 2941 14875 2975
rect 15577 2941 15611 2975
rect 15945 2941 15979 2975
rect 16497 2941 16531 2975
rect 17141 2941 17175 2975
rect 18061 2941 18095 2975
rect 20729 2941 20763 2975
rect 12909 2873 12943 2907
rect 15117 2873 15151 2907
rect 19073 2873 19107 2907
rect 20085 2873 20119 2907
rect 4169 2805 4203 2839
rect 4537 2805 4571 2839
rect 8953 2805 8987 2839
rect 11437 2805 11471 2839
rect 12449 2805 12483 2839
rect 14381 2805 14415 2839
rect 15761 2805 15795 2839
rect 18245 2805 18279 2839
rect 18705 2805 18739 2839
rect 19165 2805 19199 2839
rect 19717 2805 19751 2839
rect 20177 2805 20211 2839
rect 3525 2601 3559 2635
rect 8125 2601 8159 2635
rect 9781 2601 9815 2635
rect 10149 2601 10183 2635
rect 11345 2601 11379 2635
rect 11713 2601 11747 2635
rect 19073 2601 19107 2635
rect 10241 2533 10275 2567
rect 11805 2533 11839 2567
rect 12909 2533 12943 2567
rect 13645 2533 13679 2567
rect 15761 2533 15795 2567
rect 20453 2533 20487 2567
rect 8861 2465 8895 2499
rect 10793 2465 10827 2499
rect 12664 2465 12698 2499
rect 13277 2465 13311 2499
rect 13369 2465 13403 2499
rect 14105 2465 14139 2499
rect 14841 2465 14875 2499
rect 15485 2465 15519 2499
rect 16221 2465 16255 2499
rect 16957 2465 16991 2499
rect 17509 2465 17543 2499
rect 18337 2465 18371 2499
rect 19441 2465 19475 2499
rect 20177 2465 20211 2499
rect 8217 2397 8251 2431
rect 8309 2397 8343 2431
rect 9137 2397 9171 2431
rect 10425 2397 10459 2431
rect 11161 2397 11195 2431
rect 11897 2397 11931 2431
rect 7757 2261 7791 2295
rect 10977 2261 11011 2295
rect 11161 2261 11195 2295
rect 14381 2397 14415 2431
rect 16497 2397 16531 2431
rect 19533 2397 19567 2431
rect 19625 2397 19659 2431
rect 13277 2261 13311 2295
rect 15025 2261 15059 2295
rect 17141 2261 17175 2295
rect 17693 2261 17727 2295
rect 18521 2261 18555 2295
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 18690 19496 18696 19508
rect 18651 19468 18696 19496
rect 18690 19456 18696 19468
rect 18748 19456 18754 19508
rect 20714 19496 20720 19508
rect 20675 19468 20720 19496
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19261 1823 19295
rect 1765 19255 1823 19261
rect 2317 19295 2375 19301
rect 2317 19261 2329 19295
rect 2363 19292 2375 19295
rect 3418 19292 3424 19304
rect 2363 19264 3424 19292
rect 2363 19261 2375 19264
rect 2317 19255 2375 19261
rect 1780 19224 1808 19255
rect 3418 19252 3424 19264
rect 3476 19252 3482 19304
rect 17862 19252 17868 19304
rect 17920 19292 17926 19304
rect 18509 19295 18567 19301
rect 18509 19292 18521 19295
rect 17920 19264 18521 19292
rect 17920 19252 17926 19264
rect 18509 19261 18521 19264
rect 18555 19261 18567 19295
rect 20530 19292 20536 19304
rect 20491 19264 20536 19292
rect 18509 19255 18567 19261
rect 20530 19252 20536 19264
rect 20588 19252 20594 19304
rect 6730 19224 6736 19236
rect 1780 19196 6736 19224
rect 6730 19184 6736 19196
rect 6788 19184 6794 19236
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2774 19156 2780 19168
rect 2547 19128 2780 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2774 19116 2780 19128
rect 2832 19116 2838 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1946 18952 1952 18964
rect 1907 18924 1952 18952
rect 1946 18912 1952 18924
rect 2004 18912 2010 18964
rect 17862 18884 17868 18896
rect 17823 18856 17868 18884
rect 17862 18844 17868 18856
rect 17920 18844 17926 18896
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18816 1823 18819
rect 6178 18816 6184 18828
rect 1811 18788 6184 18816
rect 1811 18785 1823 18788
rect 1765 18779 1823 18785
rect 6178 18776 6184 18788
rect 6236 18776 6242 18828
rect 16666 18776 16672 18828
rect 16724 18816 16730 18828
rect 17589 18819 17647 18825
rect 17589 18816 17601 18819
rect 16724 18788 17601 18816
rect 16724 18776 16730 18788
rect 17589 18785 17601 18788
rect 17635 18785 17647 18819
rect 17589 18779 17647 18785
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 20714 18408 20720 18420
rect 20675 18380 20720 18408
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 20530 18204 20536 18216
rect 20491 18176 20536 18204
rect 20530 18164 20536 18176
rect 20588 18164 20594 18216
rect 16574 18096 16580 18148
rect 16632 18136 16638 18148
rect 18966 18136 18972 18148
rect 16632 18108 18972 18136
rect 16632 18096 16638 18108
rect 18966 18096 18972 18108
rect 19024 18096 19030 18148
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 2409 17799 2467 17805
rect 2409 17796 2421 17799
rect 1820 17768 2421 17796
rect 1820 17756 1826 17768
rect 2409 17765 2421 17768
rect 2455 17765 2467 17799
rect 2409 17759 2467 17765
rect 19889 17799 19947 17805
rect 19889 17765 19901 17799
rect 19935 17796 19947 17799
rect 20530 17796 20536 17808
rect 19935 17768 20536 17796
rect 19935 17765 19947 17768
rect 19889 17759 19947 17765
rect 20530 17756 20536 17768
rect 20588 17756 20594 17808
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17697 1639 17731
rect 1581 17691 1639 17697
rect 2133 17731 2191 17737
rect 2133 17697 2145 17731
rect 2179 17728 2191 17731
rect 6362 17728 6368 17740
rect 2179 17700 6368 17728
rect 2179 17697 2191 17700
rect 2133 17691 2191 17697
rect 1596 17660 1624 17691
rect 6362 17688 6368 17700
rect 6420 17688 6426 17740
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 19613 17731 19671 17737
rect 19613 17728 19625 17731
rect 17184 17700 19625 17728
rect 17184 17688 17190 17700
rect 19613 17697 19625 17700
rect 19659 17697 19671 17731
rect 19613 17691 19671 17697
rect 7374 17660 7380 17672
rect 1596 17632 7380 17660
rect 7374 17620 7380 17632
rect 7432 17620 7438 17672
rect 1670 17552 1676 17604
rect 1728 17592 1734 17604
rect 1765 17595 1823 17601
rect 1765 17592 1777 17595
rect 1728 17564 1777 17592
rect 1728 17552 1734 17564
rect 1765 17561 1777 17564
rect 1811 17561 1823 17595
rect 1765 17555 1823 17561
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 20162 17320 20168 17332
rect 20123 17292 20168 17320
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 20714 17320 20720 17332
rect 20675 17292 20720 17320
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17116 1823 17119
rect 7190 17116 7196 17128
rect 1811 17088 7196 17116
rect 1811 17085 1823 17088
rect 1765 17079 1823 17085
rect 7190 17076 7196 17088
rect 7248 17076 7254 17128
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 19981 17119 20039 17125
rect 19981 17116 19993 17119
rect 19392 17088 19993 17116
rect 19392 17076 19398 17088
rect 19981 17085 19993 17088
rect 20027 17085 20039 17119
rect 19981 17079 20039 17085
rect 20162 17076 20168 17128
rect 20220 17116 20226 17128
rect 20533 17119 20591 17125
rect 20533 17116 20545 17119
rect 20220 17088 20545 17116
rect 20220 17076 20226 17088
rect 20533 17085 20545 17088
rect 20579 17085 20591 17119
rect 20533 17079 20591 17085
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1854 16736 1860 16788
rect 1912 16776 1918 16788
rect 1949 16779 2007 16785
rect 1949 16776 1961 16779
rect 1912 16748 1961 16776
rect 1912 16736 1918 16748
rect 1949 16745 1961 16748
rect 1995 16745 2007 16779
rect 20438 16776 20444 16788
rect 20399 16748 20444 16776
rect 1949 16739 2007 16745
rect 20438 16736 20444 16748
rect 20496 16736 20502 16788
rect 1765 16643 1823 16649
rect 1765 16609 1777 16643
rect 1811 16640 1823 16643
rect 5810 16640 5816 16652
rect 1811 16612 5816 16640
rect 1811 16609 1823 16612
rect 1765 16603 1823 16609
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 20257 16643 20315 16649
rect 20257 16609 20269 16643
rect 20303 16640 20315 16643
rect 20622 16640 20628 16652
rect 20303 16612 20628 16640
rect 20303 16609 20315 16612
rect 20257 16603 20315 16609
rect 20622 16600 20628 16612
rect 20680 16600 20686 16652
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 3694 16232 3700 16244
rect 3655 16204 3700 16232
rect 3694 16192 3700 16204
rect 3752 16192 3758 16244
rect 14553 16235 14611 16241
rect 14553 16201 14565 16235
rect 14599 16232 14611 16235
rect 17954 16232 17960 16244
rect 14599 16204 17960 16232
rect 14599 16201 14611 16204
rect 14553 16195 14611 16201
rect 17954 16192 17960 16204
rect 18012 16192 18018 16244
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 16028 1823 16031
rect 3234 16028 3240 16040
rect 1811 16000 3240 16028
rect 1811 15997 1823 16000
rect 1765 15991 1823 15997
rect 3234 15988 3240 16000
rect 3292 15988 3298 16040
rect 3510 16028 3516 16040
rect 3471 16000 3516 16028
rect 3510 15988 3516 16000
rect 3568 15988 3574 16040
rect 13722 15988 13728 16040
rect 13780 16028 13786 16040
rect 14369 16031 14427 16037
rect 14369 16028 14381 16031
rect 13780 16000 14381 16028
rect 13780 15988 13786 16000
rect 14369 15997 14381 16000
rect 14415 15997 14427 16031
rect 20530 16028 20536 16040
rect 20491 16000 20536 16028
rect 14369 15991 14427 15997
rect 20530 15988 20536 16000
rect 20588 15988 20594 16040
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 2498 15688 2504 15700
rect 2459 15660 2504 15688
rect 2498 15648 2504 15660
rect 2556 15648 2562 15700
rect 19886 15688 19892 15700
rect 19847 15660 19892 15688
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 20254 15648 20260 15700
rect 20312 15688 20318 15700
rect 20441 15691 20499 15697
rect 20441 15688 20453 15691
rect 20312 15660 20453 15688
rect 20312 15648 20318 15660
rect 20441 15657 20453 15660
rect 20487 15657 20499 15691
rect 20441 15651 20499 15657
rect 3510 15580 3516 15632
rect 3568 15620 3574 15632
rect 4341 15623 4399 15629
rect 4341 15620 4353 15623
rect 3568 15592 4353 15620
rect 3568 15580 3574 15592
rect 4341 15589 4353 15592
rect 4387 15589 4399 15623
rect 13722 15620 13728 15632
rect 13683 15592 13728 15620
rect 4341 15583 4399 15589
rect 13722 15580 13728 15592
rect 13780 15580 13786 15632
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15552 1823 15555
rect 1854 15552 1860 15564
rect 1811 15524 1860 15552
rect 1811 15521 1823 15524
rect 1765 15515 1823 15521
rect 1854 15512 1860 15524
rect 1912 15512 1918 15564
rect 2317 15555 2375 15561
rect 2317 15521 2329 15555
rect 2363 15552 2375 15555
rect 3970 15552 3976 15564
rect 2363 15524 3976 15552
rect 2363 15521 2375 15524
rect 2317 15515 2375 15521
rect 3970 15512 3976 15524
rect 4028 15512 4034 15564
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4246 15552 4252 15564
rect 4111 15524 4252 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 13262 15512 13268 15564
rect 13320 15552 13326 15564
rect 13449 15555 13507 15561
rect 13449 15552 13461 15555
rect 13320 15524 13461 15552
rect 13320 15512 13326 15524
rect 13449 15521 13461 15524
rect 13495 15521 13507 15555
rect 13449 15515 13507 15521
rect 19426 15512 19432 15564
rect 19484 15552 19490 15564
rect 19705 15555 19763 15561
rect 19705 15552 19717 15555
rect 19484 15524 19717 15552
rect 19484 15512 19490 15524
rect 19705 15521 19717 15524
rect 19751 15521 19763 15555
rect 19705 15515 19763 15521
rect 19794 15512 19800 15564
rect 19852 15552 19858 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 19852 15524 20269 15552
rect 19852 15512 19858 15524
rect 20257 15521 20269 15524
rect 20303 15521 20315 15555
rect 20257 15515 20315 15521
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15144 2559 15147
rect 2774 15144 2780 15156
rect 2547 15116 2780 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 2774 15104 2780 15116
rect 2832 15104 2838 15156
rect 3050 15144 3056 15156
rect 3011 15116 3056 15144
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 3602 15144 3608 15156
rect 3563 15116 3608 15144
rect 3602 15104 3608 15116
rect 3660 15104 3666 15156
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 6181 15147 6239 15153
rect 6181 15144 6193 15147
rect 4120 15116 6193 15144
rect 4120 15104 4126 15116
rect 6181 15113 6193 15116
rect 6227 15113 6239 15147
rect 6181 15107 6239 15113
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 20717 15147 20775 15153
rect 20717 15144 20729 15147
rect 20404 15116 20729 15144
rect 20404 15104 20410 15116
rect 20717 15113 20729 15116
rect 20763 15113 20775 15147
rect 20717 15107 20775 15113
rect 1946 15076 1952 15088
rect 1907 15048 1952 15076
rect 1946 15036 1952 15048
rect 2004 15036 2010 15088
rect 11793 15079 11851 15085
rect 11793 15045 11805 15079
rect 11839 15076 11851 15079
rect 17954 15076 17960 15088
rect 11839 15048 17960 15076
rect 11839 15045 11851 15048
rect 11793 15039 11851 15045
rect 17954 15036 17960 15048
rect 18012 15036 18018 15088
rect 5626 15008 5632 15020
rect 2332 14980 5632 15008
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 2332 14949 2360 14980
rect 5626 14968 5632 14980
rect 5684 14968 5690 15020
rect 7558 15008 7564 15020
rect 5828 14980 7564 15008
rect 2317 14943 2375 14949
rect 2317 14909 2329 14943
rect 2363 14909 2375 14943
rect 2317 14903 2375 14909
rect 2869 14943 2927 14949
rect 2869 14909 2881 14943
rect 2915 14909 2927 14943
rect 2869 14903 2927 14909
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14940 3479 14943
rect 5828 14940 5856 14980
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 15008 14335 15011
rect 14366 15008 14372 15020
rect 14323 14980 14372 15008
rect 14323 14977 14335 14980
rect 14277 14971 14335 14977
rect 14366 14968 14372 14980
rect 14424 14968 14430 15020
rect 5994 14940 6000 14952
rect 3467 14912 5856 14940
rect 5955 14912 6000 14940
rect 3467 14909 3479 14912
rect 3421 14903 3479 14909
rect 2884 14872 2912 14903
rect 5994 14900 6000 14912
rect 6052 14900 6058 14952
rect 11606 14940 11612 14952
rect 11567 14912 11612 14940
rect 11606 14900 11612 14912
rect 11664 14900 11670 14952
rect 14093 14943 14151 14949
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 14458 14940 14464 14952
rect 14139 14912 14464 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 14458 14900 14464 14912
rect 14516 14940 14522 14952
rect 19334 14940 19340 14952
rect 14516 14912 19340 14940
rect 14516 14900 14522 14912
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 19429 14943 19487 14949
rect 19429 14909 19441 14943
rect 19475 14940 19487 14943
rect 19702 14940 19708 14952
rect 19475 14912 19708 14940
rect 19475 14909 19487 14912
rect 19429 14903 19487 14909
rect 19702 14900 19708 14912
rect 19760 14900 19766 14952
rect 19981 14943 20039 14949
rect 19981 14909 19993 14943
rect 20027 14940 20039 14943
rect 20438 14940 20444 14952
rect 20027 14912 20444 14940
rect 20027 14909 20039 14912
rect 19981 14903 20039 14909
rect 20438 14900 20444 14912
rect 20496 14900 20502 14952
rect 20533 14943 20591 14949
rect 20533 14909 20545 14943
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 5350 14872 5356 14884
rect 2884 14844 5356 14872
rect 5350 14832 5356 14844
rect 5408 14832 5414 14884
rect 17034 14832 17040 14884
rect 17092 14872 17098 14884
rect 20548 14872 20576 14903
rect 17092 14844 20576 14872
rect 17092 14832 17098 14844
rect 13630 14804 13636 14816
rect 13591 14776 13636 14804
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 13998 14804 14004 14816
rect 13959 14776 14004 14804
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 16942 14804 16948 14816
rect 16903 14776 16948 14804
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 19242 14764 19248 14816
rect 19300 14804 19306 14816
rect 19613 14807 19671 14813
rect 19613 14804 19625 14807
rect 19300 14776 19625 14804
rect 19300 14764 19306 14776
rect 19613 14773 19625 14776
rect 19659 14773 19671 14807
rect 19613 14767 19671 14773
rect 20165 14807 20223 14813
rect 20165 14773 20177 14807
rect 20211 14804 20223 14807
rect 20254 14804 20260 14816
rect 20211 14776 20260 14804
rect 20211 14773 20223 14776
rect 20165 14767 20223 14773
rect 20254 14764 20260 14776
rect 20312 14764 20318 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 9125 14603 9183 14609
rect 9125 14600 9137 14603
rect 7708 14572 9137 14600
rect 7708 14560 7714 14572
rect 9125 14569 9137 14572
rect 9171 14600 9183 14603
rect 16574 14600 16580 14612
rect 9171 14572 16580 14600
rect 9171 14569 9183 14572
rect 9125 14563 9183 14569
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 17497 14603 17555 14609
rect 17497 14569 17509 14603
rect 17543 14569 17555 14603
rect 19886 14600 19892 14612
rect 19847 14572 19892 14600
rect 17497 14563 17555 14569
rect 1762 14492 1768 14544
rect 1820 14532 1826 14544
rect 2133 14535 2191 14541
rect 2133 14532 2145 14535
rect 1820 14504 2145 14532
rect 1820 14492 1826 14504
rect 2133 14501 2145 14504
rect 2179 14501 2191 14535
rect 2133 14495 2191 14501
rect 2961 14535 3019 14541
rect 2961 14501 2973 14535
rect 3007 14532 3019 14535
rect 3050 14532 3056 14544
rect 3007 14504 3056 14532
rect 3007 14501 3019 14504
rect 2961 14495 3019 14501
rect 3050 14492 3056 14504
rect 3108 14492 3114 14544
rect 3142 14492 3148 14544
rect 3200 14492 3206 14544
rect 5994 14492 6000 14544
rect 6052 14532 6058 14544
rect 6641 14535 6699 14541
rect 6641 14532 6653 14535
rect 6052 14504 6653 14532
rect 6052 14492 6058 14504
rect 6641 14501 6653 14504
rect 6687 14501 6699 14535
rect 6641 14495 6699 14501
rect 7742 14492 7748 14544
rect 7800 14532 7806 14544
rect 7990 14535 8048 14541
rect 7990 14532 8002 14535
rect 7800 14504 8002 14532
rect 7800 14492 7806 14504
rect 7990 14501 8002 14504
rect 8036 14501 8048 14535
rect 7990 14495 8048 14501
rect 11146 14492 11152 14544
rect 11204 14532 11210 14544
rect 11578 14535 11636 14541
rect 11578 14532 11590 14535
rect 11204 14504 11590 14532
rect 11204 14492 11210 14504
rect 11578 14501 11590 14504
rect 11624 14501 11636 14535
rect 17512 14532 17540 14563
rect 19886 14560 19892 14572
rect 19944 14560 19950 14612
rect 19978 14560 19984 14612
rect 20036 14560 20042 14612
rect 20346 14560 20352 14612
rect 20404 14600 20410 14612
rect 20441 14603 20499 14609
rect 20441 14600 20453 14603
rect 20404 14572 20453 14600
rect 20404 14560 20410 14572
rect 20441 14569 20453 14572
rect 20487 14569 20499 14603
rect 20441 14563 20499 14569
rect 17586 14532 17592 14544
rect 17499 14504 17592 14532
rect 11578 14495 11636 14501
rect 17586 14492 17592 14504
rect 17644 14532 17650 14544
rect 18018 14535 18076 14541
rect 18018 14532 18030 14535
rect 17644 14504 18030 14532
rect 17644 14492 17650 14504
rect 18018 14501 18030 14504
rect 18064 14501 18076 14535
rect 19996 14532 20024 14560
rect 19996 14504 20392 14532
rect 18018 14495 18076 14501
rect 1857 14467 1915 14473
rect 1857 14433 1869 14467
rect 1903 14464 1915 14467
rect 2866 14464 2872 14476
rect 1903 14436 2872 14464
rect 1903 14433 1915 14436
rect 1857 14427 1915 14433
rect 2866 14424 2872 14436
rect 2924 14424 2930 14476
rect 3160 14464 3188 14492
rect 20364 14476 20392 14504
rect 4890 14464 4896 14476
rect 3068 14436 4896 14464
rect 3068 14405 3096 14436
rect 4890 14424 4896 14436
rect 4948 14424 4954 14476
rect 6365 14467 6423 14473
rect 6365 14433 6377 14467
rect 6411 14464 6423 14467
rect 7006 14464 7012 14476
rect 6411 14436 7012 14464
rect 6411 14433 6423 14436
rect 6365 14427 6423 14433
rect 7006 14424 7012 14436
rect 7064 14424 7070 14476
rect 10686 14464 10692 14476
rect 10647 14436 10692 14464
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 11333 14467 11391 14473
rect 11333 14433 11345 14467
rect 11379 14464 11391 14467
rect 12434 14464 12440 14476
rect 11379 14436 12440 14464
rect 11379 14433 11391 14436
rect 11333 14427 11391 14433
rect 12434 14424 12440 14436
rect 12492 14464 12498 14476
rect 12989 14467 13047 14473
rect 12989 14464 13001 14467
rect 12492 14436 13001 14464
rect 12492 14424 12498 14436
rect 12989 14433 13001 14436
rect 13035 14433 13047 14467
rect 13256 14467 13314 14473
rect 13256 14464 13268 14467
rect 12989 14427 13047 14433
rect 13096 14436 13268 14464
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14365 3111 14399
rect 3053 14359 3111 14365
rect 3145 14399 3203 14405
rect 3145 14365 3157 14399
rect 3191 14365 3203 14399
rect 3145 14359 3203 14365
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14365 7803 14399
rect 10778 14396 10784 14408
rect 10739 14368 10784 14396
rect 7745 14359 7803 14365
rect 2682 14288 2688 14340
rect 2740 14328 2746 14340
rect 3160 14328 3188 14359
rect 2740 14300 3188 14328
rect 2740 14288 2746 14300
rect 2222 14220 2228 14272
rect 2280 14260 2286 14272
rect 2593 14263 2651 14269
rect 2593 14260 2605 14263
rect 2280 14232 2605 14260
rect 2280 14220 2286 14232
rect 2593 14229 2605 14232
rect 2639 14229 2651 14263
rect 7760 14260 7788 14359
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 10873 14399 10931 14405
rect 10873 14365 10885 14399
rect 10919 14365 10931 14399
rect 13096 14396 13124 14436
rect 13256 14433 13268 14436
rect 13302 14464 13314 14467
rect 15102 14464 15108 14476
rect 13302 14436 15108 14464
rect 13302 14433 13314 14436
rect 13256 14427 13314 14433
rect 15102 14424 15108 14436
rect 15160 14424 15166 14476
rect 16390 14473 16396 14476
rect 16384 14427 16396 14473
rect 16448 14464 16454 14476
rect 19705 14467 19763 14473
rect 16448 14436 16484 14464
rect 16390 14424 16396 14427
rect 16448 14424 16454 14436
rect 19705 14433 19717 14467
rect 19751 14464 19763 14467
rect 19978 14464 19984 14476
rect 19751 14436 19984 14464
rect 19751 14433 19763 14436
rect 19705 14427 19763 14433
rect 19978 14424 19984 14436
rect 20036 14424 20042 14476
rect 20257 14467 20315 14473
rect 20257 14433 20269 14467
rect 20303 14433 20315 14467
rect 20257 14427 20315 14433
rect 10873 14359 10931 14365
rect 12728 14368 13124 14396
rect 10042 14288 10048 14340
rect 10100 14328 10106 14340
rect 10888 14328 10916 14359
rect 12728 14337 12756 14368
rect 15378 14356 15384 14408
rect 15436 14396 15442 14408
rect 16117 14399 16175 14405
rect 16117 14396 16129 14399
rect 15436 14368 16129 14396
rect 15436 14356 15442 14368
rect 16117 14365 16129 14368
rect 16163 14365 16175 14399
rect 17770 14396 17776 14408
rect 17731 14368 17776 14396
rect 16117 14359 16175 14365
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 18966 14356 18972 14408
rect 19024 14396 19030 14408
rect 20272 14396 20300 14427
rect 20346 14424 20352 14476
rect 20404 14424 20410 14476
rect 19024 14368 20300 14396
rect 19024 14356 19030 14368
rect 10100 14300 10916 14328
rect 12713 14331 12771 14337
rect 10100 14288 10106 14300
rect 12713 14297 12725 14331
rect 12759 14297 12771 14331
rect 12713 14291 12771 14297
rect 19886 14288 19892 14340
rect 19944 14328 19950 14340
rect 20162 14328 20168 14340
rect 19944 14300 20168 14328
rect 19944 14288 19950 14300
rect 20162 14288 20168 14300
rect 20220 14288 20226 14340
rect 8662 14260 8668 14272
rect 7760 14232 8668 14260
rect 2593 14223 2651 14229
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 10318 14260 10324 14272
rect 10279 14232 10324 14260
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 14366 14260 14372 14272
rect 14327 14232 14372 14260
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 18506 14220 18512 14272
rect 18564 14260 18570 14272
rect 19153 14263 19211 14269
rect 19153 14260 19165 14263
rect 18564 14232 19165 14260
rect 18564 14220 18570 14232
rect 19153 14229 19165 14232
rect 19199 14229 19211 14263
rect 19153 14223 19211 14229
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 2593 14059 2651 14065
rect 2593 14025 2605 14059
rect 2639 14056 2651 14059
rect 2774 14056 2780 14068
rect 2639 14028 2780 14056
rect 2639 14025 2651 14028
rect 2593 14019 2651 14025
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 6270 14056 6276 14068
rect 2976 14028 6276 14056
rect 2976 13988 3004 14028
rect 6270 14016 6276 14028
rect 6328 14016 6334 14068
rect 7006 14056 7012 14068
rect 6967 14028 7012 14056
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 16390 14016 16396 14068
rect 16448 14056 16454 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 16448 14028 16681 14056
rect 16448 14016 16454 14028
rect 16669 14025 16681 14028
rect 16715 14025 16727 14059
rect 16669 14019 16727 14025
rect 2424 13960 3004 13988
rect 10321 13991 10379 13997
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 1762 13852 1768 13864
rect 1719 13824 1768 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 2424 13861 2452 13960
rect 10321 13957 10333 13991
rect 10367 13988 10379 13991
rect 16945 13991 17003 13997
rect 10367 13960 11376 13988
rect 10367 13957 10379 13960
rect 10321 13951 10379 13957
rect 4062 13880 4068 13932
rect 4120 13920 4126 13932
rect 5169 13923 5227 13929
rect 5169 13920 5181 13923
rect 4120 13892 5181 13920
rect 4120 13880 4126 13892
rect 5169 13889 5181 13892
rect 5215 13889 5227 13923
rect 7650 13920 7656 13932
rect 7611 13892 7656 13920
rect 5169 13883 5227 13889
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 10962 13920 10968 13932
rect 10923 13892 10968 13920
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 2409 13855 2467 13861
rect 2409 13821 2421 13855
rect 2455 13821 2467 13855
rect 2409 13815 2467 13821
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13852 3019 13855
rect 4154 13852 4160 13864
rect 3007 13824 4160 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 7558 13812 7564 13864
rect 7616 13852 7622 13864
rect 7616 13824 8156 13852
rect 7616 13812 7622 13824
rect 3228 13787 3286 13793
rect 3228 13753 3240 13787
rect 3274 13784 3286 13787
rect 4062 13784 4068 13796
rect 3274 13756 4068 13784
rect 3274 13753 3286 13756
rect 3228 13747 3286 13753
rect 4062 13744 4068 13756
rect 4120 13744 4126 13796
rect 4985 13787 5043 13793
rect 4985 13753 4997 13787
rect 5031 13784 5043 13787
rect 5718 13784 5724 13796
rect 5031 13756 5724 13784
rect 5031 13753 5043 13756
rect 4985 13747 5043 13753
rect 5718 13744 5724 13756
rect 5776 13744 5782 13796
rect 7006 13744 7012 13796
rect 7064 13784 7070 13796
rect 8021 13787 8079 13793
rect 8021 13784 8033 13787
rect 7064 13756 8033 13784
rect 7064 13744 7070 13756
rect 8021 13753 8033 13756
rect 8067 13753 8079 13787
rect 8128 13784 8156 13824
rect 10318 13812 10324 13864
rect 10376 13852 10382 13864
rect 10689 13855 10747 13861
rect 10689 13852 10701 13855
rect 10376 13824 10701 13852
rect 10376 13812 10382 13824
rect 10689 13821 10701 13824
rect 10735 13821 10747 13855
rect 10689 13815 10747 13821
rect 10781 13855 10839 13861
rect 10781 13821 10793 13855
rect 10827 13852 10839 13855
rect 11238 13852 11244 13864
rect 10827 13824 11244 13852
rect 10827 13821 10839 13824
rect 10781 13815 10839 13821
rect 11238 13812 11244 13824
rect 11296 13812 11302 13864
rect 11348 13861 11376 13960
rect 16945 13957 16957 13991
rect 16991 13988 17003 13991
rect 20714 13988 20720 14000
rect 16991 13960 18092 13988
rect 16991 13957 17003 13960
rect 16945 13951 17003 13957
rect 11606 13920 11612 13932
rect 11567 13892 11612 13920
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 13998 13880 14004 13932
rect 14056 13920 14062 13932
rect 14461 13923 14519 13929
rect 14461 13920 14473 13923
rect 14056 13892 14473 13920
rect 14056 13880 14062 13892
rect 14461 13889 14473 13892
rect 14507 13889 14519 13923
rect 17586 13920 17592 13932
rect 17547 13892 17592 13920
rect 14461 13883 14519 13889
rect 17586 13880 17592 13892
rect 17644 13880 17650 13932
rect 11333 13855 11391 13861
rect 11333 13821 11345 13855
rect 11379 13821 11391 13855
rect 11333 13815 11391 13821
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12492 13824 12817 13852
rect 12492 13812 12498 13824
rect 12805 13821 12817 13824
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 13072 13855 13130 13861
rect 13072 13821 13084 13855
rect 13118 13852 13130 13855
rect 14366 13852 14372 13864
rect 13118 13824 14372 13852
rect 13118 13821 13130 13824
rect 13072 13815 13130 13821
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15378 13852 15384 13864
rect 15335 13824 15384 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 15556 13855 15614 13861
rect 15556 13821 15568 13855
rect 15602 13852 15614 13855
rect 15930 13852 15936 13864
rect 15602 13824 15936 13852
rect 15602 13821 15614 13824
rect 15556 13815 15614 13821
rect 15930 13812 15936 13824
rect 15988 13812 15994 13864
rect 18064 13861 18092 13960
rect 18984 13960 20720 13988
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18325 13855 18383 13861
rect 18325 13821 18337 13855
rect 18371 13852 18383 13855
rect 18782 13852 18788 13864
rect 18371 13824 18788 13852
rect 18371 13821 18383 13824
rect 18325 13815 18383 13821
rect 18782 13812 18788 13824
rect 18840 13812 18846 13864
rect 18984 13861 19012 13960
rect 20714 13948 20720 13960
rect 20772 13948 20778 14000
rect 19702 13920 19708 13932
rect 19663 13892 19708 13920
rect 19702 13880 19708 13892
rect 19760 13880 19766 13932
rect 20438 13920 20444 13932
rect 20399 13892 20444 13920
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 18969 13855 19027 13861
rect 18969 13821 18981 13855
rect 19015 13821 19027 13855
rect 18969 13815 19027 13821
rect 19242 13812 19248 13864
rect 19300 13852 19306 13864
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19300 13824 19533 13852
rect 19300 13812 19306 13824
rect 19521 13821 19533 13824
rect 19567 13821 19579 13855
rect 20257 13855 20315 13861
rect 20257 13852 20269 13855
rect 19521 13815 19579 13821
rect 19628 13824 20269 13852
rect 8128 13756 17908 13784
rect 8021 13747 8079 13753
rect 4338 13716 4344 13728
rect 4299 13688 4344 13716
rect 4338 13676 4344 13688
rect 4396 13676 4402 13728
rect 4614 13716 4620 13728
rect 4575 13688 4620 13716
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 5074 13676 5080 13728
rect 5132 13716 5138 13728
rect 5132 13688 5177 13716
rect 5132 13676 5138 13688
rect 6638 13676 6644 13728
rect 6696 13716 6702 13728
rect 7377 13719 7435 13725
rect 7377 13716 7389 13719
rect 6696 13688 7389 13716
rect 6696 13676 6702 13688
rect 7377 13685 7389 13688
rect 7423 13685 7435 13719
rect 7377 13679 7435 13685
rect 7466 13676 7472 13728
rect 7524 13716 7530 13728
rect 14182 13716 14188 13728
rect 7524 13688 7569 13716
rect 14143 13688 14188 13716
rect 7524 13676 7530 13688
rect 14182 13676 14188 13688
rect 14240 13676 14246 13728
rect 16758 13676 16764 13728
rect 16816 13716 16822 13728
rect 17313 13719 17371 13725
rect 17313 13716 17325 13719
rect 16816 13688 17325 13716
rect 16816 13676 16822 13688
rect 17313 13685 17325 13688
rect 17359 13685 17371 13719
rect 17313 13679 17371 13685
rect 17402 13676 17408 13728
rect 17460 13716 17466 13728
rect 17880 13716 17908 13756
rect 17954 13744 17960 13796
rect 18012 13784 18018 13796
rect 19628 13784 19656 13824
rect 20257 13821 20269 13824
rect 20303 13821 20315 13855
rect 20257 13815 20315 13821
rect 18012 13756 19656 13784
rect 18012 13744 18018 13756
rect 18874 13716 18880 13728
rect 17460 13688 17505 13716
rect 17880 13688 18880 13716
rect 17460 13676 17466 13688
rect 18874 13676 18880 13688
rect 18932 13676 18938 13728
rect 19150 13716 19156 13728
rect 19111 13688 19156 13716
rect 19150 13676 19156 13688
rect 19208 13676 19214 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 2961 13515 3019 13521
rect 2961 13512 2973 13515
rect 2924 13484 2973 13512
rect 2924 13472 2930 13484
rect 2961 13481 2973 13484
rect 3007 13481 3019 13515
rect 2961 13475 3019 13481
rect 3421 13515 3479 13521
rect 3421 13481 3433 13515
rect 3467 13512 3479 13515
rect 4614 13512 4620 13524
rect 3467 13484 4620 13512
rect 3467 13481 3479 13484
rect 3421 13475 3479 13481
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 6638 13512 6644 13524
rect 6599 13484 6644 13512
rect 6638 13472 6644 13484
rect 6696 13472 6702 13524
rect 7006 13512 7012 13524
rect 6967 13484 7012 13512
rect 7006 13472 7012 13484
rect 7064 13472 7070 13524
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 7653 13515 7711 13521
rect 7653 13512 7665 13515
rect 7524 13484 7665 13512
rect 7524 13472 7530 13484
rect 7653 13481 7665 13484
rect 7699 13481 7711 13515
rect 7653 13475 7711 13481
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 11149 13515 11207 13521
rect 11149 13512 11161 13515
rect 11020 13484 11161 13512
rect 11020 13472 11026 13484
rect 11149 13481 11161 13484
rect 11195 13481 11207 13515
rect 11149 13475 11207 13481
rect 11238 13472 11244 13524
rect 11296 13512 11302 13524
rect 11425 13515 11483 13521
rect 11425 13512 11437 13515
rect 11296 13484 11437 13512
rect 11296 13472 11302 13484
rect 11425 13481 11437 13484
rect 11471 13481 11483 13515
rect 11425 13475 11483 13481
rect 12897 13515 12955 13521
rect 12897 13481 12909 13515
rect 12943 13512 12955 13515
rect 13630 13512 13636 13524
rect 12943 13484 13636 13512
rect 12943 13481 12955 13484
rect 12897 13475 12955 13481
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 15565 13515 15623 13521
rect 15565 13481 15577 13515
rect 15611 13481 15623 13515
rect 15565 13475 15623 13481
rect 16577 13515 16635 13521
rect 16577 13481 16589 13515
rect 16623 13512 16635 13515
rect 16758 13512 16764 13524
rect 16623 13484 16764 13512
rect 16623 13481 16635 13484
rect 16577 13475 16635 13481
rect 2317 13447 2375 13453
rect 2317 13413 2329 13447
rect 2363 13444 2375 13447
rect 3510 13444 3516 13456
rect 2363 13416 3516 13444
rect 2363 13413 2375 13416
rect 2317 13407 2375 13413
rect 3510 13404 3516 13416
rect 3568 13404 3574 13456
rect 4338 13404 4344 13456
rect 4396 13453 4402 13456
rect 4396 13447 4460 13453
rect 4396 13413 4414 13447
rect 4448 13413 4460 13447
rect 4396 13407 4460 13413
rect 8113 13447 8171 13453
rect 8113 13413 8125 13447
rect 8159 13444 8171 13447
rect 8202 13444 8208 13456
rect 8159 13416 8208 13444
rect 8159 13413 8171 13416
rect 8113 13407 8171 13413
rect 4396 13404 4402 13407
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 8294 13404 8300 13456
rect 8352 13444 8358 13456
rect 12802 13444 12808 13456
rect 8352 13416 12808 13444
rect 8352 13404 8358 13416
rect 12802 13404 12808 13416
rect 12860 13404 12866 13456
rect 12986 13444 12992 13456
rect 12947 13416 12992 13444
rect 12986 13404 12992 13416
rect 13044 13404 13050 13456
rect 13446 13404 13452 13456
rect 13504 13444 13510 13456
rect 13808 13447 13866 13453
rect 13808 13444 13820 13447
rect 13504 13416 13820 13444
rect 13504 13404 13510 13416
rect 13808 13413 13820 13416
rect 13854 13444 13866 13447
rect 14182 13444 14188 13456
rect 13854 13416 14188 13444
rect 13854 13413 13866 13416
rect 13808 13407 13866 13413
rect 14182 13404 14188 13416
rect 14240 13404 14246 13456
rect 15580 13444 15608 13475
rect 16758 13472 16764 13484
rect 16816 13472 16822 13524
rect 16942 13512 16948 13524
rect 16903 13484 16948 13512
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 17034 13472 17040 13524
rect 17092 13512 17098 13524
rect 17092 13484 17137 13512
rect 17092 13472 17098 13484
rect 18874 13472 18880 13524
rect 18932 13512 18938 13524
rect 20257 13515 20315 13521
rect 20257 13512 20269 13515
rect 18932 13484 20269 13512
rect 18932 13472 18938 13484
rect 20257 13481 20269 13484
rect 20303 13481 20315 13515
rect 20257 13475 20315 13481
rect 17402 13444 17408 13456
rect 15580 13416 17408 13444
rect 17402 13404 17408 13416
rect 17460 13404 17466 13456
rect 18132 13447 18190 13453
rect 18132 13413 18144 13447
rect 18178 13444 18190 13447
rect 18506 13444 18512 13456
rect 18178 13416 18512 13444
rect 18178 13413 18190 13416
rect 18132 13407 18190 13413
rect 18506 13404 18512 13416
rect 18564 13404 18570 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13345 1455 13379
rect 1397 13339 1455 13345
rect 1412 13240 1440 13339
rect 2038 13336 2044 13388
rect 2096 13376 2102 13388
rect 3329 13379 3387 13385
rect 3329 13376 3341 13379
rect 2096 13348 3341 13376
rect 2096 13336 2102 13348
rect 3329 13345 3341 13348
rect 3375 13345 3387 13379
rect 4356 13376 4384 13404
rect 3329 13339 3387 13345
rect 3620 13348 4384 13376
rect 8021 13379 8079 13385
rect 2314 13268 2320 13320
rect 2372 13308 2378 13320
rect 2409 13311 2467 13317
rect 2409 13308 2421 13311
rect 2372 13280 2421 13308
rect 2372 13268 2378 13280
rect 2409 13277 2421 13280
rect 2455 13277 2467 13311
rect 2590 13308 2596 13320
rect 2551 13280 2596 13308
rect 2409 13271 2467 13277
rect 2590 13268 2596 13280
rect 2648 13268 2654 13320
rect 3620 13317 3648 13348
rect 8021 13345 8033 13379
rect 8067 13376 8079 13379
rect 8754 13376 8760 13388
rect 8067 13348 8760 13376
rect 8067 13345 8079 13348
rect 8021 13339 8079 13345
rect 8754 13336 8760 13348
rect 8812 13336 8818 13388
rect 10042 13385 10048 13388
rect 10036 13376 10048 13385
rect 10003 13348 10048 13376
rect 10036 13339 10048 13348
rect 10100 13376 10106 13388
rect 11790 13376 11796 13388
rect 10100 13348 10804 13376
rect 11751 13348 11796 13376
rect 10042 13336 10048 13339
rect 10100 13336 10106 13348
rect 3605 13311 3663 13317
rect 3605 13277 3617 13311
rect 3651 13277 3663 13311
rect 4154 13308 4160 13320
rect 4115 13280 4160 13308
rect 3605 13271 3663 13277
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 7101 13311 7159 13317
rect 7101 13308 7113 13311
rect 7024 13280 7113 13308
rect 7024 13252 7052 13280
rect 7101 13277 7113 13280
rect 7147 13277 7159 13311
rect 7101 13271 7159 13277
rect 7285 13311 7343 13317
rect 7285 13277 7297 13311
rect 7331 13308 7343 13311
rect 7742 13308 7748 13320
rect 7331 13280 7748 13308
rect 7331 13277 7343 13280
rect 7285 13271 7343 13277
rect 7742 13268 7748 13280
rect 7800 13308 7806 13320
rect 8205 13311 8263 13317
rect 8205 13308 8217 13311
rect 7800 13280 8217 13308
rect 7800 13268 7806 13280
rect 8205 13277 8217 13280
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 8662 13268 8668 13320
rect 8720 13308 8726 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 8720 13280 9781 13308
rect 8720 13268 8726 13280
rect 9769 13277 9781 13280
rect 9815 13277 9827 13311
rect 10776 13308 10804 13348
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 11885 13379 11943 13385
rect 11885 13345 11897 13379
rect 11931 13376 11943 13379
rect 12894 13376 12900 13388
rect 11931 13348 12900 13376
rect 11931 13345 11943 13348
rect 11885 13339 11943 13345
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 13541 13379 13599 13385
rect 13541 13376 13553 13379
rect 13004 13348 13553 13376
rect 11977 13311 12035 13317
rect 11977 13308 11989 13311
rect 10776 13280 11989 13308
rect 9769 13271 9827 13277
rect 11977 13277 11989 13280
rect 12023 13277 12035 13311
rect 11977 13271 12035 13277
rect 12434 13268 12440 13320
rect 12492 13308 12498 13320
rect 13004 13308 13032 13348
rect 13541 13345 13553 13348
rect 13587 13345 13599 13379
rect 13541 13339 13599 13345
rect 15286 13336 15292 13388
rect 15344 13376 15350 13388
rect 15933 13379 15991 13385
rect 15933 13376 15945 13379
rect 15344 13348 15945 13376
rect 15344 13336 15350 13348
rect 15933 13345 15945 13348
rect 15979 13345 15991 13379
rect 15933 13339 15991 13345
rect 16025 13379 16083 13385
rect 16025 13345 16037 13379
rect 16071 13376 16083 13379
rect 16298 13376 16304 13388
rect 16071 13348 16304 13376
rect 16071 13345 16083 13348
rect 16025 13339 16083 13345
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 20162 13376 20168 13388
rect 20123 13348 20168 13376
rect 20162 13336 20168 13348
rect 20220 13336 20226 13388
rect 12492 13280 13032 13308
rect 13173 13311 13231 13317
rect 12492 13268 12498 13280
rect 13173 13277 13185 13311
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 16209 13311 16267 13317
rect 16209 13277 16221 13311
rect 16255 13308 16267 13311
rect 16390 13308 16396 13320
rect 16255 13280 16396 13308
rect 16255 13277 16267 13280
rect 16209 13271 16267 13277
rect 3326 13240 3332 13252
rect 1412 13212 3332 13240
rect 3326 13200 3332 13212
rect 3384 13200 3390 13252
rect 7006 13200 7012 13252
rect 7064 13200 7070 13252
rect 13188 13240 13216 13271
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 17129 13311 17187 13317
rect 17129 13277 17141 13311
rect 17175 13277 17187 13311
rect 17129 13271 17187 13277
rect 13446 13240 13452 13252
rect 13188 13212 13452 13240
rect 13446 13200 13452 13212
rect 13504 13200 13510 13252
rect 16408 13240 16436 13268
rect 17144 13240 17172 13271
rect 17770 13268 17776 13320
rect 17828 13308 17834 13320
rect 17865 13311 17923 13317
rect 17865 13308 17877 13311
rect 17828 13280 17877 13308
rect 17828 13268 17834 13280
rect 17865 13277 17877 13280
rect 17911 13277 17923 13311
rect 17865 13271 17923 13277
rect 16408 13212 17172 13240
rect 1949 13175 2007 13181
rect 1949 13141 1961 13175
rect 1995 13172 2007 13175
rect 2130 13172 2136 13184
rect 1995 13144 2136 13172
rect 1995 13141 2007 13144
rect 1949 13135 2007 13141
rect 2130 13132 2136 13144
rect 2188 13132 2194 13184
rect 5534 13172 5540 13184
rect 5495 13144 5540 13172
rect 5534 13132 5540 13144
rect 5592 13132 5598 13184
rect 6086 13132 6092 13184
rect 6144 13172 6150 13184
rect 11146 13172 11152 13184
rect 6144 13144 11152 13172
rect 6144 13132 6150 13144
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 12529 13175 12587 13181
rect 12529 13141 12541 13175
rect 12575 13172 12587 13175
rect 14274 13172 14280 13184
rect 12575 13144 14280 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 14918 13172 14924 13184
rect 14879 13144 14924 13172
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 16758 13132 16764 13184
rect 16816 13172 16822 13184
rect 17126 13172 17132 13184
rect 16816 13144 17132 13172
rect 16816 13132 16822 13144
rect 17126 13132 17132 13144
rect 17184 13132 17190 13184
rect 17880 13172 17908 13271
rect 20346 13268 20352 13320
rect 20404 13308 20410 13320
rect 20404 13280 20449 13308
rect 20404 13268 20410 13280
rect 18598 13172 18604 13184
rect 17880 13144 18604 13172
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 19150 13132 19156 13184
rect 19208 13172 19214 13184
rect 19245 13175 19303 13181
rect 19245 13172 19257 13175
rect 19208 13144 19257 13172
rect 19208 13132 19214 13144
rect 19245 13141 19257 13144
rect 19291 13141 19303 13175
rect 19245 13135 19303 13141
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 19797 13175 19855 13181
rect 19797 13172 19809 13175
rect 19392 13144 19809 13172
rect 19392 13132 19398 13144
rect 19797 13141 19809 13144
rect 19843 13141 19855 13175
rect 19797 13135 19855 13141
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1765 12971 1823 12977
rect 1765 12937 1777 12971
rect 1811 12968 1823 12971
rect 2038 12968 2044 12980
rect 1811 12940 2044 12968
rect 1811 12937 1823 12940
rect 1765 12931 1823 12937
rect 2038 12928 2044 12940
rect 2096 12928 2102 12980
rect 4062 12968 4068 12980
rect 2792 12940 4068 12968
rect 2222 12832 2228 12844
rect 2183 12804 2228 12832
rect 2222 12792 2228 12804
rect 2280 12792 2286 12844
rect 2409 12835 2467 12841
rect 2409 12801 2421 12835
rect 2455 12832 2467 12835
rect 2792 12832 2820 12940
rect 4062 12928 4068 12940
rect 4120 12968 4126 12980
rect 4157 12971 4215 12977
rect 4157 12968 4169 12971
rect 4120 12940 4169 12968
rect 4120 12928 4126 12940
rect 4157 12937 4169 12940
rect 4203 12937 4215 12971
rect 4157 12931 4215 12937
rect 4709 12971 4767 12977
rect 4709 12937 4721 12971
rect 4755 12968 4767 12971
rect 5074 12968 5080 12980
rect 4755 12940 5080 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 5718 12968 5724 12980
rect 5679 12940 5724 12968
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 7800 12940 8217 12968
rect 7800 12928 7806 12940
rect 8205 12937 8217 12940
rect 8251 12937 8263 12971
rect 10042 12968 10048 12980
rect 10003 12940 10048 12968
rect 8205 12931 8263 12937
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 13909 12971 13967 12977
rect 13909 12937 13921 12971
rect 13955 12968 13967 12971
rect 17954 12968 17960 12980
rect 13955 12940 17960 12968
rect 13955 12937 13967 12940
rect 13909 12931 13967 12937
rect 17954 12928 17960 12940
rect 18012 12928 18018 12980
rect 18874 12928 18880 12980
rect 18932 12968 18938 12980
rect 20257 12971 20315 12977
rect 18932 12940 20208 12968
rect 18932 12928 18938 12940
rect 12897 12903 12955 12909
rect 12897 12869 12909 12903
rect 12943 12900 12955 12903
rect 12943 12872 14412 12900
rect 12943 12869 12955 12872
rect 12897 12863 12955 12869
rect 2455 12804 2820 12832
rect 4617 12835 4675 12841
rect 2455 12801 2467 12804
rect 2409 12795 2467 12801
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 5353 12835 5411 12841
rect 5353 12832 5365 12835
rect 4663 12804 5365 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 5353 12801 5365 12804
rect 5399 12832 5411 12835
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 5399 12804 6377 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 6365 12801 6377 12804
rect 6411 12832 6423 12835
rect 6454 12832 6460 12844
rect 6411 12804 6460 12832
rect 6411 12801 6423 12804
rect 6365 12795 6423 12801
rect 6454 12792 6460 12804
rect 6512 12792 6518 12844
rect 8662 12832 8668 12844
rect 8623 12804 8668 12832
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 10410 12792 10416 12844
rect 10468 12832 10474 12844
rect 10689 12835 10747 12841
rect 10689 12832 10701 12835
rect 10468 12804 10701 12832
rect 10468 12792 10474 12804
rect 10689 12801 10701 12804
rect 10735 12801 10747 12835
rect 13446 12832 13452 12844
rect 13407 12804 13452 12832
rect 10689 12795 10747 12801
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 14384 12841 14412 12872
rect 16482 12860 16488 12912
rect 16540 12900 16546 12912
rect 16945 12903 17003 12909
rect 16945 12900 16957 12903
rect 16540 12872 16957 12900
rect 16540 12860 16546 12872
rect 16945 12869 16957 12872
rect 16991 12869 17003 12903
rect 16945 12863 17003 12869
rect 14369 12835 14427 12841
rect 14369 12801 14381 12835
rect 14415 12801 14427 12835
rect 14369 12795 14427 12801
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12832 14611 12835
rect 14918 12832 14924 12844
rect 14599 12804 14924 12832
rect 14599 12801 14611 12804
rect 14553 12795 14611 12801
rect 14918 12792 14924 12804
rect 14976 12832 14982 12844
rect 17497 12835 17555 12841
rect 17497 12832 17509 12835
rect 14976 12804 15424 12832
rect 14976 12792 14982 12804
rect 2130 12764 2136 12776
rect 2091 12736 2136 12764
rect 2130 12724 2136 12736
rect 2188 12724 2194 12776
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12764 2835 12767
rect 2866 12764 2872 12776
rect 2823 12736 2872 12764
rect 2823 12733 2835 12736
rect 2777 12727 2835 12733
rect 2866 12724 2872 12736
rect 2924 12764 2930 12776
rect 4154 12764 4160 12776
rect 2924 12736 4160 12764
rect 2924 12724 2930 12736
rect 4154 12724 4160 12736
rect 4212 12724 4218 12776
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5258 12764 5264 12776
rect 5123 12736 5264 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 6086 12764 6092 12776
rect 6047 12736 6092 12764
rect 6086 12724 6092 12736
rect 6144 12724 6150 12776
rect 6638 12724 6644 12776
rect 6696 12764 6702 12776
rect 10962 12773 10968 12776
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6696 12736 6837 12764
rect 6696 12724 6702 12736
rect 6825 12733 6837 12736
rect 6871 12733 6883 12767
rect 10956 12764 10968 12773
rect 6825 12727 6883 12733
rect 6932 12736 10824 12764
rect 10923 12736 10968 12764
rect 3044 12699 3102 12705
rect 3044 12665 3056 12699
rect 3090 12665 3102 12699
rect 3044 12659 3102 12665
rect 2590 12588 2596 12640
rect 2648 12628 2654 12640
rect 3059 12628 3087 12659
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 6932 12696 6960 12736
rect 4120 12668 6960 12696
rect 7092 12699 7150 12705
rect 4120 12656 4126 12668
rect 7092 12665 7104 12699
rect 7138 12696 7150 12699
rect 7282 12696 7288 12708
rect 7138 12668 7288 12696
rect 7138 12665 7150 12668
rect 7092 12659 7150 12665
rect 7282 12656 7288 12668
rect 7340 12656 7346 12708
rect 8932 12699 8990 12705
rect 8932 12665 8944 12699
rect 8978 12696 8990 12699
rect 10226 12696 10232 12708
rect 8978 12668 10232 12696
rect 8978 12665 8990 12668
rect 8932 12659 8990 12665
rect 10226 12656 10232 12668
rect 10284 12656 10290 12708
rect 10796 12696 10824 12736
rect 10956 12727 10968 12736
rect 10962 12724 10968 12727
rect 11020 12724 11026 12776
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12764 13323 12767
rect 13906 12764 13912 12776
rect 13311 12736 13912 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 13906 12724 13912 12736
rect 13964 12724 13970 12776
rect 14274 12764 14280 12776
rect 14235 12736 14280 12764
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12733 15347 12767
rect 15396 12764 15424 12804
rect 16316 12804 17509 12832
rect 15545 12767 15603 12773
rect 15545 12764 15557 12767
rect 15396 12736 15557 12764
rect 15289 12727 15347 12733
rect 15545 12733 15557 12736
rect 15591 12733 15603 12767
rect 15545 12727 15603 12733
rect 12894 12696 12900 12708
rect 10796 12668 12900 12696
rect 12894 12656 12900 12668
rect 12952 12656 12958 12708
rect 15304 12696 15332 12727
rect 15378 12696 15384 12708
rect 15304 12668 15384 12696
rect 15378 12656 15384 12668
rect 15436 12656 15442 12708
rect 4617 12631 4675 12637
rect 4617 12628 4629 12631
rect 2648 12600 4629 12628
rect 2648 12588 2654 12600
rect 4617 12597 4629 12600
rect 4663 12597 4675 12631
rect 5166 12628 5172 12640
rect 5127 12600 5172 12628
rect 4617 12591 4675 12597
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 6181 12631 6239 12637
rect 6181 12597 6193 12631
rect 6227 12628 6239 12631
rect 7742 12628 7748 12640
rect 6227 12600 7748 12628
rect 6227 12597 6239 12600
rect 6181 12591 6239 12597
rect 7742 12588 7748 12600
rect 7800 12628 7806 12640
rect 8478 12628 8484 12640
rect 7800 12600 8484 12628
rect 7800 12588 7806 12600
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 12069 12631 12127 12637
rect 12069 12597 12081 12631
rect 12115 12628 12127 12631
rect 13170 12628 13176 12640
rect 12115 12600 13176 12628
rect 12115 12597 12127 12600
rect 12069 12591 12127 12597
rect 13170 12588 13176 12600
rect 13228 12588 13234 12640
rect 13357 12631 13415 12637
rect 13357 12597 13369 12631
rect 13403 12628 13415 12631
rect 13814 12628 13820 12640
rect 13403 12600 13820 12628
rect 13403 12597 13415 12600
rect 13357 12591 13415 12597
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 15102 12588 15108 12640
rect 15160 12628 15166 12640
rect 16316 12628 16344 12804
rect 17497 12801 17509 12804
rect 17543 12801 17555 12835
rect 17497 12795 17555 12801
rect 18046 12764 18052 12776
rect 18007 12736 18052 12764
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 18598 12724 18604 12776
rect 18656 12764 18662 12776
rect 19150 12773 19156 12776
rect 18877 12767 18935 12773
rect 18877 12764 18889 12767
rect 18656 12736 18889 12764
rect 18656 12724 18662 12736
rect 18877 12733 18889 12736
rect 18923 12733 18935 12767
rect 19144 12764 19156 12773
rect 19111 12736 19156 12764
rect 18877 12727 18935 12733
rect 19144 12727 19156 12736
rect 19150 12724 19156 12727
rect 19208 12724 19214 12776
rect 20180 12764 20208 12940
rect 20257 12937 20269 12971
rect 20303 12968 20315 12971
rect 20346 12968 20352 12980
rect 20303 12940 20352 12968
rect 20303 12937 20315 12940
rect 20257 12931 20315 12937
rect 20346 12928 20352 12940
rect 20404 12928 20410 12980
rect 20714 12832 20720 12844
rect 20675 12804 20720 12832
rect 20714 12792 20720 12804
rect 20772 12792 20778 12844
rect 20438 12764 20444 12776
rect 20180 12736 20444 12764
rect 20438 12724 20444 12736
rect 20496 12724 20502 12776
rect 20533 12767 20591 12773
rect 20533 12733 20545 12767
rect 20579 12733 20591 12767
rect 20533 12727 20591 12733
rect 17586 12696 17592 12708
rect 16684 12668 17592 12696
rect 16684 12637 16712 12668
rect 17586 12656 17592 12668
rect 17644 12656 17650 12708
rect 18325 12699 18383 12705
rect 18325 12665 18337 12699
rect 18371 12665 18383 12699
rect 18325 12659 18383 12665
rect 15160 12600 16344 12628
rect 16669 12631 16727 12637
rect 15160 12588 15166 12600
rect 16669 12597 16681 12631
rect 16715 12597 16727 12631
rect 17310 12628 17316 12640
rect 17271 12600 17316 12628
rect 16669 12591 16727 12597
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 18340 12628 18368 12659
rect 18690 12656 18696 12708
rect 18748 12696 18754 12708
rect 20548 12696 20576 12727
rect 18748 12668 20576 12696
rect 18748 12656 18754 12668
rect 20714 12628 20720 12640
rect 17460 12600 17505 12628
rect 18340 12600 20720 12628
rect 17460 12588 17466 12600
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 1670 12424 1676 12436
rect 1631 12396 1676 12424
rect 1670 12384 1676 12396
rect 1728 12384 1734 12436
rect 2409 12427 2467 12433
rect 2409 12393 2421 12427
rect 2455 12424 2467 12427
rect 3050 12424 3056 12436
rect 2455 12396 3056 12424
rect 2455 12393 2467 12396
rect 2409 12387 2467 12393
rect 3050 12384 3056 12396
rect 3108 12424 3114 12436
rect 3694 12424 3700 12436
rect 3108 12396 3700 12424
rect 3108 12384 3114 12396
rect 3694 12384 3700 12396
rect 3752 12384 3758 12436
rect 4065 12427 4123 12433
rect 4065 12393 4077 12427
rect 4111 12393 4123 12427
rect 4065 12387 4123 12393
rect 2498 12356 2504 12368
rect 2411 12328 2504 12356
rect 2498 12316 2504 12328
rect 2556 12356 2562 12368
rect 3326 12356 3332 12368
rect 2556 12328 3188 12356
rect 3287 12328 3332 12356
rect 2556 12316 2562 12328
rect 1489 12291 1547 12297
rect 1489 12257 1501 12291
rect 1535 12288 1547 12291
rect 1854 12288 1860 12300
rect 1535 12260 1860 12288
rect 1535 12257 1547 12260
rect 1489 12251 1547 12257
rect 1854 12248 1860 12260
rect 1912 12248 1918 12300
rect 3050 12288 3056 12300
rect 3011 12260 3056 12288
rect 3050 12248 3056 12260
rect 3108 12248 3114 12300
rect 3160 12288 3188 12328
rect 3326 12316 3332 12328
rect 3384 12316 3390 12368
rect 4080 12356 4108 12387
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4433 12427 4491 12433
rect 4433 12424 4445 12427
rect 4212 12396 4445 12424
rect 4212 12384 4218 12396
rect 4433 12393 4445 12396
rect 4479 12393 4491 12427
rect 4433 12387 4491 12393
rect 4522 12384 4528 12436
rect 4580 12424 4586 12436
rect 6454 12424 6460 12436
rect 4580 12396 5304 12424
rect 6415 12396 6460 12424
rect 4580 12384 4586 12396
rect 5166 12356 5172 12368
rect 4080 12328 4476 12356
rect 4338 12288 4344 12300
rect 3160 12260 4344 12288
rect 4338 12248 4344 12260
rect 4396 12248 4402 12300
rect 4448 12288 4476 12328
rect 4632 12328 5172 12356
rect 4632 12288 4660 12328
rect 5166 12316 5172 12328
rect 5224 12316 5230 12368
rect 5276 12356 5304 12396
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 6733 12427 6791 12433
rect 6733 12393 6745 12427
rect 6779 12424 6791 12427
rect 7006 12424 7012 12436
rect 6779 12396 7012 12424
rect 6779 12393 6791 12396
rect 6733 12387 6791 12393
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 7929 12427 7987 12433
rect 7929 12393 7941 12427
rect 7975 12424 7987 12427
rect 8202 12424 8208 12436
rect 7975 12396 8208 12424
rect 7975 12393 7987 12396
rect 7929 12387 7987 12393
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 10045 12427 10103 12433
rect 10045 12424 10057 12427
rect 8536 12396 10057 12424
rect 8536 12384 8542 12396
rect 10045 12393 10057 12396
rect 10091 12393 10103 12427
rect 10045 12387 10103 12393
rect 10689 12427 10747 12433
rect 10689 12393 10701 12427
rect 10735 12424 10747 12427
rect 10778 12424 10784 12436
rect 10735 12396 10784 12424
rect 10735 12393 10747 12396
rect 10689 12387 10747 12393
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 14185 12427 14243 12433
rect 14185 12424 14197 12427
rect 13872 12396 14197 12424
rect 13872 12384 13878 12396
rect 14185 12393 14197 12396
rect 14231 12393 14243 12427
rect 14185 12387 14243 12393
rect 14553 12427 14611 12433
rect 14553 12393 14565 12427
rect 14599 12424 14611 12427
rect 16482 12424 16488 12436
rect 14599 12396 16488 12424
rect 14599 12393 14611 12396
rect 14553 12387 14611 12393
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 17865 12427 17923 12433
rect 17865 12393 17877 12427
rect 17911 12424 17923 12427
rect 18046 12424 18052 12436
rect 17911 12396 18052 12424
rect 17911 12393 17923 12396
rect 17865 12387 17923 12393
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 18138 12384 18144 12436
rect 18196 12424 18202 12436
rect 19978 12424 19984 12436
rect 18196 12396 19984 12424
rect 18196 12384 18202 12396
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 20622 12384 20628 12436
rect 20680 12384 20686 12436
rect 7193 12359 7251 12365
rect 7193 12356 7205 12359
rect 5276 12328 7205 12356
rect 7193 12325 7205 12328
rect 7239 12325 7251 12359
rect 7193 12319 7251 12325
rect 8297 12359 8355 12365
rect 8297 12325 8309 12359
rect 8343 12356 8355 12359
rect 8343 12328 8524 12356
rect 8343 12325 8355 12328
rect 8297 12319 8355 12325
rect 8496 12300 8524 12328
rect 9214 12316 9220 12368
rect 9272 12356 9278 12368
rect 10594 12356 10600 12368
rect 9272 12328 10600 12356
rect 9272 12316 9278 12328
rect 10594 12316 10600 12328
rect 10652 12316 10658 12368
rect 14826 12316 14832 12368
rect 14884 12356 14890 12368
rect 17126 12356 17132 12368
rect 14884 12328 17132 12356
rect 14884 12316 14890 12328
rect 17126 12316 17132 12328
rect 17184 12356 17190 12368
rect 17313 12359 17371 12365
rect 17313 12356 17325 12359
rect 17184 12328 17325 12356
rect 17184 12316 17190 12328
rect 17313 12325 17325 12328
rect 17359 12325 17371 12359
rect 18506 12356 18512 12368
rect 17313 12319 17371 12325
rect 17512 12328 18512 12356
rect 5333 12291 5391 12297
rect 5333 12288 5345 12291
rect 4448 12260 4660 12288
rect 4724 12260 5345 12288
rect 4724 12232 4752 12260
rect 5333 12257 5345 12260
rect 5379 12257 5391 12291
rect 5333 12251 5391 12257
rect 6454 12248 6460 12300
rect 6512 12288 6518 12300
rect 7101 12291 7159 12297
rect 7101 12288 7113 12291
rect 6512 12260 7113 12288
rect 6512 12248 6518 12260
rect 7101 12257 7113 12260
rect 7147 12257 7159 12291
rect 7101 12251 7159 12257
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 8386 12288 8392 12300
rect 7432 12260 8392 12288
rect 7432 12248 7438 12260
rect 8386 12248 8392 12260
rect 8444 12248 8450 12300
rect 8478 12248 8484 12300
rect 8536 12248 8542 12300
rect 8662 12248 8668 12300
rect 8720 12288 8726 12300
rect 8849 12291 8907 12297
rect 8849 12288 8861 12291
rect 8720 12260 8861 12288
rect 8720 12248 8726 12260
rect 8849 12257 8861 12260
rect 8895 12257 8907 12291
rect 8849 12251 8907 12257
rect 8938 12248 8944 12300
rect 8996 12288 9002 12300
rect 9125 12291 9183 12297
rect 9125 12288 9137 12291
rect 8996 12260 9137 12288
rect 8996 12248 9002 12260
rect 9125 12257 9137 12260
rect 9171 12257 9183 12291
rect 10137 12291 10195 12297
rect 10137 12288 10149 12291
rect 9125 12251 9183 12257
rect 9232 12260 10149 12288
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12189 2743 12223
rect 2685 12183 2743 12189
rect 2700 12152 2728 12183
rect 3234 12180 3240 12232
rect 3292 12220 3298 12232
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 3292 12192 4537 12220
rect 3292 12180 3298 12192
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 4706 12220 4712 12232
rect 4619 12192 4712 12220
rect 4525 12183 4583 12189
rect 2774 12152 2780 12164
rect 2700 12124 2780 12152
rect 2774 12112 2780 12124
rect 2832 12112 2838 12164
rect 4540 12152 4568 12183
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 5074 12220 5080 12232
rect 5035 12192 5080 12220
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 8202 12220 8208 12232
rect 7340 12192 8208 12220
rect 7340 12180 7346 12192
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 8570 12220 8576 12232
rect 8531 12192 8576 12220
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 4798 12152 4804 12164
rect 4540 12124 4804 12152
rect 4798 12112 4804 12124
rect 4856 12112 4862 12164
rect 9232 12152 9260 12260
rect 10137 12257 10149 12260
rect 10183 12257 10195 12291
rect 10137 12251 10195 12257
rect 11057 12291 11115 12297
rect 11057 12257 11069 12291
rect 11103 12288 11115 12291
rect 12066 12288 12072 12300
rect 11103 12260 12072 12288
rect 11103 12257 11115 12260
rect 11057 12251 11115 12257
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 12437 12291 12495 12297
rect 12437 12257 12449 12291
rect 12483 12288 12495 12291
rect 12710 12288 12716 12300
rect 12483 12260 12716 12288
rect 12483 12257 12495 12260
rect 12437 12251 12495 12257
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 12897 12291 12955 12297
rect 12897 12257 12909 12291
rect 12943 12288 12955 12291
rect 13541 12291 13599 12297
rect 13541 12288 13553 12291
rect 12943 12260 13553 12288
rect 12943 12257 12955 12260
rect 12897 12251 12955 12257
rect 13541 12257 13553 12260
rect 13587 12257 13599 12291
rect 13541 12251 13599 12257
rect 14366 12248 14372 12300
rect 14424 12288 14430 12300
rect 15657 12291 15715 12297
rect 14424 12260 14872 12288
rect 14424 12248 14430 12260
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 10042 12220 10048 12232
rect 9456 12192 10048 12220
rect 9456 12180 9462 12192
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10226 12220 10232 12232
rect 10187 12192 10232 12220
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 11146 12220 11152 12232
rect 11107 12192 11152 12220
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 11333 12223 11391 12229
rect 11333 12189 11345 12223
rect 11379 12220 11391 12223
rect 11517 12223 11575 12229
rect 11517 12220 11529 12223
rect 11379 12192 11529 12220
rect 11379 12189 11391 12192
rect 11333 12183 11391 12189
rect 11517 12189 11529 12192
rect 11563 12189 11575 12223
rect 11698 12220 11704 12232
rect 11659 12192 11704 12220
rect 11517 12183 11575 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 12618 12180 12624 12232
rect 12676 12220 12682 12232
rect 12989 12223 13047 12229
rect 12989 12220 13001 12223
rect 12676 12192 13001 12220
rect 12676 12180 12682 12192
rect 12989 12189 13001 12192
rect 13035 12189 13047 12223
rect 13170 12220 13176 12232
rect 13083 12192 13176 12220
rect 12989 12183 13047 12189
rect 13170 12180 13176 12192
rect 13228 12220 13234 12232
rect 13446 12220 13452 12232
rect 13228 12192 13452 12220
rect 13228 12180 13234 12192
rect 13446 12180 13452 12192
rect 13504 12180 13510 12232
rect 14642 12220 14648 12232
rect 14603 12192 14648 12220
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 14844 12229 14872 12260
rect 15657 12257 15669 12291
rect 15703 12288 15715 12291
rect 16022 12288 16028 12300
rect 15703 12260 16028 12288
rect 15703 12257 15715 12260
rect 15657 12251 15715 12257
rect 16022 12248 16028 12260
rect 16080 12248 16086 12300
rect 16942 12248 16948 12300
rect 17000 12288 17006 12300
rect 17221 12291 17279 12297
rect 17221 12288 17233 12291
rect 17000 12260 17233 12288
rect 17000 12248 17006 12260
rect 17221 12257 17233 12260
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 15286 12180 15292 12232
rect 15344 12220 15350 12232
rect 15749 12223 15807 12229
rect 15749 12220 15761 12223
rect 15344 12192 15761 12220
rect 15344 12180 15350 12192
rect 15749 12189 15761 12192
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 15933 12223 15991 12229
rect 15933 12189 15945 12223
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 6012 12124 9260 12152
rect 9677 12155 9735 12161
rect 2041 12087 2099 12093
rect 2041 12053 2053 12087
rect 2087 12084 2099 12087
rect 3418 12084 3424 12096
rect 2087 12056 3424 12084
rect 2087 12053 2099 12056
rect 2041 12047 2099 12053
rect 3418 12044 3424 12056
rect 3476 12044 3482 12096
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 3786 12084 3792 12096
rect 3660 12056 3792 12084
rect 3660 12044 3666 12056
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 4982 12044 4988 12096
rect 5040 12084 5046 12096
rect 5258 12084 5264 12096
rect 5040 12056 5264 12084
rect 5040 12044 5046 12056
rect 5258 12044 5264 12056
rect 5316 12084 5322 12096
rect 6012 12084 6040 12124
rect 9677 12121 9689 12155
rect 9723 12152 9735 12155
rect 11790 12152 11796 12164
rect 9723 12124 11796 12152
rect 9723 12121 9735 12124
rect 9677 12115 9735 12121
rect 11790 12112 11796 12124
rect 11848 12112 11854 12164
rect 15948 12152 15976 12183
rect 16206 12180 16212 12232
rect 16264 12220 16270 12232
rect 17402 12220 17408 12232
rect 16264 12192 17408 12220
rect 16264 12180 16270 12192
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 17512 12229 17540 12328
rect 18506 12316 18512 12328
rect 18564 12316 18570 12368
rect 17954 12248 17960 12300
rect 18012 12288 18018 12300
rect 18233 12291 18291 12297
rect 18233 12288 18245 12291
rect 18012 12260 18245 12288
rect 18012 12248 18018 12260
rect 18233 12257 18245 12260
rect 18279 12257 18291 12291
rect 19150 12288 19156 12300
rect 18233 12251 18291 12257
rect 18524 12260 19156 12288
rect 18524 12229 18552 12260
rect 19150 12248 19156 12260
rect 19208 12248 19214 12300
rect 19981 12291 20039 12297
rect 19981 12257 19993 12291
rect 20027 12288 20039 12291
rect 20027 12260 20208 12288
rect 20027 12257 20039 12260
rect 19981 12251 20039 12257
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12189 17555 12223
rect 17497 12183 17555 12189
rect 18325 12223 18383 12229
rect 18325 12189 18337 12223
rect 18371 12189 18383 12223
rect 18325 12183 18383 12189
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12189 18567 12223
rect 18874 12220 18880 12232
rect 18835 12192 18880 12220
rect 18509 12183 18567 12189
rect 16482 12152 16488 12164
rect 11900 12124 16488 12152
rect 8846 12084 8852 12096
rect 5316 12056 6040 12084
rect 8759 12056 8852 12084
rect 5316 12044 5322 12056
rect 8846 12044 8852 12056
rect 8904 12084 8910 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8904 12056 8953 12084
rect 8904 12044 8910 12056
rect 8941 12053 8953 12056
rect 8987 12053 8999 12087
rect 8941 12047 8999 12053
rect 10226 12044 10232 12096
rect 10284 12084 10290 12096
rect 11054 12084 11060 12096
rect 10284 12056 11060 12084
rect 10284 12044 10290 12056
rect 11054 12044 11060 12056
rect 11112 12084 11118 12096
rect 11517 12087 11575 12093
rect 11517 12084 11529 12087
rect 11112 12056 11529 12084
rect 11112 12044 11118 12056
rect 11517 12053 11529 12056
rect 11563 12084 11575 12087
rect 11900 12084 11928 12124
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 16853 12155 16911 12161
rect 16853 12121 16865 12155
rect 16899 12152 16911 12155
rect 18340 12152 18368 12183
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 19794 12152 19800 12164
rect 16899 12124 18368 12152
rect 19444 12124 19800 12152
rect 16899 12121 16911 12124
rect 16853 12115 16911 12121
rect 19444 12096 19472 12124
rect 19794 12112 19800 12124
rect 19852 12152 19858 12164
rect 20088 12152 20116 12183
rect 19852 12124 20116 12152
rect 19852 12112 19858 12124
rect 11563 12056 11928 12084
rect 12253 12087 12311 12093
rect 11563 12053 11575 12056
rect 11517 12047 11575 12053
rect 12253 12053 12265 12087
rect 12299 12084 12311 12087
rect 12342 12084 12348 12096
rect 12299 12056 12348 12084
rect 12299 12053 12311 12056
rect 12253 12047 12311 12053
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 12526 12084 12532 12096
rect 12487 12056 12532 12084
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 15289 12087 15347 12093
rect 15289 12084 15301 12087
rect 13136 12056 15301 12084
rect 13136 12044 13142 12056
rect 15289 12053 15301 12056
rect 15335 12053 15347 12087
rect 15289 12047 15347 12053
rect 15746 12044 15752 12096
rect 15804 12084 15810 12096
rect 17218 12084 17224 12096
rect 15804 12056 17224 12084
rect 15804 12044 15810 12056
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 19426 12084 19432 12096
rect 19387 12056 19432 12084
rect 19426 12044 19432 12056
rect 19484 12044 19490 12096
rect 19518 12044 19524 12096
rect 19576 12084 19582 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19576 12056 19625 12084
rect 19576 12044 19582 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 20180 12084 20208 12260
rect 20257 12223 20315 12229
rect 20257 12189 20269 12223
rect 20303 12220 20315 12223
rect 20530 12220 20536 12232
rect 20303 12192 20536 12220
rect 20303 12189 20315 12192
rect 20257 12183 20315 12189
rect 20530 12180 20536 12192
rect 20588 12180 20594 12232
rect 20438 12112 20444 12164
rect 20496 12152 20502 12164
rect 20640 12152 20668 12384
rect 20496 12124 20668 12152
rect 20496 12112 20502 12124
rect 20898 12084 20904 12096
rect 20180 12056 20904 12084
rect 19613 12047 19671 12053
rect 20898 12044 20904 12056
rect 20956 12044 20962 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 4706 11880 4712 11892
rect 4028 11852 4292 11880
rect 4667 11852 4712 11880
rect 4028 11840 4034 11852
rect 1949 11815 2007 11821
rect 1949 11781 1961 11815
rect 1995 11812 2007 11815
rect 3326 11812 3332 11824
rect 1995 11784 3332 11812
rect 1995 11781 2007 11784
rect 1949 11775 2007 11781
rect 3326 11772 3332 11784
rect 3384 11772 3390 11824
rect 4264 11812 4292 11852
rect 4706 11840 4712 11852
rect 4764 11840 4770 11892
rect 4816 11852 8064 11880
rect 4816 11812 4844 11852
rect 4264 11784 4844 11812
rect 8036 11812 8064 11852
rect 8202 11840 8208 11892
rect 8260 11880 8266 11892
rect 8481 11883 8539 11889
rect 8481 11880 8493 11883
rect 8260 11852 8493 11880
rect 8260 11840 8266 11852
rect 8481 11849 8493 11852
rect 8527 11880 8539 11883
rect 8570 11880 8576 11892
rect 8527 11852 8576 11880
rect 8527 11849 8539 11852
rect 8481 11843 8539 11849
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 8754 11880 8760 11892
rect 8715 11852 8760 11880
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 10502 11880 10508 11892
rect 9088 11852 10508 11880
rect 9088 11840 9094 11852
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 10686 11880 10692 11892
rect 10647 11852 10692 11880
rect 10686 11840 10692 11852
rect 10744 11840 10750 11892
rect 11146 11840 11152 11892
rect 11204 11880 11210 11892
rect 11790 11880 11796 11892
rect 11204 11852 11796 11880
rect 11204 11840 11210 11852
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 12437 11883 12495 11889
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 12483 11852 13124 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 10594 11812 10600 11824
rect 8036 11784 10600 11812
rect 10594 11772 10600 11784
rect 10652 11772 10658 11824
rect 11054 11772 11060 11824
rect 11112 11812 11118 11824
rect 13096 11812 13124 11852
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 13449 11883 13507 11889
rect 13449 11880 13461 11883
rect 13412 11852 13461 11880
rect 13412 11840 13418 11852
rect 13449 11849 13461 11852
rect 13495 11849 13507 11883
rect 15286 11880 15292 11892
rect 15247 11852 15292 11880
rect 13449 11843 13507 11849
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 15654 11840 15660 11892
rect 15712 11880 15718 11892
rect 16206 11880 16212 11892
rect 15712 11852 16212 11880
rect 15712 11840 15718 11852
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 16482 11840 16488 11892
rect 16540 11880 16546 11892
rect 17681 11883 17739 11889
rect 17681 11880 17693 11883
rect 16540 11852 17693 11880
rect 16540 11840 16546 11852
rect 17681 11849 17693 11852
rect 17727 11849 17739 11883
rect 17681 11843 17739 11849
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 18049 11883 18107 11889
rect 18049 11880 18061 11883
rect 18012 11852 18061 11880
rect 18012 11840 18018 11852
rect 18049 11849 18061 11852
rect 18095 11849 18107 11883
rect 18049 11843 18107 11849
rect 20530 11840 20536 11892
rect 20588 11880 20594 11892
rect 20993 11883 21051 11889
rect 20993 11880 21005 11883
rect 20588 11852 21005 11880
rect 20588 11840 20594 11852
rect 20993 11849 21005 11852
rect 21039 11849 21051 11883
rect 20993 11843 21051 11849
rect 11112 11784 11284 11812
rect 13096 11784 13492 11812
rect 11112 11772 11118 11784
rect 2590 11744 2596 11756
rect 2551 11716 2596 11744
rect 2590 11704 2596 11716
rect 2648 11744 2654 11756
rect 2774 11744 2780 11756
rect 2648 11716 2780 11744
rect 2648 11704 2654 11716
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 5721 11747 5779 11753
rect 5721 11744 5733 11747
rect 5592 11716 5733 11744
rect 5592 11704 5598 11716
rect 5721 11713 5733 11716
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7156 11716 7201 11744
rect 7156 11704 7162 11716
rect 8570 11704 8576 11756
rect 8628 11744 8634 11756
rect 11256 11753 11284 11784
rect 13464 11756 13492 11784
rect 17402 11772 17408 11824
rect 17460 11812 17466 11824
rect 18138 11812 18144 11824
rect 17460 11784 18144 11812
rect 17460 11772 17466 11784
rect 18138 11772 18144 11784
rect 18196 11772 18202 11824
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 8628 11716 9321 11744
rect 8628 11704 8634 11716
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 9309 11707 9367 11713
rect 11241 11747 11299 11753
rect 11241 11713 11253 11747
rect 11287 11713 11299 11747
rect 12894 11744 12900 11756
rect 12855 11716 12900 11744
rect 11241 11707 11299 11713
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 12986 11704 12992 11756
rect 13044 11744 13050 11756
rect 13044 11716 13089 11744
rect 13044 11704 13050 11716
rect 13446 11704 13452 11756
rect 13504 11704 13510 11756
rect 14093 11747 14151 11753
rect 14093 11713 14105 11747
rect 14139 11744 14151 11747
rect 14366 11744 14372 11756
rect 14139 11716 14372 11744
rect 14139 11713 14151 11716
rect 14093 11707 14151 11713
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 15194 11744 15200 11756
rect 14700 11716 15200 11744
rect 14700 11704 14706 11716
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 15746 11744 15752 11756
rect 15707 11716 15752 11744
rect 15746 11704 15752 11716
rect 15804 11704 15810 11756
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11744 15991 11747
rect 15979 11716 16436 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 16408 11688 16436 11716
rect 18506 11704 18512 11756
rect 18564 11744 18570 11756
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 18564 11716 18613 11744
rect 18564 11704 18570 11716
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 2958 11636 2964 11688
rect 3016 11676 3022 11688
rect 3142 11676 3148 11688
rect 3016 11648 3148 11676
rect 3016 11636 3022 11648
rect 3142 11636 3148 11648
rect 3200 11676 3206 11688
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 3200 11648 3341 11676
rect 3200 11636 3206 11648
rect 3329 11645 3341 11648
rect 3375 11645 3387 11679
rect 3329 11639 3387 11645
rect 4062 11636 4068 11688
rect 4120 11676 4126 11688
rect 9030 11676 9036 11688
rect 4120 11648 9036 11676
rect 4120 11636 4126 11648
rect 9030 11636 9036 11648
rect 9088 11636 9094 11688
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11676 9275 11679
rect 9950 11676 9956 11688
rect 9263 11648 9956 11676
rect 9263 11645 9275 11648
rect 9217 11639 9275 11645
rect 9950 11636 9956 11648
rect 10008 11676 10014 11688
rect 10962 11676 10968 11688
rect 10008 11648 10968 11676
rect 10008 11636 10014 11648
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 11698 11676 11704 11688
rect 11103 11648 11704 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 16301 11679 16359 11685
rect 16301 11645 16313 11679
rect 16347 11645 16359 11679
rect 16301 11639 16359 11645
rect 2317 11611 2375 11617
rect 2317 11577 2329 11611
rect 2363 11608 2375 11611
rect 2866 11608 2872 11620
rect 2363 11580 2872 11608
rect 2363 11577 2375 11580
rect 2317 11571 2375 11577
rect 2866 11568 2872 11580
rect 2924 11568 2930 11620
rect 3234 11568 3240 11620
rect 3292 11608 3298 11620
rect 3574 11611 3632 11617
rect 3574 11608 3586 11611
rect 3292 11580 3586 11608
rect 3292 11568 3298 11580
rect 3574 11577 3586 11580
rect 3620 11577 3632 11611
rect 3574 11571 3632 11577
rect 5350 11568 5356 11620
rect 5408 11608 5414 11620
rect 5537 11611 5595 11617
rect 5537 11608 5549 11611
rect 5408 11580 5549 11608
rect 5408 11568 5414 11580
rect 5537 11577 5549 11580
rect 5583 11577 5595 11611
rect 5537 11571 5595 11577
rect 5629 11611 5687 11617
rect 5629 11577 5641 11611
rect 5675 11608 5687 11611
rect 5810 11608 5816 11620
rect 5675 11580 5816 11608
rect 5675 11577 5687 11580
rect 5629 11571 5687 11577
rect 5810 11568 5816 11580
rect 5868 11568 5874 11620
rect 7346 11611 7404 11617
rect 7346 11608 7358 11611
rect 7116 11580 7358 11608
rect 7116 11552 7144 11580
rect 7346 11577 7358 11580
rect 7392 11577 7404 11611
rect 7346 11571 7404 11577
rect 9125 11611 9183 11617
rect 9125 11577 9137 11611
rect 9171 11608 9183 11611
rect 11885 11611 11943 11617
rect 9171 11580 11836 11608
rect 9171 11577 9183 11580
rect 9125 11571 9183 11577
rect 2409 11543 2467 11549
rect 2409 11509 2421 11543
rect 2455 11540 2467 11543
rect 3786 11540 3792 11552
rect 2455 11512 3792 11540
rect 2455 11509 2467 11512
rect 2409 11503 2467 11509
rect 3786 11500 3792 11512
rect 3844 11500 3850 11552
rect 5169 11543 5227 11549
rect 5169 11509 5181 11543
rect 5215 11540 5227 11543
rect 5258 11540 5264 11552
rect 5215 11512 5264 11540
rect 5215 11509 5227 11512
rect 5169 11503 5227 11509
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 7098 11500 7104 11552
rect 7156 11500 7162 11552
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 10778 11540 10784 11552
rect 8444 11512 10784 11540
rect 8444 11500 8450 11512
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 11146 11540 11152 11552
rect 11107 11512 11152 11540
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 11808 11540 11836 11580
rect 11885 11577 11897 11611
rect 11931 11608 11943 11611
rect 12805 11611 12863 11617
rect 12805 11608 12817 11611
rect 11931 11580 12817 11608
rect 11931 11577 11943 11580
rect 11885 11571 11943 11577
rect 12805 11577 12817 11580
rect 12851 11577 12863 11611
rect 13909 11611 13967 11617
rect 13909 11608 13921 11611
rect 12805 11571 12863 11577
rect 13087 11580 13921 11608
rect 12894 11540 12900 11552
rect 11808 11512 12900 11540
rect 12894 11500 12900 11512
rect 12952 11540 12958 11552
rect 13087 11540 13115 11580
rect 13909 11577 13921 11580
rect 13955 11577 13967 11611
rect 13909 11571 13967 11577
rect 12952 11512 13115 11540
rect 13817 11543 13875 11549
rect 12952 11500 12958 11512
rect 13817 11509 13829 11543
rect 13863 11540 13875 11543
rect 14090 11540 14096 11552
rect 13863 11512 14096 11540
rect 13863 11509 13875 11512
rect 13817 11503 13875 11509
rect 14090 11500 14096 11512
rect 14148 11540 14154 11552
rect 15010 11540 15016 11552
rect 14148 11512 15016 11540
rect 14148 11500 14154 11512
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 15654 11540 15660 11552
rect 15615 11512 15660 11540
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 16316 11540 16344 11639
rect 16390 11636 16396 11688
rect 16448 11636 16454 11688
rect 18417 11679 18475 11685
rect 18417 11645 18429 11679
rect 18463 11676 18475 11679
rect 18874 11676 18880 11688
rect 18463 11648 18880 11676
rect 18463 11645 18475 11648
rect 18417 11639 18475 11645
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 19613 11679 19671 11685
rect 19613 11645 19625 11679
rect 19659 11676 19671 11679
rect 19702 11676 19708 11688
rect 19659 11648 19708 11676
rect 19659 11645 19671 11648
rect 19613 11639 19671 11645
rect 19702 11636 19708 11648
rect 19760 11636 19766 11688
rect 19880 11679 19938 11685
rect 19880 11645 19892 11679
rect 19926 11676 19938 11679
rect 20254 11676 20260 11688
rect 19926 11648 20260 11676
rect 19926 11645 19938 11648
rect 19880 11639 19938 11645
rect 20254 11636 20260 11648
rect 20312 11636 20318 11688
rect 16574 11617 16580 11620
rect 16568 11571 16580 11617
rect 16632 11608 16638 11620
rect 16850 11608 16856 11620
rect 16632 11580 16856 11608
rect 16574 11568 16580 11571
rect 16632 11568 16638 11580
rect 16850 11568 16856 11580
rect 16908 11568 16914 11620
rect 18509 11611 18567 11617
rect 18509 11577 18521 11611
rect 18555 11608 18567 11611
rect 18966 11608 18972 11620
rect 18555 11580 18972 11608
rect 18555 11577 18567 11580
rect 18509 11571 18567 11577
rect 18966 11568 18972 11580
rect 19024 11568 19030 11620
rect 16482 11540 16488 11552
rect 16316 11512 16488 11540
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 19426 11540 19432 11552
rect 17092 11512 19432 11540
rect 17092 11500 17098 11512
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 2041 11339 2099 11345
rect 2041 11305 2053 11339
rect 2087 11336 2099 11339
rect 3050 11336 3056 11348
rect 2087 11308 3056 11336
rect 2087 11305 2099 11308
rect 2041 11299 2099 11305
rect 3050 11296 3056 11308
rect 3108 11296 3114 11348
rect 5258 11336 5264 11348
rect 5219 11308 5264 11336
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 6362 11296 6368 11348
rect 6420 11336 6426 11348
rect 6457 11339 6515 11345
rect 6457 11336 6469 11339
rect 6420 11308 6469 11336
rect 6420 11296 6426 11308
rect 6457 11305 6469 11308
rect 6503 11305 6515 11339
rect 6457 11299 6515 11305
rect 7558 11296 7564 11348
rect 7616 11336 7622 11348
rect 7837 11339 7895 11345
rect 7837 11336 7849 11339
rect 7616 11308 7849 11336
rect 7616 11296 7622 11308
rect 7837 11305 7849 11308
rect 7883 11305 7895 11339
rect 7837 11299 7895 11305
rect 8573 11339 8631 11345
rect 8573 11305 8585 11339
rect 8619 11336 8631 11339
rect 10045 11339 10103 11345
rect 10045 11336 10057 11339
rect 8619 11308 10057 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 10045 11305 10057 11308
rect 10091 11305 10103 11339
rect 10045 11299 10103 11305
rect 10962 11296 10968 11348
rect 11020 11336 11026 11348
rect 12529 11339 12587 11345
rect 11020 11308 11560 11336
rect 11020 11296 11026 11308
rect 1394 11228 1400 11280
rect 1452 11268 1458 11280
rect 3329 11271 3387 11277
rect 3329 11268 3341 11271
rect 1452 11240 3341 11268
rect 1452 11228 1458 11240
rect 3329 11237 3341 11240
rect 3375 11237 3387 11271
rect 3329 11231 3387 11237
rect 4154 11228 4160 11280
rect 4212 11268 4218 11280
rect 9033 11271 9091 11277
rect 9033 11268 9045 11271
rect 4212 11240 9045 11268
rect 4212 11228 4218 11240
rect 9033 11237 9045 11240
rect 9079 11237 9091 11271
rect 9033 11231 9091 11237
rect 9122 11228 9128 11280
rect 9180 11268 9186 11280
rect 10870 11268 10876 11280
rect 9180 11240 10876 11268
rect 9180 11228 9186 11240
rect 10870 11228 10876 11240
rect 10928 11228 10934 11280
rect 11146 11228 11152 11280
rect 11204 11268 11210 11280
rect 11394 11271 11452 11277
rect 11394 11268 11406 11271
rect 11204 11240 11406 11268
rect 11204 11228 11210 11240
rect 11394 11237 11406 11240
rect 11440 11237 11452 11271
rect 11532 11268 11560 11308
rect 12529 11305 12541 11339
rect 12575 11336 12587 11339
rect 12986 11336 12992 11348
rect 12575 11308 12992 11336
rect 12575 11305 12587 11308
rect 12529 11299 12587 11305
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 13173 11339 13231 11345
rect 13173 11305 13185 11339
rect 13219 11336 13231 11339
rect 13446 11336 13452 11348
rect 13219 11308 13452 11336
rect 13219 11305 13231 11308
rect 13173 11299 13231 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 13817 11339 13875 11345
rect 13817 11305 13829 11339
rect 13863 11336 13875 11339
rect 13906 11336 13912 11348
rect 13863 11308 13912 11336
rect 13863 11305 13875 11308
rect 13817 11299 13875 11305
rect 13906 11296 13912 11308
rect 13964 11296 13970 11348
rect 14829 11339 14887 11345
rect 14829 11336 14841 11339
rect 14384 11308 14841 11336
rect 14185 11271 14243 11277
rect 14185 11268 14197 11271
rect 11532 11240 14197 11268
rect 11394 11231 11452 11237
rect 14185 11237 14197 11240
rect 14231 11237 14243 11271
rect 14185 11231 14243 11237
rect 1854 11160 1860 11212
rect 1912 11200 1918 11212
rect 2409 11203 2467 11209
rect 2409 11200 2421 11203
rect 1912 11172 2421 11200
rect 1912 11160 1918 11172
rect 2409 11169 2421 11172
rect 2455 11169 2467 11203
rect 2409 11163 2467 11169
rect 2501 11203 2559 11209
rect 2501 11169 2513 11203
rect 2547 11200 2559 11203
rect 2866 11200 2872 11212
rect 2547 11172 2872 11200
rect 2547 11169 2559 11172
rect 2501 11163 2559 11169
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 3050 11200 3056 11212
rect 3011 11172 3056 11200
rect 3050 11160 3056 11172
rect 3108 11160 3114 11212
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11200 5227 11203
rect 5534 11200 5540 11212
rect 5215 11172 5540 11200
rect 5215 11169 5227 11172
rect 5169 11163 5227 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 6822 11200 6828 11212
rect 6783 11172 6828 11200
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 7929 11203 7987 11209
rect 7929 11200 7941 11203
rect 7340 11172 7941 11200
rect 7340 11160 7346 11172
rect 7929 11169 7941 11172
rect 7975 11200 7987 11203
rect 8202 11200 8208 11212
rect 7975 11172 8208 11200
rect 7975 11169 7987 11172
rect 7929 11163 7987 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 8941 11203 8999 11209
rect 8941 11169 8953 11203
rect 8987 11200 8999 11203
rect 9674 11200 9680 11212
rect 8987 11172 9680 11200
rect 8987 11169 8999 11172
rect 8941 11163 8999 11169
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 12434 11200 12440 11212
rect 11164 11172 12440 11200
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11132 2743 11135
rect 3234 11132 3240 11144
rect 2731 11104 3240 11132
rect 2731 11101 2743 11104
rect 2685 11095 2743 11101
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11101 5503 11135
rect 5445 11095 5503 11101
rect 2498 11024 2504 11076
rect 2556 11064 2562 11076
rect 2774 11064 2780 11076
rect 2556 11036 2780 11064
rect 2556 11024 2562 11036
rect 2774 11024 2780 11036
rect 2832 11024 2838 11076
rect 4798 11064 4804 11076
rect 4759 11036 4804 11064
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 5460 10996 5488 11095
rect 5626 11092 5632 11144
rect 5684 11132 5690 11144
rect 5810 11132 5816 11144
rect 5684 11104 5816 11132
rect 5684 11092 5690 11104
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 6914 11132 6920 11144
rect 6875 11104 6920 11132
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 7098 11132 7104 11144
rect 7059 11104 7104 11132
rect 7098 11092 7104 11104
rect 7156 11092 7162 11144
rect 7558 11092 7564 11144
rect 7616 11132 7622 11144
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 7616 11104 8033 11132
rect 7616 11092 7622 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11132 9275 11135
rect 9766 11132 9772 11144
rect 9263 11104 9772 11132
rect 9263 11101 9275 11104
rect 9217 11095 9275 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 10134 11132 10140 11144
rect 10095 11104 10140 11132
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 10284 11104 10329 11132
rect 10284 11092 10290 11104
rect 10502 11092 10508 11144
rect 10560 11132 10566 11144
rect 11164 11141 11192 11172
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 12710 11160 12716 11212
rect 12768 11200 12774 11212
rect 14384 11200 14412 11308
rect 14829 11305 14841 11308
rect 14875 11305 14887 11339
rect 14829 11299 14887 11305
rect 15841 11339 15899 11345
rect 15841 11305 15853 11339
rect 15887 11336 15899 11339
rect 16758 11336 16764 11348
rect 15887 11308 16764 11336
rect 15887 11305 15899 11308
rect 15841 11299 15899 11305
rect 14844 11268 14872 11299
rect 16758 11296 16764 11308
rect 16816 11296 16822 11348
rect 16850 11296 16856 11348
rect 16908 11336 16914 11348
rect 18509 11339 18567 11345
rect 18509 11336 18521 11339
rect 16908 11308 18521 11336
rect 16908 11296 16914 11308
rect 18509 11305 18521 11308
rect 18555 11305 18567 11339
rect 19518 11336 19524 11348
rect 19479 11308 19524 11336
rect 18509 11299 18567 11305
rect 19518 11296 19524 11308
rect 19576 11296 19582 11348
rect 20346 11296 20352 11348
rect 20404 11336 20410 11348
rect 20441 11339 20499 11345
rect 20441 11336 20453 11339
rect 20404 11308 20453 11336
rect 20404 11296 20410 11308
rect 20441 11305 20453 11308
rect 20487 11305 20499 11339
rect 20898 11336 20904 11348
rect 20859 11308 20904 11336
rect 20441 11299 20499 11305
rect 20898 11296 20904 11308
rect 20956 11296 20962 11348
rect 14844 11240 15792 11268
rect 15010 11200 15016 11212
rect 12768 11172 14412 11200
rect 14971 11172 15016 11200
rect 12768 11160 12774 11172
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 15764 11209 15792 11240
rect 16298 11228 16304 11280
rect 16356 11268 16362 11280
rect 20622 11268 20628 11280
rect 16356 11240 20628 11268
rect 16356 11228 16362 11240
rect 20622 11228 20628 11240
rect 20680 11228 20686 11280
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11169 15807 11203
rect 16206 11200 16212 11212
rect 16167 11172 16212 11200
rect 15749 11163 15807 11169
rect 16206 11160 16212 11172
rect 16264 11160 16270 11212
rect 17396 11203 17454 11209
rect 17396 11169 17408 11203
rect 17442 11200 17454 11203
rect 17862 11200 17868 11212
rect 17442 11172 17868 11200
rect 17442 11169 17454 11172
rect 17396 11163 17454 11169
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 20254 11200 20260 11212
rect 20215 11172 20260 11200
rect 20254 11160 20260 11172
rect 20312 11160 20318 11212
rect 11149 11135 11207 11141
rect 11149 11132 11161 11135
rect 10560 11104 11161 11132
rect 10560 11092 10566 11104
rect 11149 11101 11161 11104
rect 11195 11101 11207 11135
rect 11149 11095 11207 11101
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 13265 11135 13323 11141
rect 13265 11132 13277 11135
rect 12676 11104 13277 11132
rect 12676 11092 12682 11104
rect 13265 11101 13277 11104
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11132 13507 11135
rect 13722 11132 13728 11144
rect 13495 11104 13728 11132
rect 13495 11101 13507 11104
rect 13449 11095 13507 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 14274 11132 14280 11144
rect 14235 11104 14280 11132
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 14366 11092 14372 11144
rect 14424 11132 14430 11144
rect 14424 11104 14469 11132
rect 14424 11092 14430 11104
rect 15654 11092 15660 11144
rect 15712 11132 15718 11144
rect 16301 11135 16359 11141
rect 16301 11132 16313 11135
rect 15712 11104 16313 11132
rect 15712 11092 15718 11104
rect 16301 11101 16313 11104
rect 16347 11101 16359 11135
rect 16301 11095 16359 11101
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11132 16543 11135
rect 16850 11132 16856 11144
rect 16531 11104 16856 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 16850 11092 16856 11104
rect 16908 11092 16914 11144
rect 17126 11132 17132 11144
rect 17087 11104 17132 11132
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 19426 11092 19432 11144
rect 19484 11132 19490 11144
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 19484 11104 19625 11132
rect 19484 11092 19490 11104
rect 19613 11101 19625 11104
rect 19659 11101 19671 11135
rect 19613 11095 19671 11101
rect 19797 11135 19855 11141
rect 19797 11101 19809 11135
rect 19843 11132 19855 11135
rect 19886 11132 19892 11144
rect 19843 11104 19892 11132
rect 19843 11101 19855 11104
rect 19797 11095 19855 11101
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 7374 11024 7380 11076
rect 7432 11064 7438 11076
rect 7469 11067 7527 11073
rect 7469 11064 7481 11067
rect 7432 11036 7481 11064
rect 7432 11024 7438 11036
rect 7469 11033 7481 11036
rect 7515 11033 7527 11067
rect 7469 11027 7527 11033
rect 8202 11024 8208 11076
rect 8260 11064 8266 11076
rect 9677 11067 9735 11073
rect 8260 11036 9628 11064
rect 8260 11024 8266 11036
rect 5626 10996 5632 11008
rect 5460 10968 5632 10996
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 9490 10996 9496 11008
rect 6788 10968 9496 10996
rect 6788 10956 6794 10968
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 9600 10996 9628 11036
rect 9677 11033 9689 11067
rect 9723 11064 9735 11067
rect 11054 11064 11060 11076
rect 9723 11036 11060 11064
rect 9723 11033 9735 11036
rect 9677 11027 9735 11033
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 12805 11067 12863 11073
rect 12805 11033 12817 11067
rect 12851 11064 12863 11067
rect 14182 11064 14188 11076
rect 12851 11036 14188 11064
rect 12851 11033 12863 11036
rect 12805 11027 12863 11033
rect 14182 11024 14188 11036
rect 14240 11024 14246 11076
rect 15562 11024 15568 11076
rect 15620 11064 15626 11076
rect 16574 11064 16580 11076
rect 15620 11036 16580 11064
rect 15620 11024 15626 11036
rect 16574 11024 16580 11036
rect 16632 11064 16638 11076
rect 17144 11064 17172 11092
rect 16632 11036 17172 11064
rect 16632 11024 16638 11036
rect 18138 11024 18144 11076
rect 18196 11064 18202 11076
rect 18874 11064 18880 11076
rect 18196 11036 18880 11064
rect 18196 11024 18202 11036
rect 18874 11024 18880 11036
rect 18932 11024 18938 11076
rect 19058 11024 19064 11076
rect 19116 11064 19122 11076
rect 19153 11067 19211 11073
rect 19153 11064 19165 11067
rect 19116 11036 19165 11064
rect 19116 11024 19122 11036
rect 19153 11033 19165 11036
rect 19199 11033 19211 11067
rect 19153 11027 19211 11033
rect 10410 10996 10416 11008
rect 9600 10968 10416 10996
rect 10410 10956 10416 10968
rect 10468 10956 10474 11008
rect 16482 10956 16488 11008
rect 16540 10996 16546 11008
rect 18598 10996 18604 11008
rect 16540 10968 18604 10996
rect 16540 10956 16546 10968
rect 18598 10956 18604 10968
rect 18656 10956 18662 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 3234 10792 3240 10804
rect 3195 10764 3240 10792
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 7156 10764 8217 10792
rect 7156 10752 7162 10764
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 10226 10792 10232 10804
rect 10187 10764 10232 10792
rect 8205 10755 8263 10761
rect 10226 10752 10232 10764
rect 10284 10752 10290 10804
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 10468 10764 11560 10792
rect 10468 10752 10474 10764
rect 5813 10727 5871 10733
rect 5813 10693 5825 10727
rect 5859 10724 5871 10727
rect 5994 10724 6000 10736
rect 5859 10696 6000 10724
rect 5859 10693 5871 10696
rect 5813 10687 5871 10693
rect 5994 10684 6000 10696
rect 6052 10684 6058 10736
rect 3510 10656 3516 10668
rect 3471 10628 3516 10656
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 6638 10616 6644 10668
rect 6696 10656 6702 10668
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6696 10628 6837 10656
rect 6696 10616 6702 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 8846 10656 8852 10668
rect 8807 10628 8852 10656
rect 6825 10619 6883 10625
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 10244 10656 10272 10752
rect 11532 10656 11560 10764
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 14093 10795 14151 10801
rect 11664 10764 14044 10792
rect 11664 10752 11670 10764
rect 14016 10724 14044 10764
rect 14093 10761 14105 10795
rect 14139 10792 14151 10795
rect 14274 10792 14280 10804
rect 14139 10764 14280 10792
rect 14139 10761 14151 10764
rect 14093 10755 14151 10761
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 15105 10795 15163 10801
rect 15105 10761 15117 10795
rect 15151 10792 15163 10795
rect 16206 10792 16212 10804
rect 15151 10764 16212 10792
rect 15151 10761 15163 10764
rect 15105 10755 15163 10761
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 16298 10752 16304 10804
rect 16356 10792 16362 10804
rect 19794 10792 19800 10804
rect 16356 10764 19800 10792
rect 16356 10752 16362 10764
rect 19794 10752 19800 10764
rect 19852 10752 19858 10804
rect 14016 10696 17264 10724
rect 10244 10628 10640 10656
rect 11532 10628 12572 10656
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 1857 10591 1915 10597
rect 1857 10588 1869 10591
rect 1728 10560 1869 10588
rect 1728 10548 1734 10560
rect 1857 10557 1869 10560
rect 1903 10588 1915 10591
rect 3142 10588 3148 10600
rect 1903 10560 3148 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 3142 10548 3148 10560
rect 3200 10588 3206 10600
rect 4154 10588 4160 10600
rect 3200 10560 4160 10588
rect 3200 10548 3206 10560
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 4424 10591 4482 10597
rect 4424 10557 4436 10591
rect 4470 10588 4482 10591
rect 5442 10588 5448 10600
rect 4470 10560 5448 10588
rect 4470 10557 4482 10560
rect 4424 10551 4482 10557
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 5997 10591 6055 10597
rect 5997 10557 6009 10591
rect 6043 10588 6055 10591
rect 7650 10588 7656 10600
rect 6043 10560 7656 10588
rect 6043 10557 6055 10560
rect 5997 10551 6055 10557
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 8478 10548 8484 10600
rect 8536 10588 8542 10600
rect 10321 10591 10379 10597
rect 10321 10588 10333 10591
rect 8536 10560 10333 10588
rect 8536 10548 8542 10560
rect 10321 10557 10333 10560
rect 10367 10557 10379 10591
rect 10502 10588 10508 10600
rect 10463 10560 10508 10588
rect 10321 10551 10379 10557
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 10612 10588 10640 10628
rect 10761 10591 10819 10597
rect 10761 10588 10773 10591
rect 10612 10560 10773 10588
rect 10761 10557 10773 10560
rect 10807 10557 10819 10591
rect 12434 10588 12440 10600
rect 12395 10560 12440 10588
rect 10761 10551 10819 10557
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 2124 10523 2182 10529
rect 2124 10489 2136 10523
rect 2170 10520 2182 10523
rect 2498 10520 2504 10532
rect 2170 10492 2504 10520
rect 2170 10489 2182 10492
rect 2124 10483 2182 10489
rect 2498 10480 2504 10492
rect 2556 10480 2562 10532
rect 3970 10480 3976 10532
rect 4028 10520 4034 10532
rect 7092 10523 7150 10529
rect 4028 10492 5764 10520
rect 4028 10480 4034 10492
rect 1946 10412 1952 10464
rect 2004 10452 2010 10464
rect 3234 10452 3240 10464
rect 2004 10424 3240 10452
rect 2004 10412 2010 10424
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 5537 10455 5595 10461
rect 5537 10421 5549 10455
rect 5583 10452 5595 10455
rect 5626 10452 5632 10464
rect 5583 10424 5632 10452
rect 5583 10421 5595 10424
rect 5537 10415 5595 10421
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 5736 10452 5764 10492
rect 7092 10489 7104 10523
rect 7138 10520 7150 10523
rect 7466 10520 7472 10532
rect 7138 10492 7472 10520
rect 7138 10489 7150 10492
rect 7092 10483 7150 10489
rect 7466 10480 7472 10492
rect 7524 10480 7530 10532
rect 9116 10523 9174 10529
rect 9116 10489 9128 10523
rect 9162 10520 9174 10523
rect 9766 10520 9772 10532
rect 9162 10492 9772 10520
rect 9162 10489 9174 10492
rect 9116 10483 9174 10489
rect 9766 10480 9772 10492
rect 9824 10480 9830 10532
rect 12544 10520 12572 10628
rect 14458 10616 14464 10668
rect 14516 10656 14522 10668
rect 14645 10659 14703 10665
rect 14645 10656 14657 10659
rect 14516 10628 14657 10656
rect 14516 10616 14522 10628
rect 14645 10625 14657 10628
rect 14691 10656 14703 10659
rect 15102 10656 15108 10668
rect 14691 10628 15108 10656
rect 14691 10625 14703 10628
rect 14645 10619 14703 10625
rect 15102 10616 15108 10628
rect 15160 10616 15166 10668
rect 15562 10656 15568 10668
rect 15523 10628 15568 10656
rect 15562 10616 15568 10628
rect 15620 10616 15626 10668
rect 15746 10656 15752 10668
rect 15707 10628 15752 10656
rect 15746 10616 15752 10628
rect 15804 10616 15810 10668
rect 16482 10616 16488 10668
rect 16540 10656 16546 10668
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 16540 10628 16681 10656
rect 16540 10616 16546 10628
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 12710 10597 12716 10600
rect 12704 10588 12716 10597
rect 12623 10560 12716 10588
rect 12704 10551 12716 10560
rect 12768 10588 12774 10600
rect 12986 10588 12992 10600
rect 12768 10560 12992 10588
rect 12710 10548 12716 10551
rect 12768 10548 12774 10560
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 17037 10591 17095 10597
rect 17037 10588 17049 10591
rect 13096 10560 17049 10588
rect 13096 10520 13124 10560
rect 17037 10557 17049 10560
rect 17083 10557 17095 10591
rect 17037 10551 17095 10557
rect 14461 10523 14519 10529
rect 14461 10520 14473 10523
rect 10971 10492 12020 10520
rect 12544 10492 13124 10520
rect 13188 10492 14473 10520
rect 10226 10452 10232 10464
rect 5736 10424 10232 10452
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 10321 10455 10379 10461
rect 10321 10421 10333 10455
rect 10367 10452 10379 10455
rect 10971 10452 10999 10492
rect 10367 10424 10999 10452
rect 10367 10421 10379 10424
rect 10321 10415 10379 10421
rect 11238 10412 11244 10464
rect 11296 10452 11302 10464
rect 11885 10455 11943 10461
rect 11885 10452 11897 10455
rect 11296 10424 11897 10452
rect 11296 10412 11302 10424
rect 11885 10421 11897 10424
rect 11931 10421 11943 10455
rect 11992 10452 12020 10492
rect 13188 10452 13216 10492
rect 14461 10489 14473 10492
rect 14507 10489 14519 10523
rect 14461 10483 14519 10489
rect 15473 10523 15531 10529
rect 15473 10489 15485 10523
rect 15519 10520 15531 10523
rect 16485 10523 16543 10529
rect 15519 10492 16160 10520
rect 15519 10489 15531 10492
rect 15473 10483 15531 10489
rect 11992 10424 13216 10452
rect 11885 10415 11943 10421
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13780 10424 13829 10452
rect 13780 10412 13786 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 13817 10415 13875 10421
rect 14553 10455 14611 10461
rect 14553 10421 14565 10455
rect 14599 10452 14611 10455
rect 16022 10452 16028 10464
rect 14599 10424 16028 10452
rect 14599 10421 14611 10424
rect 14553 10415 14611 10421
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 16132 10461 16160 10492
rect 16485 10489 16497 10523
rect 16531 10520 16543 10523
rect 17129 10523 17187 10529
rect 17129 10520 17141 10523
rect 16531 10492 17141 10520
rect 16531 10489 16543 10492
rect 16485 10483 16543 10489
rect 17129 10489 17141 10492
rect 17175 10489 17187 10523
rect 17236 10520 17264 10696
rect 19794 10616 19800 10668
rect 19852 10656 19858 10668
rect 19978 10656 19984 10668
rect 19852 10628 19984 10656
rect 19852 10616 19858 10628
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 20622 10656 20628 10668
rect 20583 10628 20628 10656
rect 20622 10616 20628 10628
rect 20680 10616 20686 10668
rect 20717 10659 20775 10665
rect 20717 10625 20729 10659
rect 20763 10625 20775 10659
rect 20717 10619 20775 10625
rect 18417 10591 18475 10597
rect 18417 10557 18429 10591
rect 18463 10588 18475 10591
rect 18506 10588 18512 10600
rect 18463 10560 18512 10588
rect 18463 10557 18475 10560
rect 18417 10551 18475 10557
rect 18506 10548 18512 10560
rect 18564 10548 18570 10600
rect 18776 10591 18834 10597
rect 18776 10557 18788 10591
rect 18822 10588 18834 10591
rect 19518 10588 19524 10600
rect 18822 10560 19524 10588
rect 18822 10557 18834 10560
rect 18776 10551 18834 10557
rect 19518 10548 19524 10560
rect 19576 10588 19582 10600
rect 20438 10588 20444 10600
rect 19576 10560 20444 10588
rect 19576 10548 19582 10560
rect 20438 10548 20444 10560
rect 20496 10548 20502 10600
rect 20530 10548 20536 10600
rect 20588 10588 20594 10600
rect 20732 10588 20760 10619
rect 20588 10560 20760 10588
rect 20588 10548 20594 10560
rect 17236 10492 20576 10520
rect 17129 10483 17187 10489
rect 16117 10455 16175 10461
rect 16117 10421 16129 10455
rect 16163 10421 16175 10455
rect 16574 10452 16580 10464
rect 16535 10424 16580 10452
rect 16117 10415 16175 10421
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 17037 10455 17095 10461
rect 17037 10421 17049 10455
rect 17083 10452 17095 10455
rect 18322 10452 18328 10464
rect 17083 10424 18328 10452
rect 17083 10421 17095 10424
rect 17037 10415 17095 10421
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 18417 10455 18475 10461
rect 18417 10421 18429 10455
rect 18463 10452 18475 10455
rect 19150 10452 19156 10464
rect 18463 10424 19156 10452
rect 18463 10421 18475 10424
rect 18417 10415 18475 10421
rect 19150 10412 19156 10424
rect 19208 10452 19214 10464
rect 19702 10452 19708 10464
rect 19208 10424 19708 10452
rect 19208 10412 19214 10424
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 19886 10452 19892 10464
rect 19847 10424 19892 10452
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 20162 10452 20168 10464
rect 20123 10424 20168 10452
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 20548 10461 20576 10492
rect 20533 10455 20591 10461
rect 20533 10421 20545 10455
rect 20579 10421 20591 10455
rect 20533 10415 20591 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 2498 10208 2504 10260
rect 2556 10248 2562 10260
rect 3053 10251 3111 10257
rect 3053 10248 3065 10251
rect 2556 10220 3065 10248
rect 2556 10208 2562 10220
rect 3053 10217 3065 10220
rect 3099 10217 3111 10251
rect 3053 10211 3111 10217
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 7377 10251 7435 10257
rect 4120 10220 5764 10248
rect 4120 10208 4126 10220
rect 4608 10183 4666 10189
rect 4608 10149 4620 10183
rect 4654 10180 4666 10183
rect 5626 10180 5632 10192
rect 4654 10152 5632 10180
rect 4654 10149 4666 10152
rect 4608 10143 4666 10149
rect 5626 10140 5632 10152
rect 5684 10140 5690 10192
rect 5736 10180 5764 10220
rect 7377 10217 7389 10251
rect 7423 10248 7435 10251
rect 7558 10248 7564 10260
rect 7423 10220 7564 10248
rect 7423 10217 7435 10220
rect 7377 10211 7435 10217
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 7650 10208 7656 10260
rect 7708 10248 7714 10260
rect 8938 10248 8944 10260
rect 7708 10220 8944 10248
rect 7708 10208 7714 10220
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9674 10248 9680 10260
rect 9635 10220 9680 10248
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 10597 10251 10655 10257
rect 10597 10217 10609 10251
rect 10643 10248 10655 10251
rect 12069 10251 12127 10257
rect 12069 10248 12081 10251
rect 10643 10220 12081 10248
rect 10643 10217 10655 10220
rect 10597 10211 10655 10217
rect 12069 10217 12081 10220
rect 12115 10217 12127 10251
rect 16850 10248 16856 10260
rect 16811 10220 16856 10248
rect 12069 10211 12127 10217
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 5736 10152 10640 10180
rect 1940 10115 1998 10121
rect 1940 10081 1952 10115
rect 1986 10112 1998 10115
rect 2222 10112 2228 10124
rect 1986 10084 2228 10112
rect 1986 10081 1998 10084
rect 1940 10075 1998 10081
rect 2222 10072 2228 10084
rect 2280 10072 2286 10124
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 4341 10115 4399 10121
rect 4341 10112 4353 10115
rect 4212 10084 4353 10112
rect 4212 10072 4218 10084
rect 4341 10081 4353 10084
rect 4387 10112 4399 10115
rect 5074 10112 5080 10124
rect 4387 10084 5080 10112
rect 4387 10081 4399 10084
rect 4341 10075 4399 10081
rect 5074 10072 5080 10084
rect 5132 10112 5138 10124
rect 5132 10084 5396 10112
rect 5132 10072 5138 10084
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 5368 10044 5396 10084
rect 5718 10072 5724 10124
rect 5776 10112 5782 10124
rect 6253 10115 6311 10121
rect 6253 10112 6265 10115
rect 5776 10084 6265 10112
rect 5776 10072 5782 10084
rect 6253 10081 6265 10084
rect 6299 10081 6311 10115
rect 6253 10075 6311 10081
rect 7742 10072 7748 10124
rect 7800 10112 7806 10124
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 7800 10084 7849 10112
rect 7800 10072 7806 10084
rect 7837 10081 7849 10084
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 8196 10115 8254 10121
rect 8196 10081 8208 10115
rect 8242 10112 8254 10115
rect 9490 10112 9496 10124
rect 8242 10084 9496 10112
rect 8242 10081 8254 10084
rect 8196 10075 8254 10081
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 9950 10112 9956 10124
rect 9732 10084 9956 10112
rect 9732 10072 9738 10084
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 5994 10044 6000 10056
rect 5368 10016 6000 10044
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 7926 10044 7932 10056
rect 7887 10016 7932 10044
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 9950 9976 9956 9988
rect 5276 9948 5856 9976
rect 3602 9868 3608 9920
rect 3660 9908 3666 9920
rect 4062 9908 4068 9920
rect 3660 9880 4068 9908
rect 3660 9868 3666 9880
rect 4062 9868 4068 9880
rect 4120 9908 4126 9920
rect 5276 9908 5304 9948
rect 5718 9908 5724 9920
rect 4120 9880 5304 9908
rect 5679 9880 5724 9908
rect 4120 9868 4126 9880
rect 5718 9868 5724 9880
rect 5776 9868 5782 9920
rect 5828 9908 5856 9948
rect 8864 9948 9956 9976
rect 8864 9908 8892 9948
rect 9950 9936 9956 9948
rect 10008 9936 10014 9988
rect 5828 9880 8892 9908
rect 9309 9911 9367 9917
rect 9309 9877 9321 9911
rect 9355 9908 9367 9911
rect 9766 9908 9772 9920
rect 9355 9880 9772 9908
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 9766 9868 9772 9880
rect 9824 9908 9830 9920
rect 10226 9908 10232 9920
rect 9824 9880 10232 9908
rect 9824 9868 9830 9880
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 10612 9908 10640 10152
rect 10686 10140 10692 10192
rect 10744 10180 10750 10192
rect 11057 10183 11115 10189
rect 11057 10180 11069 10183
rect 10744 10152 11069 10180
rect 10744 10140 10750 10152
rect 11057 10149 11069 10152
rect 11103 10149 11115 10183
rect 12710 10180 12716 10192
rect 11057 10143 11115 10149
rect 12360 10152 12716 10180
rect 10965 10115 11023 10121
rect 10965 10081 10977 10115
rect 11011 10112 11023 10115
rect 11146 10112 11152 10124
rect 11011 10084 11152 10112
rect 11011 10081 11023 10084
rect 10965 10075 11023 10081
rect 11146 10072 11152 10084
rect 11204 10112 11210 10124
rect 11606 10112 11612 10124
rect 11204 10084 11612 10112
rect 11204 10072 11210 10084
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 11974 10112 11980 10124
rect 11935 10084 11980 10112
rect 11974 10072 11980 10084
rect 12032 10072 12038 10124
rect 12360 10112 12388 10152
rect 12710 10140 12716 10152
rect 12768 10140 12774 10192
rect 12888 10183 12946 10189
rect 12888 10149 12900 10183
rect 12934 10180 12946 10183
rect 13722 10180 13728 10192
rect 12934 10152 13728 10180
rect 12934 10149 12946 10152
rect 12888 10143 12946 10149
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 13814 10140 13820 10192
rect 13872 10180 13878 10192
rect 16298 10180 16304 10192
rect 13872 10152 16304 10180
rect 13872 10140 13878 10152
rect 16298 10140 16304 10152
rect 16356 10140 16362 10192
rect 16868 10180 16896 10208
rect 17374 10183 17432 10189
rect 17374 10180 17386 10183
rect 16868 10152 17386 10180
rect 17374 10149 17386 10152
rect 17420 10149 17432 10183
rect 17374 10143 17432 10149
rect 19420 10183 19478 10189
rect 19420 10149 19432 10183
rect 19466 10180 19478 10183
rect 19886 10180 19892 10192
rect 19466 10152 19892 10180
rect 19466 10149 19478 10152
rect 19420 10143 19478 10149
rect 19886 10140 19892 10152
rect 19944 10140 19950 10192
rect 12268 10084 12388 10112
rect 11238 10044 11244 10056
rect 11199 10016 11244 10044
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 12268 10053 12296 10084
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 12621 10115 12679 10121
rect 12621 10112 12633 10115
rect 12492 10084 12633 10112
rect 12492 10072 12498 10084
rect 12621 10081 12633 10084
rect 12667 10112 12679 10115
rect 13998 10112 14004 10124
rect 12667 10084 14004 10112
rect 12667 10081 12679 10084
rect 12621 10075 12679 10081
rect 13998 10072 14004 10084
rect 14056 10072 14062 10124
rect 14182 10072 14188 10124
rect 14240 10112 14246 10124
rect 14277 10115 14335 10121
rect 14277 10112 14289 10115
rect 14240 10084 14289 10112
rect 14240 10072 14246 10084
rect 14277 10081 14289 10084
rect 14323 10081 14335 10115
rect 14277 10075 14335 10081
rect 15378 10072 15384 10124
rect 15436 10112 15442 10124
rect 15746 10121 15752 10124
rect 15729 10115 15752 10121
rect 15729 10112 15741 10115
rect 15436 10084 15741 10112
rect 15436 10072 15442 10084
rect 15729 10081 15741 10084
rect 15804 10112 15810 10124
rect 15804 10084 15877 10112
rect 15729 10075 15752 10081
rect 15746 10072 15752 10075
rect 15804 10072 15810 10084
rect 16022 10072 16028 10124
rect 16080 10112 16086 10124
rect 16758 10112 16764 10124
rect 16080 10084 16764 10112
rect 16080 10072 16086 10084
rect 16758 10072 16764 10084
rect 16816 10072 16822 10124
rect 17126 10112 17132 10124
rect 17039 10084 17132 10112
rect 17126 10072 17132 10084
rect 17184 10112 17190 10124
rect 17184 10084 19196 10112
rect 17184 10072 17190 10084
rect 19168 10056 19196 10084
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 14553 10047 14611 10053
rect 14553 10013 14565 10047
rect 14599 10044 14611 10047
rect 15102 10044 15108 10056
rect 14599 10016 15108 10044
rect 14599 10013 14611 10016
rect 14553 10007 14611 10013
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 15470 10044 15476 10056
rect 15431 10016 15476 10044
rect 15470 10004 15476 10016
rect 15528 10004 15534 10056
rect 19150 10044 19156 10056
rect 19111 10016 19156 10044
rect 19150 10004 19156 10016
rect 19208 10004 19214 10056
rect 11609 9979 11667 9985
rect 11609 9945 11621 9979
rect 11655 9976 11667 9979
rect 12618 9976 12624 9988
rect 11655 9948 12624 9976
rect 11655 9945 11667 9948
rect 11609 9939 11667 9945
rect 12618 9936 12624 9948
rect 12676 9936 12682 9988
rect 12894 9908 12900 9920
rect 10612 9880 12900 9908
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 13354 9868 13360 9920
rect 13412 9908 13418 9920
rect 14001 9911 14059 9917
rect 14001 9908 14013 9911
rect 13412 9880 14013 9908
rect 13412 9868 13418 9880
rect 14001 9877 14013 9880
rect 14047 9877 14059 9911
rect 14001 9871 14059 9877
rect 18509 9911 18567 9917
rect 18509 9877 18521 9911
rect 18555 9908 18567 9911
rect 18598 9908 18604 9920
rect 18555 9880 18604 9908
rect 18555 9877 18567 9880
rect 18509 9871 18567 9877
rect 18598 9868 18604 9880
rect 18656 9868 18662 9920
rect 20530 9908 20536 9920
rect 20491 9880 20536 9908
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 5552 9676 6132 9704
rect 1854 9636 1860 9648
rect 1815 9608 1860 9636
rect 1854 9596 1860 9608
rect 1912 9596 1918 9648
rect 2866 9636 2872 9648
rect 2827 9608 2872 9636
rect 2866 9596 2872 9608
rect 2924 9596 2930 9648
rect 4246 9596 4252 9648
rect 4304 9636 4310 9648
rect 4433 9639 4491 9645
rect 4433 9636 4445 9639
rect 4304 9608 4445 9636
rect 4304 9596 4310 9608
rect 4433 9605 4445 9608
rect 4479 9605 4491 9639
rect 5552 9636 5580 9676
rect 4433 9599 4491 9605
rect 4540 9608 5580 9636
rect 2498 9568 2504 9580
rect 2459 9540 2504 9568
rect 2498 9528 2504 9540
rect 2556 9568 2562 9580
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 2556 9540 3433 9568
rect 2556 9528 2562 9540
rect 3421 9537 3433 9540
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 3878 9528 3884 9580
rect 3936 9568 3942 9580
rect 4540 9568 4568 9608
rect 5626 9596 5632 9648
rect 5684 9636 5690 9648
rect 5684 9608 6040 9636
rect 5684 9596 5690 9608
rect 3936 9540 4568 9568
rect 3936 9528 3942 9540
rect 4798 9528 4804 9580
rect 4856 9568 4862 9580
rect 4893 9571 4951 9577
rect 4893 9568 4905 9571
rect 4856 9540 4905 9568
rect 4856 9528 4862 9540
rect 4893 9537 4905 9540
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9568 5135 9571
rect 5718 9568 5724 9580
rect 5123 9540 5724 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 6012 9577 6040 9608
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 3510 9460 3516 9512
rect 3568 9500 3574 9512
rect 3786 9500 3792 9512
rect 3568 9472 3792 9500
rect 3568 9460 3574 9472
rect 3786 9460 3792 9472
rect 3844 9500 3850 9512
rect 5166 9500 5172 9512
rect 3844 9472 5172 9500
rect 3844 9460 3850 9472
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 5350 9460 5356 9512
rect 5408 9500 5414 9512
rect 5905 9503 5963 9509
rect 5905 9500 5917 9503
rect 5408 9472 5917 9500
rect 5408 9460 5414 9472
rect 5905 9469 5917 9472
rect 5951 9469 5963 9503
rect 6104 9500 6132 9676
rect 7926 9664 7932 9716
rect 7984 9704 7990 9716
rect 8662 9704 8668 9716
rect 7984 9676 8668 9704
rect 7984 9664 7990 9676
rect 8662 9664 8668 9676
rect 8720 9664 8726 9716
rect 8754 9664 8760 9716
rect 8812 9664 8818 9716
rect 9490 9664 9496 9716
rect 9548 9704 9554 9716
rect 9548 9676 9720 9704
rect 9548 9664 9554 9676
rect 6914 9636 6920 9648
rect 6875 9608 6920 9636
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 8772 9636 8800 9664
rect 7208 9608 8800 9636
rect 9692 9636 9720 9676
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 13814 9704 13820 9716
rect 10008 9676 13820 9704
rect 10008 9664 10014 9676
rect 13814 9664 13820 9676
rect 13872 9664 13878 9716
rect 15378 9704 15384 9716
rect 14016 9676 14964 9704
rect 15339 9676 15384 9704
rect 10137 9639 10195 9645
rect 10137 9636 10149 9639
rect 9692 9608 10149 9636
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 7208 9568 7236 9608
rect 10137 9605 10149 9608
rect 10183 9636 10195 9639
rect 10183 9608 11008 9636
rect 10183 9605 10195 9608
rect 10137 9599 10195 9605
rect 7374 9568 7380 9580
rect 6871 9540 7236 9568
rect 7335 9540 7380 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 7466 9528 7472 9580
rect 7524 9568 7530 9580
rect 7524 9540 7569 9568
rect 7524 9528 7530 9540
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 8570 9568 8576 9580
rect 7892 9540 8576 9568
rect 7892 9528 7898 9540
rect 8570 9528 8576 9540
rect 8628 9528 8634 9580
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 10980 9577 11008 9608
rect 11054 9596 11060 9648
rect 11112 9636 11118 9648
rect 11333 9639 11391 9645
rect 11333 9636 11345 9639
rect 11112 9608 11345 9636
rect 11112 9596 11118 9608
rect 11333 9605 11345 9608
rect 11379 9605 11391 9639
rect 11333 9599 11391 9605
rect 12805 9639 12863 9645
rect 12805 9605 12817 9639
rect 12851 9636 12863 9639
rect 13262 9636 13268 9648
rect 12851 9608 13268 9636
rect 12851 9605 12863 9608
rect 12805 9599 12863 9605
rect 13262 9596 13268 9608
rect 13320 9596 13326 9648
rect 13722 9636 13728 9648
rect 13372 9608 13728 9636
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 8720 9540 8769 9568
rect 8720 9528 8726 9540
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 10965 9571 11023 9577
rect 10965 9537 10977 9571
rect 11011 9537 11023 9571
rect 13372 9568 13400 9608
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 13906 9596 13912 9648
rect 13964 9636 13970 9648
rect 14016 9636 14044 9676
rect 13964 9608 14044 9636
rect 14936 9636 14964 9676
rect 15378 9664 15384 9676
rect 15436 9704 15442 9716
rect 15436 9676 16252 9704
rect 15436 9664 15442 9676
rect 15654 9636 15660 9648
rect 14936 9608 15056 9636
rect 15615 9608 15660 9636
rect 13964 9596 13970 9608
rect 10965 9531 11023 9537
rect 11072 9540 13400 9568
rect 13449 9571 13507 9577
rect 10594 9500 10600 9512
rect 6104 9472 10600 9500
rect 5905 9463 5963 9469
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 10781 9503 10839 9509
rect 10781 9500 10793 9503
rect 10744 9472 10793 9500
rect 10744 9460 10750 9472
rect 10781 9469 10793 9472
rect 10827 9500 10839 9503
rect 11072 9500 11100 9540
rect 13449 9537 13461 9571
rect 13495 9568 13507 9571
rect 13814 9568 13820 9580
rect 13495 9540 13820 9568
rect 13495 9537 13507 9540
rect 13449 9531 13507 9537
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 13998 9568 14004 9580
rect 13959 9540 14004 9568
rect 13998 9528 14004 9540
rect 14056 9528 14062 9580
rect 15028 9568 15056 9608
rect 15654 9596 15660 9608
rect 15712 9596 15718 9648
rect 16224 9577 16252 9676
rect 16298 9664 16304 9716
rect 16356 9704 16362 9716
rect 17954 9704 17960 9716
rect 16356 9676 17960 9704
rect 16356 9664 16362 9676
rect 17954 9664 17960 9676
rect 18012 9664 18018 9716
rect 18509 9639 18567 9645
rect 18509 9605 18521 9639
rect 18555 9605 18567 9639
rect 19426 9636 19432 9648
rect 18509 9599 18567 9605
rect 18984 9608 19432 9636
rect 16209 9571 16267 9577
rect 15028 9540 16160 9568
rect 10827 9472 11100 9500
rect 11333 9503 11391 9509
rect 10827 9469 10839 9472
rect 10781 9463 10839 9469
rect 11333 9469 11345 9503
rect 11379 9500 11391 9503
rect 11425 9503 11483 9509
rect 11425 9500 11437 9503
rect 11379 9472 11437 9500
rect 11379 9469 11391 9472
rect 11333 9463 11391 9469
rect 11425 9469 11437 9472
rect 11471 9469 11483 9503
rect 16025 9503 16083 9509
rect 16025 9500 16037 9503
rect 11425 9463 11483 9469
rect 11532 9472 16037 9500
rect 3237 9435 3295 9441
rect 3237 9401 3249 9435
rect 3283 9432 3295 9435
rect 4706 9432 4712 9444
rect 3283 9404 4712 9432
rect 3283 9401 3295 9404
rect 3237 9395 3295 9401
rect 4706 9392 4712 9404
rect 4764 9392 4770 9444
rect 4801 9435 4859 9441
rect 4801 9401 4813 9435
rect 4847 9432 4859 9435
rect 4847 9404 5488 9432
rect 4847 9401 4859 9404
rect 4801 9395 4859 9401
rect 1394 9364 1400 9376
rect 1355 9336 1400 9364
rect 1394 9324 1400 9336
rect 1452 9324 1458 9376
rect 1946 9324 1952 9376
rect 2004 9364 2010 9376
rect 2225 9367 2283 9373
rect 2225 9364 2237 9367
rect 2004 9336 2237 9364
rect 2004 9324 2010 9336
rect 2225 9333 2237 9336
rect 2271 9333 2283 9367
rect 2225 9327 2283 9333
rect 2317 9367 2375 9373
rect 2317 9333 2329 9367
rect 2363 9364 2375 9367
rect 2774 9364 2780 9376
rect 2363 9336 2780 9364
rect 2363 9333 2375 9336
rect 2317 9327 2375 9333
rect 2774 9324 2780 9336
rect 2832 9324 2838 9376
rect 3329 9367 3387 9373
rect 3329 9333 3341 9367
rect 3375 9364 3387 9367
rect 4062 9364 4068 9376
rect 3375 9336 4068 9364
rect 3375 9333 3387 9336
rect 3329 9327 3387 9333
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 5460 9373 5488 9404
rect 6178 9392 6184 9444
rect 6236 9432 6242 9444
rect 8294 9432 8300 9444
rect 6236 9404 8300 9432
rect 6236 9392 6242 9404
rect 8294 9392 8300 9404
rect 8352 9392 8358 9444
rect 9024 9435 9082 9441
rect 9024 9401 9036 9435
rect 9070 9432 9082 9435
rect 9306 9432 9312 9444
rect 9070 9404 9312 9432
rect 9070 9401 9082 9404
rect 9024 9395 9082 9401
rect 9306 9392 9312 9404
rect 9364 9392 9370 9444
rect 9398 9392 9404 9444
rect 9456 9432 9462 9444
rect 11532 9432 11560 9472
rect 16025 9469 16037 9472
rect 16071 9469 16083 9503
rect 16132 9500 16160 9540
rect 16209 9537 16221 9571
rect 16255 9537 16267 9571
rect 16209 9531 16267 9537
rect 16482 9528 16488 9580
rect 16540 9568 16546 9580
rect 17221 9571 17279 9577
rect 17221 9568 17233 9571
rect 16540 9540 17233 9568
rect 16540 9528 16546 9540
rect 17221 9537 17233 9540
rect 17267 9537 17279 9571
rect 18524 9568 18552 9599
rect 18984 9568 19012 9608
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 19518 9596 19524 9648
rect 19576 9596 19582 9648
rect 18524 9540 19012 9568
rect 19107 9571 19165 9577
rect 17221 9531 17279 9537
rect 19107 9537 19119 9571
rect 19153 9568 19165 9571
rect 19536 9568 19564 9596
rect 19153 9540 19564 9568
rect 19153 9537 19165 9540
rect 19107 9531 19165 9537
rect 17954 9500 17960 9512
rect 16132 9472 17960 9500
rect 16025 9463 16083 9469
rect 17954 9460 17960 9472
rect 18012 9460 18018 9512
rect 18969 9503 19027 9509
rect 18969 9469 18981 9503
rect 19015 9500 19027 9503
rect 19334 9500 19340 9512
rect 19015 9472 19340 9500
rect 19015 9469 19027 9472
rect 18969 9463 19027 9469
rect 19334 9460 19340 9472
rect 19392 9460 19398 9512
rect 19521 9503 19579 9509
rect 19521 9469 19533 9503
rect 19567 9469 19579 9503
rect 19521 9463 19579 9469
rect 19788 9503 19846 9509
rect 19788 9469 19800 9503
rect 19834 9500 19846 9503
rect 20530 9500 20536 9512
rect 19834 9472 20536 9500
rect 19834 9469 19846 9472
rect 19788 9463 19846 9469
rect 9456 9404 11560 9432
rect 11701 9435 11759 9441
rect 9456 9392 9462 9404
rect 11701 9401 11713 9435
rect 11747 9432 11759 9435
rect 12894 9432 12900 9444
rect 11747 9404 12900 9432
rect 11747 9401 11759 9404
rect 11701 9395 11759 9401
rect 12894 9392 12900 9404
rect 12952 9392 12958 9444
rect 13170 9432 13176 9444
rect 13131 9404 13176 9432
rect 13170 9392 13176 9404
rect 13228 9392 13234 9444
rect 13998 9392 14004 9444
rect 14056 9432 14062 9444
rect 14246 9435 14304 9441
rect 14246 9432 14258 9435
rect 14056 9404 14258 9432
rect 14056 9392 14062 9404
rect 14246 9401 14258 9404
rect 14292 9401 14304 9435
rect 18877 9435 18935 9441
rect 18877 9432 18889 9435
rect 14246 9395 14304 9401
rect 14384 9404 18889 9432
rect 5445 9367 5503 9373
rect 5445 9333 5457 9367
rect 5491 9333 5503 9367
rect 5810 9364 5816 9376
rect 5771 9336 5816 9364
rect 5445 9327 5503 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 6825 9367 6883 9373
rect 6825 9364 6837 9367
rect 5960 9336 6837 9364
rect 5960 9324 5966 9336
rect 6825 9333 6837 9336
rect 6871 9333 6883 9367
rect 7282 9364 7288 9376
rect 7243 9336 7288 9364
rect 6825 9327 6883 9333
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 10410 9364 10416 9376
rect 10371 9336 10416 9364
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 10870 9364 10876 9376
rect 10783 9336 10876 9364
rect 10870 9324 10876 9336
rect 10928 9364 10934 9376
rect 13078 9364 13084 9376
rect 10928 9336 13084 9364
rect 10928 9324 10934 9336
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 13262 9364 13268 9376
rect 13223 9336 13268 9364
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 14384 9364 14412 9404
rect 18877 9401 18889 9404
rect 18923 9401 18935 9435
rect 18877 9395 18935 9401
rect 19150 9392 19156 9444
rect 19208 9432 19214 9444
rect 19536 9432 19564 9463
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 19208 9404 19564 9432
rect 19208 9392 19214 9404
rect 13780 9336 14412 9364
rect 16117 9367 16175 9373
rect 13780 9324 13786 9336
rect 16117 9333 16129 9367
rect 16163 9364 16175 9367
rect 16669 9367 16727 9373
rect 16669 9364 16681 9367
rect 16163 9336 16681 9364
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 16669 9333 16681 9336
rect 16715 9333 16727 9367
rect 17034 9364 17040 9376
rect 16995 9336 17040 9364
rect 16669 9327 16727 9333
rect 17034 9324 17040 9336
rect 17092 9324 17098 9376
rect 17129 9367 17187 9373
rect 17129 9333 17141 9367
rect 17175 9364 17187 9367
rect 17678 9364 17684 9376
rect 17175 9336 17684 9364
rect 17175 9333 17187 9336
rect 17129 9327 17187 9333
rect 17678 9324 17684 9336
rect 17736 9324 17742 9376
rect 18966 9324 18972 9376
rect 19024 9364 19030 9376
rect 20346 9364 20352 9376
rect 19024 9336 20352 9364
rect 19024 9324 19030 9336
rect 20346 9324 20352 9336
rect 20404 9324 20410 9376
rect 20438 9324 20444 9376
rect 20496 9364 20502 9376
rect 20901 9367 20959 9373
rect 20901 9364 20913 9367
rect 20496 9336 20913 9364
rect 20496 9324 20502 9336
rect 20901 9333 20913 9336
rect 20947 9333 20959 9367
rect 20901 9327 20959 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2832 9132 2973 9160
rect 2832 9120 2838 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 3326 9160 3332 9172
rect 3287 9132 3332 9160
rect 2961 9123 3019 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 4062 9160 4068 9172
rect 3476 9132 3521 9160
rect 4023 9132 4068 9160
rect 3476 9120 3482 9132
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 5077 9163 5135 9169
rect 5077 9160 5089 9163
rect 4764 9132 5089 9160
rect 4764 9120 4770 9132
rect 5077 9129 5089 9132
rect 5123 9129 5135 9163
rect 5077 9123 5135 9129
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 8113 9163 8171 9169
rect 8113 9160 8125 9163
rect 5491 9132 8125 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 8113 9129 8125 9132
rect 8159 9129 8171 9163
rect 8113 9123 8171 9129
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 13998 9160 14004 9172
rect 8536 9132 14004 9160
rect 8536 9120 8542 9132
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14093 9163 14151 9169
rect 14093 9129 14105 9163
rect 14139 9160 14151 9163
rect 14550 9160 14556 9172
rect 14139 9132 14556 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 14550 9120 14556 9132
rect 14608 9160 14614 9172
rect 15010 9160 15016 9172
rect 14608 9132 15016 9160
rect 14608 9120 14614 9132
rect 15010 9120 15016 9132
rect 15068 9120 15074 9172
rect 15289 9163 15347 9169
rect 15289 9129 15301 9163
rect 15335 9160 15347 9163
rect 15562 9160 15568 9172
rect 15335 9132 15568 9160
rect 15335 9129 15347 9132
rect 15289 9123 15347 9129
rect 15562 9120 15568 9132
rect 15620 9120 15626 9172
rect 15657 9163 15715 9169
rect 15657 9129 15669 9163
rect 15703 9160 15715 9163
rect 16206 9160 16212 9172
rect 15703 9132 16212 9160
rect 15703 9129 15715 9132
rect 15657 9123 15715 9129
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 16669 9163 16727 9169
rect 16669 9129 16681 9163
rect 16715 9160 16727 9163
rect 17678 9160 17684 9172
rect 16715 9132 17684 9160
rect 16715 9129 16727 9132
rect 16669 9123 16727 9129
rect 17678 9120 17684 9132
rect 17736 9120 17742 9172
rect 17862 9120 17868 9172
rect 17920 9160 17926 9172
rect 18785 9163 18843 9169
rect 18785 9160 18797 9163
rect 17920 9132 18797 9160
rect 17920 9120 17926 9132
rect 18785 9129 18797 9132
rect 18831 9129 18843 9163
rect 18785 9123 18843 9129
rect 18874 9120 18880 9172
rect 18932 9160 18938 9172
rect 18932 9132 19932 9160
rect 18932 9120 18938 9132
rect 1394 9052 1400 9104
rect 1452 9092 1458 9104
rect 2317 9095 2375 9101
rect 2317 9092 2329 9095
rect 1452 9064 2329 9092
rect 1452 9052 1458 9064
rect 2317 9061 2329 9064
rect 2363 9061 2375 9095
rect 4893 9095 4951 9101
rect 2317 9055 2375 9061
rect 3712 9064 4568 9092
rect 2222 8984 2228 9036
rect 2280 9024 2286 9036
rect 3712 9024 3740 9064
rect 2280 8996 2544 9024
rect 2280 8984 2286 8996
rect 2406 8956 2412 8968
rect 2367 8928 2412 8956
rect 2406 8916 2412 8928
rect 2464 8916 2470 8968
rect 2516 8965 2544 8996
rect 3528 8996 3740 9024
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 2682 8956 2688 8968
rect 2547 8928 2688 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 2682 8916 2688 8928
rect 2740 8956 2746 8968
rect 3528 8965 3556 8996
rect 4246 8984 4252 9036
rect 4304 9024 4310 9036
rect 4433 9027 4491 9033
rect 4433 9024 4445 9027
rect 4304 8996 4445 9024
rect 4304 8984 4310 8996
rect 4433 8993 4445 8996
rect 4479 8993 4491 9027
rect 4540 9024 4568 9064
rect 4893 9061 4905 9095
rect 4939 9092 4951 9095
rect 12618 9092 12624 9104
rect 4939 9064 12624 9092
rect 4939 9061 4951 9064
rect 4893 9055 4951 9061
rect 12618 9052 12624 9064
rect 12676 9052 12682 9104
rect 13078 9052 13084 9104
rect 13136 9092 13142 9104
rect 13136 9064 14412 9092
rect 13136 9052 13142 9064
rect 4540 8996 5672 9024
rect 4433 8987 4491 8993
rect 3513 8959 3571 8965
rect 3513 8956 3525 8959
rect 2740 8928 3525 8956
rect 2740 8916 2746 8928
rect 3513 8925 3525 8928
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 4724 8965 4752 8996
rect 4525 8959 4583 8965
rect 4525 8956 4537 8959
rect 3660 8928 4537 8956
rect 3660 8916 3666 8928
rect 4525 8925 4537 8928
rect 4571 8925 4583 8959
rect 4525 8919 4583 8925
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 5644 8965 5672 8996
rect 5994 8984 6000 9036
rect 6052 9024 6058 9036
rect 6457 9027 6515 9033
rect 6457 9024 6469 9027
rect 6052 8996 6469 9024
rect 6052 8984 6058 8996
rect 6457 8993 6469 8996
rect 6503 8993 6515 9027
rect 6457 8987 6515 8993
rect 6724 9027 6782 9033
rect 6724 8993 6736 9027
rect 6770 9024 6782 9027
rect 7190 9024 7196 9036
rect 6770 8996 7196 9024
rect 6770 8993 6782 8996
rect 6724 8987 6782 8993
rect 7190 8984 7196 8996
rect 7248 9024 7254 9036
rect 7558 9024 7564 9036
rect 7248 8996 7564 9024
rect 7248 8984 7254 8996
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 8202 8984 8208 9036
rect 8260 9024 8266 9036
rect 8481 9027 8539 9033
rect 8481 9024 8493 9027
rect 8260 8996 8493 9024
rect 8260 8984 8266 8996
rect 8481 8993 8493 8996
rect 8527 8993 8539 9027
rect 8481 8987 8539 8993
rect 8570 8984 8576 9036
rect 8628 9024 8634 9036
rect 10594 9024 10600 9036
rect 8628 8996 8673 9024
rect 10555 8996 10600 9024
rect 8628 8984 8634 8996
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 12342 8984 12348 9036
rect 12400 9024 12406 9036
rect 12704 9027 12762 9033
rect 12704 9024 12716 9027
rect 12400 8996 12716 9024
rect 12400 8984 12406 8996
rect 12704 8993 12716 8996
rect 12750 9024 12762 9027
rect 13538 9024 13544 9036
rect 12750 8996 13544 9024
rect 12750 8993 12762 8996
rect 12704 8987 12762 8993
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 14277 9027 14335 9033
rect 14277 8993 14289 9027
rect 14323 8993 14335 9027
rect 14277 8987 14335 8993
rect 5537 8959 5595 8965
rect 5537 8956 5549 8959
rect 4856 8928 5549 8956
rect 4856 8916 4862 8928
rect 5537 8925 5549 8928
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8925 5687 8959
rect 5629 8919 5687 8925
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 7708 8928 7972 8956
rect 7708 8916 7714 8928
rect 3970 8848 3976 8900
rect 4028 8888 4034 8900
rect 4893 8891 4951 8897
rect 4893 8888 4905 8891
rect 4028 8860 4905 8888
rect 4028 8848 4034 8860
rect 4893 8857 4905 8860
rect 4939 8857 4951 8891
rect 4893 8851 4951 8857
rect 7466 8848 7472 8900
rect 7524 8888 7530 8900
rect 7837 8891 7895 8897
rect 7837 8888 7849 8891
rect 7524 8860 7849 8888
rect 7524 8848 7530 8860
rect 7837 8857 7849 8860
rect 7883 8857 7895 8891
rect 7944 8888 7972 8928
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8665 8959 8723 8965
rect 8665 8956 8677 8959
rect 8352 8928 8677 8956
rect 8352 8916 8358 8928
rect 8665 8925 8677 8928
rect 8711 8925 8723 8959
rect 8665 8919 8723 8925
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 12158 8956 12164 8968
rect 8812 8928 12164 8956
rect 8812 8916 8818 8928
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 12434 8956 12440 8968
rect 12395 8928 12440 8956
rect 12434 8916 12440 8928
rect 12492 8916 12498 8968
rect 12250 8888 12256 8900
rect 7944 8860 12256 8888
rect 7837 8851 7895 8857
rect 12250 8848 12256 8860
rect 12308 8848 12314 8900
rect 14292 8888 14320 8987
rect 13372 8860 14320 8888
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 9490 8820 9496 8832
rect 4120 8792 9496 8820
rect 4120 8780 4126 8792
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 11882 8820 11888 8832
rect 11843 8792 11888 8820
rect 11882 8780 11888 8792
rect 11940 8820 11946 8832
rect 13372 8820 13400 8860
rect 11940 8792 13400 8820
rect 11940 8780 11946 8792
rect 13722 8780 13728 8832
rect 13780 8820 13786 8832
rect 13817 8823 13875 8829
rect 13817 8820 13829 8823
rect 13780 8792 13829 8820
rect 13780 8780 13786 8792
rect 13817 8789 13829 8792
rect 13863 8789 13875 8823
rect 14384 8820 14412 9064
rect 14458 9052 14464 9104
rect 14516 9092 14522 9104
rect 14516 9064 16896 9092
rect 14516 9052 14522 9064
rect 14642 8984 14648 9036
rect 14700 9024 14706 9036
rect 16574 9024 16580 9036
rect 14700 8996 16580 9024
rect 14700 8984 14706 8996
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 15436 8928 15761 8956
rect 15436 8916 15442 8928
rect 15749 8925 15761 8928
rect 15795 8925 15807 8959
rect 15749 8919 15807 8925
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 16482 8956 16488 8968
rect 15896 8928 16488 8956
rect 15896 8916 15902 8928
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 16868 8965 16896 9064
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 17310 9092 17316 9104
rect 17092 9064 17316 9092
rect 17092 9052 17098 9064
rect 17310 9052 17316 9064
rect 17368 9092 17374 9104
rect 19794 9092 19800 9104
rect 17368 9064 19800 9092
rect 17368 9052 17374 9064
rect 19794 9052 19800 9064
rect 19852 9052 19858 9104
rect 19904 9092 19932 9132
rect 20162 9120 20168 9172
rect 20220 9160 20226 9172
rect 20257 9163 20315 9169
rect 20257 9160 20269 9163
rect 20220 9132 20269 9160
rect 20220 9120 20226 9132
rect 20257 9129 20269 9132
rect 20303 9129 20315 9163
rect 20257 9123 20315 9129
rect 20346 9092 20352 9104
rect 19904 9064 20352 9092
rect 20346 9052 20352 9064
rect 20404 9052 20410 9104
rect 17672 9027 17730 9033
rect 17672 8993 17684 9027
rect 17718 9024 17730 9027
rect 17954 9024 17960 9036
rect 17718 8996 17960 9024
rect 17718 8993 17730 8996
rect 17672 8987 17730 8993
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 19058 9024 19064 9036
rect 19019 8996 19064 9024
rect 19058 8984 19064 8996
rect 19116 8984 19122 9036
rect 20165 9027 20223 9033
rect 20165 8993 20177 9027
rect 20211 9024 20223 9027
rect 20901 9027 20959 9033
rect 20901 9024 20913 9027
rect 20211 8996 20913 9024
rect 20211 8993 20223 8996
rect 20165 8987 20223 8993
rect 20901 8993 20913 8996
rect 20947 8993 20959 9027
rect 20901 8987 20959 8993
rect 16761 8959 16819 8965
rect 16761 8925 16773 8959
rect 16807 8925 16819 8959
rect 16761 8919 16819 8925
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8925 16911 8959
rect 17402 8956 17408 8968
rect 17363 8928 17408 8956
rect 16853 8919 16911 8925
rect 15194 8848 15200 8900
rect 15252 8888 15258 8900
rect 16301 8891 16359 8897
rect 16301 8888 16313 8891
rect 15252 8860 16313 8888
rect 15252 8848 15258 8860
rect 16301 8857 16313 8860
rect 16347 8857 16359 8891
rect 16776 8888 16804 8919
rect 17402 8916 17408 8928
rect 17460 8916 17466 8968
rect 19334 8956 19340 8968
rect 19295 8928 19340 8956
rect 19334 8916 19340 8928
rect 19392 8916 19398 8968
rect 20438 8956 20444 8968
rect 20399 8928 20444 8956
rect 20438 8916 20444 8928
rect 20496 8916 20502 8968
rect 16942 8888 16948 8900
rect 16776 8860 16948 8888
rect 16301 8851 16359 8857
rect 16942 8848 16948 8860
rect 17000 8888 17006 8900
rect 17218 8888 17224 8900
rect 17000 8860 17224 8888
rect 17000 8848 17006 8860
rect 17218 8848 17224 8860
rect 17276 8848 17282 8900
rect 19150 8820 19156 8832
rect 14384 8792 19156 8820
rect 13817 8783 13875 8789
rect 19150 8780 19156 8792
rect 19208 8780 19214 8832
rect 19797 8823 19855 8829
rect 19797 8789 19809 8823
rect 19843 8820 19855 8823
rect 20070 8820 20076 8832
rect 19843 8792 20076 8820
rect 19843 8789 19855 8792
rect 19797 8783 19855 8789
rect 20070 8780 20076 8792
rect 20128 8780 20134 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2682 8576 2688 8628
rect 2740 8616 2746 8628
rect 3145 8619 3203 8625
rect 3145 8616 3157 8619
rect 2740 8588 3157 8616
rect 2740 8576 2746 8588
rect 3145 8585 3157 8588
rect 3191 8585 3203 8619
rect 3602 8616 3608 8628
rect 3563 8588 3608 8616
rect 3145 8579 3203 8585
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 3804 8588 4445 8616
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 3804 8548 3832 8588
rect 4433 8585 4445 8588
rect 4479 8585 4491 8619
rect 4433 8579 4491 8585
rect 4617 8619 4675 8625
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 5810 8616 5816 8628
rect 4663 8588 5816 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 6822 8616 6828 8628
rect 6783 8588 6828 8616
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7650 8616 7656 8628
rect 6932 8588 7656 8616
rect 3292 8520 3832 8548
rect 3292 8508 3298 8520
rect 3878 8508 3884 8560
rect 3936 8548 3942 8560
rect 6932 8548 6960 8588
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 9398 8616 9404 8628
rect 7883 8588 9404 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9953 8619 10011 8625
rect 9953 8585 9965 8619
rect 9999 8616 10011 8619
rect 10134 8616 10140 8628
rect 9999 8588 10140 8616
rect 9999 8585 10011 8588
rect 9953 8579 10011 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 11146 8616 11152 8628
rect 10560 8588 11152 8616
rect 10560 8576 10566 8588
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11333 8619 11391 8625
rect 11333 8585 11345 8619
rect 11379 8616 11391 8619
rect 12618 8616 12624 8628
rect 11379 8588 12624 8616
rect 11379 8585 11391 8588
rect 11333 8579 11391 8585
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 13814 8616 13820 8628
rect 13775 8588 13820 8616
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 15473 8619 15531 8625
rect 15473 8616 15485 8619
rect 14056 8588 15485 8616
rect 14056 8576 14062 8588
rect 15473 8585 15485 8588
rect 15519 8616 15531 8619
rect 15838 8616 15844 8628
rect 15519 8588 15844 8616
rect 15519 8585 15531 8588
rect 15473 8579 15531 8585
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 16850 8616 16856 8628
rect 15948 8588 16856 8616
rect 3936 8520 6960 8548
rect 3936 8508 3942 8520
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 7742 8548 7748 8560
rect 7064 8520 7748 8548
rect 7064 8508 7070 8520
rect 7742 8508 7748 8520
rect 7800 8548 7806 8560
rect 8849 8551 8907 8557
rect 8849 8548 8861 8551
rect 7800 8520 8861 8548
rect 7800 8508 7806 8520
rect 8849 8517 8861 8520
rect 8895 8517 8907 8551
rect 8849 8511 8907 8517
rect 9125 8551 9183 8557
rect 9125 8517 9137 8551
rect 9171 8548 9183 8551
rect 10042 8548 10048 8560
rect 9171 8520 10048 8548
rect 9171 8517 9183 8520
rect 9125 8511 9183 8517
rect 10042 8508 10048 8520
rect 10100 8508 10106 8560
rect 10226 8508 10232 8560
rect 10284 8548 10290 8560
rect 10284 8520 10640 8548
rect 10284 8508 10290 8520
rect 1670 8440 1676 8492
rect 1728 8480 1734 8492
rect 1765 8483 1823 8489
rect 1765 8480 1777 8483
rect 1728 8452 1777 8480
rect 1728 8440 1734 8452
rect 1765 8449 1777 8452
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 3786 8440 3792 8492
rect 3844 8480 3850 8492
rect 4157 8483 4215 8489
rect 4157 8480 4169 8483
rect 3844 8452 4169 8480
rect 3844 8440 3850 8452
rect 4157 8449 4169 8452
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8480 5135 8483
rect 5166 8480 5172 8492
rect 5123 8452 5172 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5442 8480 5448 8492
rect 5307 8452 5448 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 6178 8480 6184 8492
rect 5583 8452 6184 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 7558 8480 7564 8492
rect 7515 8452 7564 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 8478 8480 8484 8492
rect 8439 8452 8484 8480
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 9677 8483 9735 8489
rect 9677 8480 9689 8483
rect 8996 8452 9689 8480
rect 8996 8440 9002 8452
rect 9677 8449 9689 8452
rect 9723 8449 9735 8483
rect 10410 8480 10416 8492
rect 10371 8452 10416 8480
rect 9677 8443 9735 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10612 8489 10640 8520
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 11793 8483 11851 8489
rect 11793 8480 11805 8483
rect 11204 8452 11805 8480
rect 11204 8440 11210 8452
rect 11793 8449 11805 8452
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8480 12035 8483
rect 12342 8480 12348 8492
rect 12023 8452 12348 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 13832 8480 13860 8576
rect 15194 8508 15200 8560
rect 15252 8548 15258 8560
rect 15948 8548 15976 8588
rect 16850 8576 16856 8588
rect 16908 8576 16914 8628
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 19242 8616 19248 8628
rect 18932 8588 19104 8616
rect 18932 8576 18938 8588
rect 15252 8520 15976 8548
rect 16393 8551 16451 8557
rect 15252 8508 15258 8520
rect 16393 8517 16405 8551
rect 16439 8548 16451 8551
rect 17310 8548 17316 8560
rect 16439 8520 17316 8548
rect 16439 8517 16451 8520
rect 16393 8511 16451 8517
rect 17310 8508 17316 8520
rect 17368 8508 17374 8560
rect 17589 8551 17647 8557
rect 17589 8517 17601 8551
rect 17635 8548 17647 8551
rect 18969 8551 19027 8557
rect 18969 8548 18981 8551
rect 17635 8520 18981 8548
rect 17635 8517 17647 8520
rect 17589 8511 17647 8517
rect 18969 8517 18981 8520
rect 19015 8517 19027 8551
rect 18969 8511 19027 8517
rect 13832 8452 14228 8480
rect 2314 8372 2320 8424
rect 2372 8412 2378 8424
rect 2498 8412 2504 8424
rect 2372 8384 2504 8412
rect 2372 8372 2378 8384
rect 2498 8372 2504 8384
rect 2556 8412 2562 8424
rect 5997 8415 6055 8421
rect 5997 8412 6009 8415
rect 2556 8384 6009 8412
rect 2556 8372 2562 8384
rect 5997 8381 6009 8384
rect 6043 8381 6055 8415
rect 5997 8375 6055 8381
rect 6822 8372 6828 8424
rect 6880 8412 6886 8424
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 6880 8384 7297 8412
rect 6880 8372 6886 8384
rect 7285 8381 7297 8384
rect 7331 8381 7343 8415
rect 7285 8375 7343 8381
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8412 9091 8415
rect 11882 8412 11888 8424
rect 9079 8384 11888 8412
rect 9079 8381 9091 8384
rect 9033 8375 9091 8381
rect 11882 8372 11888 8384
rect 11940 8372 11946 8424
rect 12434 8412 12440 8424
rect 12347 8384 12440 8412
rect 12434 8372 12440 8384
rect 12492 8412 12498 8424
rect 14093 8415 14151 8421
rect 14093 8412 14105 8415
rect 12492 8384 14105 8412
rect 12492 8372 12498 8384
rect 14093 8381 14105 8384
rect 14139 8381 14151 8415
rect 14200 8412 14228 8452
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16816 8452 16865 8480
rect 16816 8440 16822 8452
rect 16853 8449 16865 8452
rect 16899 8480 16911 8483
rect 17037 8483 17095 8489
rect 16899 8452 16988 8480
rect 16899 8449 16911 8452
rect 16853 8443 16911 8449
rect 14349 8415 14407 8421
rect 14349 8412 14361 8415
rect 14200 8384 14361 8412
rect 14093 8375 14151 8381
rect 14349 8381 14361 8384
rect 14395 8381 14407 8415
rect 16960 8412 16988 8452
rect 17037 8449 17049 8483
rect 17083 8480 17095 8483
rect 17218 8480 17224 8492
rect 17083 8452 17224 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 17218 8440 17224 8452
rect 17276 8440 17282 8492
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 18693 8483 18751 8489
rect 18693 8480 18705 8483
rect 17920 8452 18705 8480
rect 17920 8440 17926 8452
rect 18693 8449 18705 8452
rect 18739 8449 18751 8483
rect 19076 8480 19104 8588
rect 18693 8443 18751 8449
rect 18800 8452 19104 8480
rect 19168 8588 19248 8616
rect 19168 8480 19196 8588
rect 19242 8576 19248 8588
rect 19300 8576 19306 8628
rect 19337 8619 19395 8625
rect 19337 8585 19349 8619
rect 19383 8616 19395 8619
rect 19978 8616 19984 8628
rect 19383 8588 19984 8616
rect 19383 8585 19395 8588
rect 19337 8579 19395 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 19168 8452 19288 8480
rect 17126 8412 17132 8424
rect 16960 8384 17132 8412
rect 14349 8375 14407 8381
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 17405 8415 17463 8421
rect 17405 8381 17417 8415
rect 17451 8412 17463 8415
rect 17494 8412 17500 8424
rect 17451 8384 17500 8412
rect 17451 8381 17463 8384
rect 17405 8375 17463 8381
rect 17494 8372 17500 8384
rect 17552 8372 17558 8424
rect 18601 8415 18659 8421
rect 18601 8381 18613 8415
rect 18647 8412 18659 8415
rect 18800 8412 18828 8452
rect 18647 8384 18828 8412
rect 18647 8381 18659 8384
rect 18601 8375 18659 8381
rect 18874 8372 18880 8424
rect 18932 8412 18938 8424
rect 19153 8415 19211 8421
rect 19153 8412 19165 8415
rect 18932 8384 19165 8412
rect 18932 8372 18938 8384
rect 19153 8381 19165 8384
rect 19199 8381 19211 8415
rect 19260 8412 19288 8452
rect 19260 8384 19380 8412
rect 19153 8375 19211 8381
rect 2032 8347 2090 8353
rect 2032 8313 2044 8347
rect 2078 8344 2090 8347
rect 2078 8316 2360 8344
rect 2078 8313 2090 8316
rect 2032 8307 2090 8313
rect 2332 8276 2360 8316
rect 2406 8304 2412 8356
rect 2464 8344 2470 8356
rect 6454 8344 6460 8356
rect 2464 8316 5672 8344
rect 2464 8304 2470 8316
rect 2590 8276 2596 8288
rect 2332 8248 2596 8276
rect 2590 8236 2596 8248
rect 2648 8276 2654 8288
rect 3234 8276 3240 8288
rect 2648 8248 3240 8276
rect 2648 8236 2654 8248
rect 3234 8236 3240 8248
rect 3292 8276 3298 8288
rect 3786 8276 3792 8288
rect 3292 8248 3792 8276
rect 3292 8236 3298 8248
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 3970 8276 3976 8288
rect 3931 8248 3976 8276
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 4065 8279 4123 8285
rect 4065 8245 4077 8279
rect 4111 8276 4123 8279
rect 4430 8276 4436 8288
rect 4111 8248 4436 8276
rect 4111 8245 4123 8248
rect 4065 8239 4123 8245
rect 4430 8236 4436 8248
rect 4488 8236 4494 8288
rect 4982 8276 4988 8288
rect 4943 8248 4988 8276
rect 4982 8236 4988 8248
rect 5040 8236 5046 8288
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 5644 8285 5672 8316
rect 6380 8316 6460 8344
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 5224 8248 5457 8276
rect 5224 8236 5230 8248
rect 5445 8245 5457 8248
rect 5491 8245 5503 8279
rect 5445 8239 5503 8245
rect 5629 8279 5687 8285
rect 5629 8245 5641 8279
rect 5675 8245 5687 8279
rect 5629 8239 5687 8245
rect 5810 8236 5816 8288
rect 5868 8276 5874 8288
rect 6089 8279 6147 8285
rect 6089 8276 6101 8279
rect 5868 8248 6101 8276
rect 5868 8236 5874 8248
rect 6089 8245 6101 8248
rect 6135 8276 6147 8279
rect 6380 8276 6408 8316
rect 6454 8304 6460 8316
rect 6512 8304 6518 8356
rect 6546 8304 6552 8356
rect 6604 8344 6610 8356
rect 7193 8347 7251 8353
rect 7193 8344 7205 8347
rect 6604 8316 7205 8344
rect 6604 8304 6610 8316
rect 7193 8313 7205 8316
rect 7239 8313 7251 8347
rect 7193 8307 7251 8313
rect 7374 8304 7380 8356
rect 7432 8344 7438 8356
rect 8205 8347 8263 8353
rect 8205 8344 8217 8347
rect 7432 8316 8217 8344
rect 7432 8304 7438 8316
rect 8205 8313 8217 8316
rect 8251 8313 8263 8347
rect 8205 8307 8263 8313
rect 9493 8347 9551 8353
rect 9493 8313 9505 8347
rect 9539 8344 9551 8347
rect 10686 8344 10692 8356
rect 9539 8316 10692 8344
rect 9539 8313 9551 8316
rect 9493 8307 9551 8313
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 10781 8347 10839 8353
rect 10781 8313 10793 8347
rect 10827 8344 10839 8347
rect 11054 8344 11060 8356
rect 10827 8316 11060 8344
rect 10827 8313 10839 8316
rect 10781 8307 10839 8313
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 12704 8347 12762 8353
rect 12704 8313 12716 8347
rect 12750 8344 12762 8347
rect 12802 8344 12808 8356
rect 12750 8316 12808 8344
rect 12750 8313 12762 8316
rect 12704 8307 12762 8313
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 12894 8304 12900 8356
rect 12952 8344 12958 8356
rect 16574 8344 16580 8356
rect 12952 8316 13584 8344
rect 12952 8304 12958 8316
rect 6135 8248 6408 8276
rect 6135 8245 6147 8248
rect 6089 8239 6147 8245
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 8297 8279 8355 8285
rect 8297 8276 8309 8279
rect 6696 8248 8309 8276
rect 6696 8236 6702 8248
rect 8297 8245 8309 8248
rect 8343 8245 8355 8279
rect 8297 8239 8355 8245
rect 9585 8279 9643 8285
rect 9585 8245 9597 8279
rect 9631 8276 9643 8279
rect 10226 8276 10232 8288
rect 9631 8248 10232 8276
rect 9631 8245 9643 8248
rect 9585 8239 9643 8245
rect 10226 8236 10232 8248
rect 10284 8236 10290 8288
rect 10318 8236 10324 8288
rect 10376 8276 10382 8288
rect 11701 8279 11759 8285
rect 11701 8276 11713 8279
rect 10376 8248 11713 8276
rect 10376 8236 10382 8248
rect 11701 8245 11713 8248
rect 11747 8276 11759 8279
rect 13446 8276 13452 8288
rect 11747 8248 13452 8276
rect 11747 8245 11759 8248
rect 11701 8239 11759 8245
rect 13446 8236 13452 8248
rect 13504 8236 13510 8288
rect 13556 8276 13584 8316
rect 14568 8316 16580 8344
rect 14568 8276 14596 8316
rect 16574 8304 16580 8316
rect 16632 8304 16638 8356
rect 16758 8344 16764 8356
rect 16719 8316 16764 8344
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 19058 8344 19064 8356
rect 18156 8316 19064 8344
rect 15746 8276 15752 8288
rect 13556 8248 14596 8276
rect 15707 8248 15752 8276
rect 15746 8236 15752 8248
rect 15804 8236 15810 8288
rect 15838 8236 15844 8288
rect 15896 8276 15902 8288
rect 17034 8276 17040 8288
rect 15896 8248 17040 8276
rect 15896 8236 15902 8248
rect 17034 8236 17040 8248
rect 17092 8276 17098 8288
rect 17862 8276 17868 8288
rect 17092 8248 17868 8276
rect 17092 8236 17098 8248
rect 17862 8236 17868 8248
rect 17920 8236 17926 8288
rect 18156 8285 18184 8316
rect 19058 8304 19064 8316
rect 19116 8304 19122 8356
rect 19352 8344 19380 8384
rect 19426 8372 19432 8424
rect 19484 8412 19490 8424
rect 19705 8415 19763 8421
rect 19705 8412 19717 8415
rect 19484 8384 19717 8412
rect 19484 8372 19490 8384
rect 19705 8381 19717 8384
rect 19751 8381 19763 8415
rect 19705 8375 19763 8381
rect 19972 8415 20030 8421
rect 19972 8381 19984 8415
rect 20018 8412 20030 8415
rect 20438 8412 20444 8424
rect 20018 8384 20444 8412
rect 20018 8381 20030 8384
rect 19972 8375 20030 8381
rect 20438 8372 20444 8384
rect 20496 8372 20502 8424
rect 19352 8316 21128 8344
rect 18141 8279 18199 8285
rect 18141 8245 18153 8279
rect 18187 8245 18199 8279
rect 18141 8239 18199 8245
rect 18506 8236 18512 8288
rect 18564 8276 18570 8288
rect 18969 8279 19027 8285
rect 18564 8248 18609 8276
rect 18564 8236 18570 8248
rect 18969 8245 18981 8279
rect 19015 8276 19027 8279
rect 20438 8276 20444 8288
rect 19015 8248 20444 8276
rect 19015 8245 19027 8248
rect 18969 8239 19027 8245
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 21100 8285 21128 8316
rect 21085 8279 21143 8285
rect 21085 8245 21097 8279
rect 21131 8245 21143 8279
rect 21085 8239 21143 8245
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 4982 8072 4988 8084
rect 3559 8044 4988 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5077 8075 5135 8081
rect 5077 8041 5089 8075
rect 5123 8072 5135 8075
rect 5350 8072 5356 8084
rect 5123 8044 5356 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 6546 8072 6552 8084
rect 6507 8044 6552 8072
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 9306 8072 9312 8084
rect 9267 8044 9312 8072
rect 9306 8032 9312 8044
rect 9364 8032 9370 8084
rect 10042 8072 10048 8084
rect 10003 8044 10048 8072
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 10137 8075 10195 8081
rect 10137 8041 10149 8075
rect 10183 8072 10195 8075
rect 10410 8072 10416 8084
rect 10183 8044 10416 8072
rect 10183 8041 10195 8044
rect 10137 8035 10195 8041
rect 10410 8032 10416 8044
rect 10468 8032 10474 8084
rect 10686 8072 10692 8084
rect 10647 8044 10692 8072
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 11054 8072 11060 8084
rect 11015 8044 11060 8072
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 12526 8072 12532 8084
rect 12487 8044 12532 8072
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 13173 8075 13231 8081
rect 12676 8044 12721 8072
rect 12676 8032 12682 8044
rect 13173 8041 13185 8075
rect 13219 8072 13231 8075
rect 13262 8072 13268 8084
rect 13219 8044 13268 8072
rect 13219 8041 13231 8044
rect 13173 8035 13231 8041
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 14185 8075 14243 8081
rect 14185 8072 14197 8075
rect 13679 8044 14197 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 14185 8041 14197 8044
rect 14231 8041 14243 8075
rect 14185 8035 14243 8041
rect 14458 8032 14464 8084
rect 14516 8072 14522 8084
rect 15838 8072 15844 8084
rect 14516 8044 15844 8072
rect 14516 8032 14522 8044
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 15930 8032 15936 8084
rect 15988 8072 15994 8084
rect 16390 8072 16396 8084
rect 15988 8044 16396 8072
rect 15988 8032 15994 8044
rect 16390 8032 16396 8044
rect 16448 8072 16454 8084
rect 16669 8075 16727 8081
rect 16669 8072 16681 8075
rect 16448 8044 16681 8072
rect 16448 8032 16454 8044
rect 16669 8041 16681 8044
rect 16715 8041 16727 8075
rect 17402 8072 17408 8084
rect 16669 8035 16727 8041
rect 16960 8044 17408 8072
rect 4433 8007 4491 8013
rect 4433 7973 4445 8007
rect 4479 8004 4491 8007
rect 4890 8004 4896 8016
rect 4479 7976 4896 8004
rect 4479 7973 4491 7976
rect 4433 7967 4491 7973
rect 4890 7964 4896 7976
rect 4948 7964 4954 8016
rect 5258 7964 5264 8016
rect 5316 8004 5322 8016
rect 5445 8007 5503 8013
rect 5445 8004 5457 8007
rect 5316 7976 5457 8004
rect 5316 7964 5322 7976
rect 5445 7973 5457 7976
rect 5491 7973 5503 8007
rect 5445 7967 5503 7973
rect 8196 8007 8254 8013
rect 8196 7973 8208 8007
rect 8242 8004 8254 8007
rect 8938 8004 8944 8016
rect 8242 7976 8944 8004
rect 8242 7973 8254 7976
rect 8196 7967 8254 7973
rect 8938 7964 8944 7976
rect 8996 7964 9002 8016
rect 2038 7896 2044 7948
rect 2096 7936 2102 7948
rect 2409 7939 2467 7945
rect 2409 7936 2421 7939
rect 2096 7908 2421 7936
rect 2096 7896 2102 7908
rect 2409 7905 2421 7908
rect 2455 7905 2467 7939
rect 2409 7899 2467 7905
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7936 2559 7939
rect 3418 7936 3424 7948
rect 2547 7908 3424 7936
rect 2547 7905 2559 7908
rect 2501 7899 2559 7905
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 4525 7939 4583 7945
rect 4525 7905 4537 7939
rect 4571 7936 4583 7939
rect 4982 7936 4988 7948
rect 4571 7908 4988 7936
rect 4571 7905 4583 7908
rect 4525 7899 4583 7905
rect 4982 7896 4988 7908
rect 5040 7896 5046 7948
rect 6089 7939 6147 7945
rect 6089 7905 6101 7939
rect 6135 7936 6147 7939
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 6135 7908 6929 7936
rect 6135 7905 6147 7908
rect 6089 7899 6147 7905
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7936 7987 7939
rect 9030 7936 9036 7948
rect 7975 7908 9036 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 9030 7896 9036 7908
rect 9088 7896 9094 7948
rect 9324 7936 9352 8032
rect 9490 7964 9496 8016
rect 9548 8004 9554 8016
rect 11149 8007 11207 8013
rect 11149 8004 11161 8007
rect 9548 7976 11161 8004
rect 9548 7964 9554 7976
rect 11149 7973 11161 7976
rect 11195 7973 11207 8007
rect 11149 7967 11207 7973
rect 11882 7964 11888 8016
rect 11940 8004 11946 8016
rect 15194 8004 15200 8016
rect 11940 7976 15200 8004
rect 11940 7964 11946 7976
rect 15194 7964 15200 7976
rect 15252 7964 15258 8016
rect 15562 8013 15568 8016
rect 15556 8004 15568 8013
rect 15523 7976 15568 8004
rect 15556 7967 15568 7976
rect 15562 7964 15568 7967
rect 15620 7964 15626 8016
rect 9324 7908 10272 7936
rect 2682 7868 2688 7880
rect 2643 7840 2688 7868
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 3786 7828 3792 7880
rect 3844 7868 3850 7880
rect 4709 7871 4767 7877
rect 4709 7868 4721 7871
rect 3844 7840 4721 7868
rect 3844 7828 3850 7840
rect 4709 7837 4721 7840
rect 4755 7868 4767 7871
rect 5166 7868 5172 7880
rect 4755 7840 5172 7868
rect 4755 7837 4767 7840
rect 4709 7831 4767 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 5258 7828 5264 7880
rect 5316 7868 5322 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5316 7840 5549 7868
rect 5316 7828 5322 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 5629 7831 5687 7837
rect 5736 7840 7021 7868
rect 4065 7803 4123 7809
rect 4065 7769 4077 7803
rect 4111 7800 4123 7803
rect 4798 7800 4804 7812
rect 4111 7772 4804 7800
rect 4111 7769 4123 7772
rect 4065 7763 4123 7769
rect 4798 7760 4804 7772
rect 4856 7760 4862 7812
rect 5442 7760 5448 7812
rect 5500 7800 5506 7812
rect 5644 7800 5672 7831
rect 5500 7772 5672 7800
rect 5500 7760 5506 7772
rect 2041 7735 2099 7741
rect 2041 7701 2053 7735
rect 2087 7732 2099 7735
rect 2590 7732 2596 7744
rect 2087 7704 2596 7732
rect 2087 7701 2099 7704
rect 2041 7695 2099 7701
rect 2590 7692 2596 7704
rect 2648 7692 2654 7744
rect 2958 7692 2964 7744
rect 3016 7732 3022 7744
rect 3786 7732 3792 7744
rect 3016 7704 3792 7732
rect 3016 7692 3022 7704
rect 3786 7692 3792 7704
rect 3844 7732 3850 7744
rect 5736 7732 5764 7840
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7190 7868 7196 7880
rect 7151 7840 7196 7868
rect 7009 7831 7067 7837
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 10134 7868 10140 7880
rect 9180 7840 10140 7868
rect 9180 7828 9186 7840
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10244 7877 10272 7908
rect 10962 7896 10968 7948
rect 11020 7936 11026 7948
rect 11020 7908 11284 7936
rect 11020 7896 11026 7908
rect 11256 7877 11284 7908
rect 11606 7896 11612 7948
rect 11664 7936 11670 7948
rect 12618 7936 12624 7948
rect 11664 7908 12624 7936
rect 11664 7896 11670 7908
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 12710 7896 12716 7948
rect 12768 7936 12774 7948
rect 13262 7936 13268 7948
rect 12768 7908 13268 7936
rect 12768 7896 12774 7908
rect 13262 7896 13268 7908
rect 13320 7896 13326 7948
rect 13446 7896 13452 7948
rect 13504 7936 13510 7948
rect 13541 7939 13599 7945
rect 13541 7936 13553 7939
rect 13504 7908 13553 7936
rect 13504 7896 13510 7908
rect 13541 7905 13553 7908
rect 13587 7905 13599 7939
rect 13541 7899 13599 7905
rect 14553 7939 14611 7945
rect 14553 7905 14565 7939
rect 14599 7936 14611 7939
rect 15010 7936 15016 7948
rect 14599 7908 15016 7936
rect 14599 7905 14611 7908
rect 14553 7899 14611 7905
rect 15010 7896 15016 7908
rect 15068 7896 15074 7948
rect 16960 7945 16988 8044
rect 17402 8032 17408 8044
rect 17460 8072 17466 8084
rect 18509 8075 18567 8081
rect 18509 8072 18521 8075
rect 17460 8044 18521 8072
rect 17460 8032 17466 8044
rect 18509 8041 18521 8044
rect 18555 8072 18567 8075
rect 19426 8072 19432 8084
rect 18555 8044 19432 8072
rect 18555 8041 18567 8044
rect 18509 8035 18567 8041
rect 19426 8032 19432 8044
rect 19484 8032 19490 8084
rect 19610 8032 19616 8084
rect 19668 8072 19674 8084
rect 20441 8075 20499 8081
rect 20441 8072 20453 8075
rect 19668 8044 20453 8072
rect 19668 8032 19674 8044
rect 20441 8041 20453 8044
rect 20487 8041 20499 8075
rect 20441 8035 20499 8041
rect 17218 8013 17224 8016
rect 17212 8004 17224 8013
rect 17052 7976 17224 8004
rect 15289 7939 15347 7945
rect 15289 7905 15301 7939
rect 15335 7936 15347 7939
rect 16945 7939 17003 7945
rect 16945 7936 16957 7939
rect 15335 7908 16957 7936
rect 15335 7905 15347 7908
rect 15289 7899 15347 7905
rect 16945 7905 16957 7908
rect 16991 7905 17003 7939
rect 16945 7899 17003 7905
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 12802 7868 12808 7880
rect 12715 7840 12808 7868
rect 11241 7831 11299 7837
rect 12802 7828 12808 7840
rect 12860 7868 12866 7880
rect 13722 7868 13728 7880
rect 12860 7840 13728 7868
rect 12860 7828 12866 7840
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7837 14703 7871
rect 14826 7868 14832 7880
rect 14787 7840 14832 7868
rect 14645 7831 14703 7837
rect 9677 7803 9735 7809
rect 9677 7769 9689 7803
rect 9723 7800 9735 7803
rect 12161 7803 12219 7809
rect 9723 7772 12112 7800
rect 9723 7769 9735 7772
rect 9677 7763 9735 7769
rect 3844 7704 5764 7732
rect 3844 7692 3850 7704
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 10594 7732 10600 7744
rect 6972 7704 10600 7732
rect 6972 7692 6978 7704
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 12084 7732 12112 7772
rect 12161 7769 12173 7803
rect 12207 7800 12219 7803
rect 13170 7800 13176 7812
rect 12207 7772 13176 7800
rect 12207 7769 12219 7772
rect 12161 7763 12219 7769
rect 13170 7760 13176 7772
rect 13228 7760 13234 7812
rect 13262 7760 13268 7812
rect 13320 7800 13326 7812
rect 14458 7800 14464 7812
rect 13320 7772 14464 7800
rect 13320 7760 13326 7772
rect 14458 7760 14464 7772
rect 14516 7760 14522 7812
rect 13998 7732 14004 7744
rect 12084 7704 14004 7732
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 14660 7732 14688 7831
rect 14826 7828 14832 7840
rect 14884 7828 14890 7880
rect 16850 7828 16856 7880
rect 16908 7868 16914 7880
rect 17052 7868 17080 7976
rect 17212 7967 17224 7976
rect 17218 7964 17224 7967
rect 17276 7964 17282 8016
rect 17862 7964 17868 8016
rect 17920 8004 17926 8016
rect 17920 7976 20300 8004
rect 17920 7964 17926 7976
rect 18857 7939 18915 7945
rect 18857 7936 18869 7939
rect 16908 7840 17080 7868
rect 18340 7908 18869 7936
rect 16908 7828 16914 7840
rect 17678 7732 17684 7744
rect 14660 7704 17684 7732
rect 17678 7692 17684 7704
rect 17736 7692 17742 7744
rect 17862 7692 17868 7744
rect 17920 7732 17926 7744
rect 18340 7741 18368 7908
rect 18857 7905 18869 7908
rect 18903 7936 18915 7939
rect 19150 7936 19156 7948
rect 18903 7908 19156 7936
rect 18903 7905 18915 7908
rect 18857 7899 18915 7905
rect 19150 7896 19156 7908
rect 19208 7896 19214 7948
rect 20272 7945 20300 7976
rect 20257 7939 20315 7945
rect 20257 7905 20269 7939
rect 20303 7905 20315 7939
rect 20257 7899 20315 7905
rect 18509 7871 18567 7877
rect 18509 7837 18521 7871
rect 18555 7868 18567 7871
rect 18601 7871 18659 7877
rect 18601 7868 18613 7871
rect 18555 7840 18613 7868
rect 18555 7837 18567 7840
rect 18509 7831 18567 7837
rect 18601 7837 18613 7840
rect 18647 7837 18659 7871
rect 20898 7868 20904 7880
rect 20859 7840 20904 7868
rect 18601 7831 18659 7837
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 18325 7735 18383 7741
rect 18325 7732 18337 7735
rect 17920 7704 18337 7732
rect 17920 7692 17926 7704
rect 18325 7701 18337 7704
rect 18371 7701 18383 7735
rect 18325 7695 18383 7701
rect 19242 7692 19248 7744
rect 19300 7732 19306 7744
rect 19981 7735 20039 7741
rect 19981 7732 19993 7735
rect 19300 7704 19993 7732
rect 19300 7692 19306 7704
rect 19981 7701 19993 7704
rect 20027 7701 20039 7735
rect 19981 7695 20039 7701
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 2225 7531 2283 7537
rect 2225 7497 2237 7531
rect 2271 7528 2283 7531
rect 3050 7528 3056 7540
rect 2271 7500 3056 7528
rect 2271 7497 2283 7500
rect 2225 7491 2283 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 4433 7531 4491 7537
rect 4433 7528 4445 7531
rect 4304 7500 4445 7528
rect 4304 7488 4310 7500
rect 4433 7497 4445 7500
rect 4479 7497 4491 7531
rect 5534 7528 5540 7540
rect 5495 7500 5540 7528
rect 4433 7491 4491 7497
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 6822 7528 6828 7540
rect 6783 7500 6828 7528
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 7837 7531 7895 7537
rect 7837 7528 7849 7531
rect 7340 7500 7849 7528
rect 7340 7488 7346 7500
rect 7837 7497 7849 7500
rect 7883 7497 7895 7531
rect 7837 7491 7895 7497
rect 8938 7488 8944 7540
rect 8996 7528 9002 7540
rect 8996 7500 9996 7528
rect 8996 7488 9002 7500
rect 6914 7460 6920 7472
rect 5368 7432 6920 7460
rect 2866 7392 2872 7404
rect 2827 7364 2872 7392
rect 2866 7352 2872 7364
rect 2924 7352 2930 7404
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7361 3847 7395
rect 3789 7355 3847 7361
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7392 5135 7395
rect 5166 7392 5172 7404
rect 5123 7364 5172 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 2590 7324 2596 7336
rect 2551 7296 2596 7324
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 2682 7284 2688 7336
rect 2740 7324 2746 7336
rect 3804 7324 3832 7355
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 2740 7296 3832 7324
rect 2740 7284 2746 7296
rect 4246 7284 4252 7336
rect 4304 7324 4310 7336
rect 4893 7327 4951 7333
rect 4893 7324 4905 7327
rect 4304 7296 4905 7324
rect 4304 7284 4310 7296
rect 4893 7293 4905 7296
rect 4939 7324 4951 7327
rect 5258 7324 5264 7336
rect 4939 7296 5264 7324
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 4801 7259 4859 7265
rect 4801 7225 4813 7259
rect 4847 7256 4859 7259
rect 5368 7256 5396 7432
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 8754 7460 8760 7472
rect 7116 7432 8760 7460
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 6089 7395 6147 7401
rect 6089 7392 6101 7395
rect 5500 7364 6101 7392
rect 5500 7352 5506 7364
rect 6089 7361 6101 7364
rect 6135 7361 6147 7395
rect 6089 7355 6147 7361
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 7116 7324 7144 7432
rect 8754 7420 8760 7432
rect 8812 7420 8818 7472
rect 9968 7460 9996 7500
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 10689 7531 10747 7537
rect 10689 7528 10701 7531
rect 10284 7500 10701 7528
rect 10284 7488 10290 7500
rect 10689 7497 10701 7500
rect 10735 7497 10747 7531
rect 10689 7491 10747 7497
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 12066 7528 12072 7540
rect 11112 7500 12072 7528
rect 11112 7488 11118 7500
rect 12066 7488 12072 7500
rect 12124 7528 12130 7540
rect 13262 7528 13268 7540
rect 12124 7500 13268 7528
rect 12124 7488 12130 7500
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 13446 7528 13452 7540
rect 13407 7500 13452 7528
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 13538 7488 13544 7540
rect 13596 7528 13602 7540
rect 15657 7531 15715 7537
rect 13596 7500 14136 7528
rect 13596 7488 13602 7500
rect 10318 7460 10324 7472
rect 9968 7432 10324 7460
rect 10318 7420 10324 7432
rect 10376 7460 10382 7472
rect 10413 7463 10471 7469
rect 10413 7460 10425 7463
rect 10376 7432 10425 7460
rect 10376 7420 10382 7432
rect 10413 7429 10425 7432
rect 10459 7429 10471 7463
rect 10413 7423 10471 7429
rect 10594 7420 10600 7472
rect 10652 7460 10658 7472
rect 10652 7432 11468 7460
rect 10652 7420 10658 7432
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 7248 7364 7389 7392
rect 7248 7352 7254 7364
rect 7377 7361 7389 7364
rect 7423 7392 7435 7395
rect 8389 7395 8447 7401
rect 8389 7392 8401 7395
rect 7423 7364 8401 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 8389 7361 8401 7364
rect 8435 7361 8447 7395
rect 9030 7392 9036 7404
rect 8991 7364 9036 7392
rect 8389 7355 8447 7361
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 10134 7352 10140 7404
rect 10192 7392 10198 7404
rect 11146 7392 11152 7404
rect 10192 7364 11152 7392
rect 10192 7352 10198 7364
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 11241 7395 11299 7401
rect 11241 7361 11253 7395
rect 11287 7361 11299 7395
rect 11440 7392 11468 7432
rect 11514 7420 11520 7472
rect 11572 7460 11578 7472
rect 11572 7432 13952 7460
rect 11572 7420 11578 7432
rect 13081 7395 13139 7401
rect 11440 7364 11652 7392
rect 11241 7355 11299 7361
rect 8110 7324 8116 7336
rect 5951 7296 7144 7324
rect 7208 7296 8116 7324
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 4847 7228 5396 7256
rect 4847 7225 4859 7228
rect 4801 7219 4859 7225
rect 5442 7216 5448 7268
rect 5500 7256 5506 7268
rect 7208 7265 7236 7296
rect 8110 7284 8116 7296
rect 8168 7284 8174 7336
rect 8205 7327 8263 7333
rect 8205 7293 8217 7327
rect 8251 7324 8263 7327
rect 9122 7324 9128 7336
rect 8251 7296 9128 7324
rect 8251 7293 8263 7296
rect 8205 7287 8263 7293
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 9300 7327 9358 7333
rect 9300 7293 9312 7327
rect 9346 7324 9358 7327
rect 10594 7324 10600 7336
rect 9346 7296 10600 7324
rect 9346 7293 9358 7296
rect 9300 7287 9358 7293
rect 10594 7284 10600 7296
rect 10652 7324 10658 7336
rect 10962 7324 10968 7336
rect 10652 7296 10968 7324
rect 10652 7284 10658 7296
rect 10962 7284 10968 7296
rect 11020 7324 11026 7336
rect 11256 7324 11284 7355
rect 11020 7296 11284 7324
rect 11624 7324 11652 7364
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13354 7392 13360 7404
rect 13127 7364 13360 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 13924 7401 13952 7432
rect 14108 7401 14136 7500
rect 15657 7497 15669 7531
rect 15703 7528 15715 7531
rect 16298 7528 16304 7540
rect 15703 7500 16304 7528
rect 15703 7497 15715 7500
rect 15657 7491 15715 7497
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 18141 7531 18199 7537
rect 18141 7497 18153 7531
rect 18187 7528 18199 7531
rect 18506 7528 18512 7540
rect 18187 7500 18512 7528
rect 18187 7497 18199 7500
rect 18141 7491 18199 7497
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 18966 7488 18972 7540
rect 19024 7528 19030 7540
rect 19153 7531 19211 7537
rect 19153 7528 19165 7531
rect 19024 7500 19165 7528
rect 19024 7488 19030 7500
rect 19153 7497 19165 7500
rect 19199 7497 19211 7531
rect 19153 7491 19211 7497
rect 15010 7420 15016 7472
rect 15068 7460 15074 7472
rect 20530 7460 20536 7472
rect 15068 7432 20536 7460
rect 15068 7420 15074 7432
rect 20530 7420 20536 7432
rect 20588 7420 20594 7472
rect 13909 7395 13967 7401
rect 13909 7361 13921 7395
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7392 14151 7395
rect 14826 7392 14832 7404
rect 14139 7364 14832 7392
rect 14139 7361 14151 7364
rect 14093 7355 14151 7361
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7392 15531 7395
rect 15562 7392 15568 7404
rect 15519 7364 15568 7392
rect 15519 7361 15531 7364
rect 15473 7355 15531 7361
rect 15562 7352 15568 7364
rect 15620 7392 15626 7404
rect 16022 7392 16028 7404
rect 15620 7364 16028 7392
rect 15620 7352 15626 7364
rect 16022 7352 16028 7364
rect 16080 7352 16086 7404
rect 16390 7392 16396 7404
rect 16351 7364 16396 7392
rect 16390 7352 16396 7364
rect 16448 7352 16454 7404
rect 17310 7392 17316 7404
rect 17271 7364 17316 7392
rect 17310 7352 17316 7364
rect 17368 7352 17374 7404
rect 17497 7395 17555 7401
rect 17497 7361 17509 7395
rect 17543 7392 17555 7395
rect 17862 7392 17868 7404
rect 17543 7364 17868 7392
rect 17543 7361 17555 7364
rect 17497 7355 17555 7361
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 18693 7395 18751 7401
rect 18693 7392 18705 7395
rect 18012 7364 18705 7392
rect 18012 7352 18018 7364
rect 18693 7361 18705 7364
rect 18739 7392 18751 7395
rect 19242 7392 19248 7404
rect 18739 7364 19248 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 19242 7352 19248 7364
rect 19300 7392 19306 7404
rect 19705 7395 19763 7401
rect 19705 7392 19717 7395
rect 19300 7364 19717 7392
rect 19300 7352 19306 7364
rect 19705 7361 19717 7364
rect 19751 7361 19763 7395
rect 20622 7392 20628 7404
rect 19705 7355 19763 7361
rect 19812 7364 20628 7392
rect 13817 7327 13875 7333
rect 13817 7324 13829 7327
rect 11624 7296 13829 7324
rect 11020 7284 11026 7296
rect 13817 7293 13829 7296
rect 13863 7293 13875 7327
rect 13817 7287 13875 7293
rect 14550 7284 14556 7336
rect 14608 7324 14614 7336
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 14608 7296 14657 7324
rect 14608 7284 14614 7296
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 15197 7327 15255 7333
rect 15197 7324 15209 7327
rect 14645 7287 14703 7293
rect 14752 7296 15209 7324
rect 7193 7259 7251 7265
rect 7193 7256 7205 7259
rect 5500 7228 7205 7256
rect 5500 7216 5506 7228
rect 7193 7225 7205 7228
rect 7239 7225 7251 7259
rect 7193 7219 7251 7225
rect 7285 7259 7343 7265
rect 7285 7225 7297 7259
rect 7331 7256 7343 7259
rect 12618 7256 12624 7268
rect 7331 7228 12624 7256
rect 7331 7225 7343 7228
rect 7285 7219 7343 7225
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 13446 7216 13452 7268
rect 13504 7256 13510 7268
rect 14752 7256 14780 7296
rect 15197 7293 15209 7296
rect 15243 7293 15255 7327
rect 15197 7287 15255 7293
rect 15286 7284 15292 7336
rect 15344 7324 15350 7336
rect 16209 7327 16267 7333
rect 16209 7324 16221 7327
rect 15344 7296 16221 7324
rect 15344 7284 15350 7296
rect 16209 7293 16221 7296
rect 16255 7293 16267 7327
rect 16209 7287 16267 7293
rect 16482 7284 16488 7336
rect 16540 7324 16546 7336
rect 16540 7296 19380 7324
rect 16540 7284 16546 7296
rect 16301 7259 16359 7265
rect 16301 7256 16313 7259
rect 13504 7228 14780 7256
rect 14844 7228 16313 7256
rect 13504 7216 13510 7228
rect 2685 7191 2743 7197
rect 2685 7157 2697 7191
rect 2731 7188 2743 7191
rect 3237 7191 3295 7197
rect 3237 7188 3249 7191
rect 2731 7160 3249 7188
rect 2731 7157 2743 7160
rect 2685 7151 2743 7157
rect 3237 7157 3249 7160
rect 3283 7157 3295 7191
rect 3602 7188 3608 7200
rect 3563 7160 3608 7188
rect 3237 7151 3295 7157
rect 3602 7148 3608 7160
rect 3660 7148 3666 7200
rect 3697 7191 3755 7197
rect 3697 7157 3709 7191
rect 3743 7188 3755 7191
rect 4706 7188 4712 7200
rect 3743 7160 4712 7188
rect 3743 7157 3755 7160
rect 3697 7151 3755 7157
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 5994 7188 6000 7200
rect 5955 7160 6000 7188
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 7466 7148 7472 7200
rect 7524 7188 7530 7200
rect 8297 7191 8355 7197
rect 8297 7188 8309 7191
rect 7524 7160 8309 7188
rect 7524 7148 7530 7160
rect 8297 7157 8309 7160
rect 8343 7157 8355 7191
rect 8297 7151 8355 7157
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 10410 7188 10416 7200
rect 9732 7160 10416 7188
rect 9732 7148 9738 7160
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 11054 7188 11060 7200
rect 11015 7160 11060 7188
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11149 7191 11207 7197
rect 11149 7157 11161 7191
rect 11195 7188 11207 7191
rect 11882 7188 11888 7200
rect 11195 7160 11888 7188
rect 11195 7157 11207 7160
rect 11149 7151 11207 7157
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12802 7188 12808 7200
rect 12492 7160 12537 7188
rect 12763 7160 12808 7188
rect 12492 7148 12498 7160
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 12897 7191 12955 7197
rect 12897 7157 12909 7191
rect 12943 7188 12955 7191
rect 13170 7188 13176 7200
rect 12943 7160 13176 7188
rect 12943 7157 12955 7160
rect 12897 7151 12955 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 14844 7197 14872 7228
rect 16301 7225 16313 7228
rect 16347 7225 16359 7259
rect 18601 7259 18659 7265
rect 18601 7256 18613 7259
rect 16301 7219 16359 7225
rect 16868 7228 18613 7256
rect 14461 7191 14519 7197
rect 14461 7188 14473 7191
rect 14424 7160 14473 7188
rect 14424 7148 14430 7160
rect 14461 7157 14473 7160
rect 14507 7157 14519 7191
rect 14461 7151 14519 7157
rect 14829 7191 14887 7197
rect 14829 7157 14841 7191
rect 14875 7157 14887 7191
rect 14829 7151 14887 7157
rect 15289 7191 15347 7197
rect 15289 7157 15301 7191
rect 15335 7188 15347 7191
rect 15657 7191 15715 7197
rect 15657 7188 15669 7191
rect 15335 7160 15669 7188
rect 15335 7157 15347 7160
rect 15289 7151 15347 7157
rect 15657 7157 15669 7160
rect 15703 7157 15715 7191
rect 15657 7151 15715 7157
rect 15841 7191 15899 7197
rect 15841 7157 15853 7191
rect 15887 7188 15899 7191
rect 16206 7188 16212 7200
rect 15887 7160 16212 7188
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16868 7197 16896 7228
rect 18601 7225 18613 7228
rect 18647 7225 18659 7259
rect 19352 7256 19380 7296
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 19812 7324 19840 7364
rect 20622 7352 20628 7364
rect 20680 7392 20686 7404
rect 20717 7395 20775 7401
rect 20717 7392 20729 7395
rect 20680 7364 20729 7392
rect 20680 7352 20686 7364
rect 20717 7361 20729 7364
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 19484 7296 19840 7324
rect 19484 7284 19490 7296
rect 19886 7284 19892 7336
rect 19944 7324 19950 7336
rect 19944 7296 20668 7324
rect 19944 7284 19950 7296
rect 20254 7256 20260 7268
rect 19352 7228 20260 7256
rect 18601 7219 18659 7225
rect 20254 7216 20260 7228
rect 20312 7256 20318 7268
rect 20640 7265 20668 7296
rect 20533 7259 20591 7265
rect 20533 7256 20545 7259
rect 20312 7228 20545 7256
rect 20312 7216 20318 7228
rect 20533 7225 20545 7228
rect 20579 7225 20591 7259
rect 20533 7219 20591 7225
rect 20625 7259 20683 7265
rect 20625 7225 20637 7259
rect 20671 7225 20683 7259
rect 20625 7219 20683 7225
rect 16853 7191 16911 7197
rect 16853 7157 16865 7191
rect 16899 7157 16911 7191
rect 17218 7188 17224 7200
rect 17179 7160 17224 7188
rect 16853 7151 16911 7157
rect 17218 7148 17224 7160
rect 17276 7148 17282 7200
rect 18506 7188 18512 7200
rect 18467 7160 18512 7188
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 19518 7188 19524 7200
rect 19479 7160 19524 7188
rect 19518 7148 19524 7160
rect 19576 7148 19582 7200
rect 19610 7148 19616 7200
rect 19668 7188 19674 7200
rect 19668 7160 19713 7188
rect 19668 7148 19674 7160
rect 19886 7148 19892 7200
rect 19944 7188 19950 7200
rect 20165 7191 20223 7197
rect 20165 7188 20177 7191
rect 19944 7160 20177 7188
rect 19944 7148 19950 7160
rect 20165 7157 20177 7160
rect 20211 7157 20223 7191
rect 20165 7151 20223 7157
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 2038 6984 2044 6996
rect 1999 6956 2044 6984
rect 2038 6944 2044 6956
rect 2096 6944 2102 6996
rect 2958 6944 2964 6996
rect 3016 6984 3022 6996
rect 3016 6956 3556 6984
rect 3016 6944 3022 6956
rect 2409 6919 2467 6925
rect 2409 6885 2421 6919
rect 2455 6916 2467 6919
rect 3053 6919 3111 6925
rect 3053 6916 3065 6919
rect 2455 6888 3065 6916
rect 2455 6885 2467 6888
rect 2409 6879 2467 6885
rect 3053 6885 3065 6888
rect 3099 6885 3111 6919
rect 3528 6916 3556 6956
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 4065 6987 4123 6993
rect 4065 6984 4077 6987
rect 3660 6956 4077 6984
rect 3660 6944 3666 6956
rect 4065 6953 4077 6956
rect 4111 6953 4123 6987
rect 4065 6947 4123 6953
rect 4525 6987 4583 6993
rect 4525 6953 4537 6987
rect 4571 6984 4583 6987
rect 4890 6984 4896 6996
rect 4571 6956 4896 6984
rect 4571 6953 4583 6956
rect 4525 6947 4583 6953
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 5629 6987 5687 6993
rect 5629 6953 5641 6987
rect 5675 6984 5687 6987
rect 5902 6984 5908 6996
rect 5675 6956 5908 6984
rect 5675 6953 5687 6956
rect 5629 6947 5687 6953
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7282 6984 7288 6996
rect 6972 6956 7288 6984
rect 6972 6944 6978 6956
rect 7282 6944 7288 6956
rect 7340 6944 7346 6996
rect 9674 6984 9680 6996
rect 9635 6956 9680 6984
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 13173 6987 13231 6993
rect 13173 6984 13185 6987
rect 12860 6956 13185 6984
rect 12860 6944 12866 6956
rect 13173 6953 13185 6956
rect 13219 6953 13231 6987
rect 13173 6947 13231 6953
rect 13262 6944 13268 6996
rect 13320 6984 13326 6996
rect 15286 6984 15292 6996
rect 13320 6956 14412 6984
rect 15247 6956 15292 6984
rect 13320 6944 13326 6956
rect 3528 6888 3924 6916
rect 3053 6879 3111 6885
rect 3896 6848 3924 6888
rect 3970 6876 3976 6928
rect 4028 6916 4034 6928
rect 7098 6916 7104 6928
rect 4028 6888 6776 6916
rect 7059 6888 7104 6916
rect 4028 6876 4034 6888
rect 4433 6851 4491 6857
rect 4433 6848 4445 6851
rect 3896 6820 4445 6848
rect 4433 6817 4445 6820
rect 4479 6848 4491 6851
rect 5442 6848 5448 6860
rect 4479 6820 5448 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 5721 6851 5779 6857
rect 5721 6817 5733 6851
rect 5767 6848 5779 6851
rect 6362 6848 6368 6860
rect 5767 6820 6368 6848
rect 5767 6817 5779 6820
rect 5721 6811 5779 6817
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 6641 6851 6699 6857
rect 6641 6817 6653 6851
rect 6687 6817 6699 6851
rect 6748 6848 6776 6888
rect 7098 6876 7104 6888
rect 7156 6876 7162 6928
rect 7558 6876 7564 6928
rect 7616 6916 7622 6928
rect 8113 6919 8171 6925
rect 8113 6916 8125 6919
rect 7616 6888 8125 6916
rect 7616 6876 7622 6888
rect 8113 6885 8125 6888
rect 8159 6916 8171 6919
rect 11606 6916 11612 6928
rect 8159 6888 11612 6916
rect 8159 6885 8171 6888
rect 8113 6879 8171 6885
rect 11606 6876 11612 6888
rect 11664 6876 11670 6928
rect 11974 6916 11980 6928
rect 11716 6888 11980 6916
rect 7193 6851 7251 6857
rect 7193 6848 7205 6851
rect 6748 6820 7205 6848
rect 6641 6811 6699 6817
rect 7193 6817 7205 6820
rect 7239 6817 7251 6851
rect 7193 6811 7251 6817
rect 2498 6780 2504 6792
rect 2459 6752 2504 6780
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 2590 6740 2596 6792
rect 2648 6780 2654 6792
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 2648 6752 4629 6780
rect 2648 6740 2654 6752
rect 4617 6749 4629 6752
rect 4663 6749 4675 6783
rect 5902 6780 5908 6792
rect 5863 6752 5908 6780
rect 4617 6743 4675 6749
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 6656 6780 6684 6811
rect 8018 6808 8024 6860
rect 8076 6848 8082 6860
rect 8205 6851 8263 6857
rect 8205 6848 8217 6851
rect 8076 6820 8217 6848
rect 8076 6808 8082 6820
rect 8205 6817 8217 6820
rect 8251 6817 8263 6851
rect 10042 6848 10048 6860
rect 10003 6820 10048 6848
rect 8205 6811 8263 6817
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11716 6848 11744 6888
rect 11974 6876 11980 6888
rect 12032 6876 12038 6928
rect 12158 6876 12164 6928
rect 12216 6916 12222 6928
rect 14277 6919 14335 6925
rect 14277 6916 14289 6919
rect 12216 6888 14289 6916
rect 12216 6876 12222 6888
rect 14277 6885 14289 6888
rect 14323 6885 14335 6919
rect 14384 6916 14412 6956
rect 15286 6944 15292 6956
rect 15344 6944 15350 6996
rect 15657 6987 15715 6993
rect 15657 6953 15669 6987
rect 15703 6984 15715 6987
rect 15746 6984 15752 6996
rect 15703 6956 15752 6984
rect 15703 6953 15715 6956
rect 15657 6947 15715 6953
rect 15746 6944 15752 6956
rect 15804 6944 15810 6996
rect 16390 6944 16396 6996
rect 16448 6984 16454 6996
rect 17313 6987 17371 6993
rect 16448 6956 16988 6984
rect 16448 6944 16454 6956
rect 16669 6919 16727 6925
rect 16669 6916 16681 6919
rect 14384 6888 16681 6916
rect 14277 6879 14335 6885
rect 16669 6885 16681 6888
rect 16715 6885 16727 6919
rect 16669 6879 16727 6885
rect 16758 6876 16764 6928
rect 16816 6916 16822 6928
rect 16960 6916 16988 6956
rect 17313 6953 17325 6987
rect 17359 6984 17371 6987
rect 17402 6984 17408 6996
rect 17359 6956 17408 6984
rect 17359 6953 17371 6956
rect 17313 6947 17371 6953
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 17678 6944 17684 6996
rect 17736 6984 17742 6996
rect 17862 6984 17868 6996
rect 17736 6956 17868 6984
rect 17736 6944 17742 6956
rect 17862 6944 17868 6956
rect 17920 6984 17926 6996
rect 18141 6987 18199 6993
rect 18141 6984 18153 6987
rect 17920 6956 18153 6984
rect 17920 6944 17926 6956
rect 18141 6953 18153 6956
rect 18187 6953 18199 6987
rect 18141 6947 18199 6953
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 18785 6987 18843 6993
rect 18785 6984 18797 6987
rect 18564 6956 18797 6984
rect 18564 6944 18570 6956
rect 18785 6953 18797 6956
rect 18831 6953 18843 6987
rect 19426 6984 19432 6996
rect 18785 6947 18843 6953
rect 19076 6956 19432 6984
rect 18598 6916 18604 6928
rect 16816 6888 16861 6916
rect 16960 6888 18604 6916
rect 16816 6876 16822 6888
rect 18598 6876 18604 6888
rect 18656 6876 18662 6928
rect 11112 6820 11744 6848
rect 11784 6851 11842 6857
rect 11112 6808 11118 6820
rect 11784 6817 11796 6851
rect 11830 6848 11842 6851
rect 13354 6848 13360 6860
rect 11830 6820 13360 6848
rect 11830 6817 11842 6820
rect 11784 6811 11842 6817
rect 13354 6808 13360 6820
rect 13412 6808 13418 6860
rect 14458 6808 14464 6860
rect 14516 6848 14522 6860
rect 17497 6851 17555 6857
rect 17497 6848 17509 6851
rect 14516 6820 17509 6848
rect 14516 6808 14522 6820
rect 17497 6817 17509 6820
rect 17543 6817 17555 6851
rect 17497 6811 17555 6817
rect 18506 6808 18512 6860
rect 18564 6848 18570 6860
rect 18782 6848 18788 6860
rect 18564 6820 18788 6848
rect 18564 6808 18570 6820
rect 18782 6808 18788 6820
rect 18840 6808 18846 6860
rect 7006 6780 7012 6792
rect 6656 6752 7012 6780
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6780 7435 6783
rect 8294 6780 8300 6792
rect 7423 6752 8300 6780
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 8294 6740 8300 6752
rect 8352 6780 8358 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 8352 6752 8401 6780
rect 8352 6740 8358 6752
rect 8389 6749 8401 6752
rect 8435 6780 8447 6783
rect 9214 6780 9220 6792
rect 8435 6752 9220 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10318 6780 10324 6792
rect 10279 6752 10324 6780
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 6733 6715 6791 6721
rect 5184 6684 6684 6712
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 5184 6644 5212 6684
rect 4120 6616 5212 6644
rect 5261 6647 5319 6653
rect 4120 6604 4126 6616
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5442 6644 5448 6656
rect 5307 6616 5448 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 6454 6644 6460 6656
rect 5592 6616 6460 6644
rect 5592 6604 5598 6616
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 6656 6644 6684 6684
rect 6733 6681 6745 6715
rect 6779 6712 6791 6715
rect 8110 6712 8116 6724
rect 6779 6684 8116 6712
rect 6779 6681 6791 6684
rect 6733 6675 6791 6681
rect 8110 6672 8116 6684
rect 8168 6672 8174 6724
rect 8754 6672 8760 6724
rect 8812 6712 8818 6724
rect 11422 6712 11428 6724
rect 8812 6684 11428 6712
rect 8812 6672 8818 6684
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 7558 6644 7564 6656
rect 6656 6616 7564 6644
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 7742 6644 7748 6656
rect 7703 6616 7748 6644
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 7834 6604 7840 6656
rect 7892 6644 7898 6656
rect 11054 6644 11060 6656
rect 7892 6616 11060 6644
rect 7892 6604 7898 6616
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11532 6644 11560 6743
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 14369 6783 14427 6789
rect 14369 6780 14381 6783
rect 13964 6752 14381 6780
rect 13964 6740 13970 6752
rect 14369 6749 14381 6752
rect 14415 6749 14427 6783
rect 14369 6743 14427 6749
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 14826 6780 14832 6792
rect 14599 6752 14832 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 14826 6740 14832 6752
rect 14884 6740 14890 6792
rect 15654 6740 15660 6792
rect 15712 6780 15718 6792
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 15712 6752 15761 6780
rect 15712 6740 15718 6752
rect 15749 6749 15761 6752
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15933 6783 15991 6789
rect 15933 6749 15945 6783
rect 15979 6780 15991 6783
rect 16022 6780 16028 6792
rect 15979 6752 16028 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 16850 6780 16856 6792
rect 16811 6752 16856 6780
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 16942 6740 16948 6792
rect 17000 6780 17006 6792
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 17000 6752 18245 6780
rect 17000 6740 17006 6752
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 19076 6780 19104 6956
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 19797 6987 19855 6993
rect 19797 6984 19809 6987
rect 19576 6956 19809 6984
rect 19576 6944 19582 6956
rect 19797 6953 19809 6956
rect 19843 6953 19855 6987
rect 19797 6947 19855 6953
rect 19153 6919 19211 6925
rect 19153 6885 19165 6919
rect 19199 6916 19211 6919
rect 20898 6916 20904 6928
rect 19199 6888 20904 6916
rect 19199 6885 19211 6888
rect 19153 6879 19211 6885
rect 20898 6876 20904 6888
rect 20956 6876 20962 6928
rect 19245 6851 19303 6857
rect 19245 6817 19257 6851
rect 19291 6848 19303 6851
rect 19886 6848 19892 6860
rect 19291 6820 19892 6848
rect 19291 6817 19303 6820
rect 19245 6811 19303 6817
rect 19886 6808 19892 6820
rect 19944 6808 19950 6860
rect 20162 6848 20168 6860
rect 20123 6820 20168 6848
rect 20162 6808 20168 6820
rect 20220 6808 20226 6860
rect 18325 6743 18383 6749
rect 18800 6752 19104 6780
rect 12526 6672 12532 6724
rect 12584 6712 12590 6724
rect 16758 6712 16764 6724
rect 12584 6684 16764 6712
rect 12584 6672 12590 6684
rect 16758 6672 16764 6684
rect 16816 6672 16822 6724
rect 16868 6712 16896 6740
rect 18340 6712 18368 6743
rect 18800 6724 18828 6752
rect 19150 6740 19156 6792
rect 19208 6780 19214 6792
rect 19337 6783 19395 6789
rect 19337 6780 19349 6783
rect 19208 6752 19349 6780
rect 19208 6740 19214 6752
rect 19337 6749 19349 6752
rect 19383 6749 19395 6783
rect 20254 6780 20260 6792
rect 20215 6752 20260 6780
rect 19337 6743 19395 6749
rect 18782 6712 18788 6724
rect 16868 6684 18788 6712
rect 18782 6672 18788 6684
rect 18840 6672 18846 6724
rect 19352 6712 19380 6743
rect 20254 6740 20260 6752
rect 20312 6740 20318 6792
rect 20349 6783 20407 6789
rect 20349 6749 20361 6783
rect 20395 6749 20407 6783
rect 20349 6743 20407 6749
rect 20364 6712 20392 6743
rect 19352 6684 20392 6712
rect 12250 6644 12256 6656
rect 11532 6616 12256 6644
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 12860 6616 12909 6644
rect 12860 6604 12866 6616
rect 12897 6613 12909 6616
rect 12943 6613 12955 6647
rect 12897 6607 12955 6613
rect 13909 6647 13967 6653
rect 13909 6613 13921 6647
rect 13955 6644 13967 6647
rect 14642 6644 14648 6656
rect 13955 6616 14648 6644
rect 13955 6613 13967 6616
rect 13909 6607 13967 6613
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 16301 6647 16359 6653
rect 16301 6613 16313 6647
rect 16347 6644 16359 6647
rect 17218 6644 17224 6656
rect 16347 6616 17224 6644
rect 16347 6613 16359 6616
rect 16301 6607 16359 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 17773 6647 17831 6653
rect 17773 6613 17785 6647
rect 17819 6644 17831 6647
rect 19702 6644 19708 6656
rect 17819 6616 19708 6644
rect 17819 6613 17831 6616
rect 17773 6607 17831 6613
rect 19702 6604 19708 6616
rect 19760 6604 19766 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 3145 6443 3203 6449
rect 3145 6440 3157 6443
rect 2740 6412 3157 6440
rect 2740 6400 2746 6412
rect 3145 6409 3157 6412
rect 3191 6409 3203 6443
rect 3418 6440 3424 6452
rect 3379 6412 3424 6440
rect 3145 6403 3203 6409
rect 3418 6400 3424 6412
rect 3476 6400 3482 6452
rect 5534 6440 5540 6452
rect 4724 6412 5540 6440
rect 3973 6307 4031 6313
rect 3973 6273 3985 6307
rect 4019 6273 4031 6307
rect 3973 6267 4031 6273
rect 1765 6239 1823 6245
rect 1765 6205 1777 6239
rect 1811 6236 1823 6239
rect 2032 6239 2090 6245
rect 1811 6208 1992 6236
rect 1811 6205 1823 6208
rect 1765 6199 1823 6205
rect 1964 6180 1992 6208
rect 2032 6205 2044 6239
rect 2078 6236 2090 6239
rect 2590 6236 2596 6248
rect 2078 6208 2596 6236
rect 2078 6205 2090 6208
rect 2032 6199 2090 6205
rect 2590 6196 2596 6208
rect 2648 6236 2654 6248
rect 3988 6236 4016 6267
rect 4724 6245 4752 6412
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 9953 6443 10011 6449
rect 5960 6412 8524 6440
rect 5960 6400 5966 6412
rect 2648 6208 4016 6236
rect 2648 6196 2654 6208
rect 1946 6128 1952 6180
rect 2004 6128 2010 6180
rect 3326 6128 3332 6180
rect 3384 6168 3390 6180
rect 3694 6168 3700 6180
rect 3384 6140 3700 6168
rect 3384 6128 3390 6140
rect 3694 6128 3700 6140
rect 3752 6168 3758 6180
rect 3881 6171 3939 6177
rect 3881 6168 3893 6171
rect 3752 6140 3893 6168
rect 3752 6128 3758 6140
rect 3881 6137 3893 6140
rect 3927 6137 3939 6171
rect 3988 6168 4016 6208
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6205 4767 6239
rect 4709 6199 4767 6205
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 5068 6239 5126 6245
rect 4856 6208 4901 6236
rect 4856 6196 4862 6208
rect 5068 6205 5080 6239
rect 5114 6236 5126 6239
rect 5920 6236 5948 6400
rect 7116 6304 7144 6412
rect 7190 6332 7196 6384
rect 7248 6372 7254 6384
rect 8018 6372 8024 6384
rect 7248 6344 8024 6372
rect 7248 6332 7254 6344
rect 8018 6332 8024 6344
rect 8076 6332 8082 6384
rect 8202 6332 8208 6384
rect 8260 6372 8266 6384
rect 8496 6372 8524 6412
rect 9953 6409 9965 6443
rect 9999 6440 10011 6443
rect 10042 6440 10048 6452
rect 9999 6412 10048 6440
rect 9999 6409 10011 6412
rect 9953 6403 10011 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 10965 6443 11023 6449
rect 10965 6440 10977 6443
rect 10192 6412 10977 6440
rect 10192 6400 10198 6412
rect 10965 6409 10977 6412
rect 11011 6409 11023 6443
rect 10965 6403 11023 6409
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 13446 6440 13452 6452
rect 11664 6412 13452 6440
rect 11664 6400 11670 6412
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 13906 6440 13912 6452
rect 13819 6412 13912 6440
rect 13906 6400 13912 6412
rect 13964 6440 13970 6452
rect 14826 6440 14832 6452
rect 13964 6412 14832 6440
rect 13964 6400 13970 6412
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 15654 6400 15660 6452
rect 15712 6440 15718 6452
rect 16482 6440 16488 6452
rect 15712 6412 16488 6440
rect 15712 6400 15718 6412
rect 16482 6400 16488 6412
rect 16540 6400 16546 6452
rect 16666 6400 16672 6452
rect 16724 6440 16730 6452
rect 16945 6443 17003 6449
rect 16945 6440 16957 6443
rect 16724 6412 16957 6440
rect 16724 6400 16730 6412
rect 16945 6409 16957 6412
rect 16991 6409 17003 6443
rect 16945 6403 17003 6409
rect 17494 6400 17500 6452
rect 17552 6440 17558 6452
rect 18598 6440 18604 6452
rect 17552 6412 18604 6440
rect 17552 6400 17558 6412
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 19245 6443 19303 6449
rect 19245 6409 19257 6443
rect 19291 6440 19303 6443
rect 19610 6440 19616 6452
rect 19291 6412 19616 6440
rect 19291 6409 19303 6412
rect 19245 6403 19303 6409
rect 19610 6400 19616 6412
rect 19668 6400 19674 6452
rect 20254 6440 20260 6452
rect 20215 6412 20260 6440
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 10870 6372 10876 6384
rect 8260 6344 8432 6372
rect 8496 6344 10876 6372
rect 8260 6332 8266 6344
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7116 6276 7389 6304
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7742 6264 7748 6316
rect 7800 6304 7806 6316
rect 8404 6313 8432 6344
rect 10870 6332 10876 6344
rect 10928 6332 10934 6384
rect 12069 6375 12127 6381
rect 12069 6341 12081 6375
rect 12115 6372 12127 6375
rect 12342 6372 12348 6384
rect 12115 6344 12348 6372
rect 12115 6341 12127 6344
rect 12069 6335 12127 6341
rect 12342 6332 12348 6344
rect 12400 6372 12406 6384
rect 12400 6344 12572 6372
rect 12400 6332 12406 6344
rect 8297 6307 8355 6313
rect 8297 6304 8309 6307
rect 7800 6276 8309 6304
rect 7800 6264 7806 6276
rect 8297 6273 8309 6276
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 9214 6264 9220 6316
rect 9272 6304 9278 6316
rect 9401 6307 9459 6313
rect 9401 6304 9413 6307
rect 9272 6276 9413 6304
rect 9272 6264 9278 6276
rect 9401 6273 9413 6276
rect 9447 6273 9459 6307
rect 10502 6304 10508 6316
rect 9401 6267 9459 6273
rect 9600 6276 10508 6304
rect 5114 6208 5948 6236
rect 5114 6205 5126 6208
rect 5068 6199 5126 6205
rect 6822 6196 6828 6248
rect 6880 6236 6886 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 6880 6208 7297 6236
rect 6880 6196 6886 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 8110 6196 8116 6248
rect 8168 6236 8174 6248
rect 8205 6239 8263 6245
rect 8205 6236 8217 6239
rect 8168 6208 8217 6236
rect 8168 6196 8174 6208
rect 8205 6205 8217 6208
rect 8251 6205 8263 6239
rect 8205 6199 8263 6205
rect 8478 6196 8484 6248
rect 8536 6236 8542 6248
rect 9309 6239 9367 6245
rect 9309 6236 9321 6239
rect 8536 6208 9321 6236
rect 8536 6196 8542 6208
rect 9309 6205 9321 6208
rect 9355 6236 9367 6239
rect 9600 6236 9628 6276
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 10594 6264 10600 6316
rect 10652 6304 10658 6316
rect 10962 6304 10968 6316
rect 10652 6276 10968 6304
rect 10652 6264 10658 6276
rect 10962 6264 10968 6276
rect 11020 6304 11026 6316
rect 12544 6313 12572 6344
rect 14550 6332 14556 6384
rect 14608 6372 14614 6384
rect 16577 6375 16635 6381
rect 14608 6344 14780 6372
rect 14608 6332 14614 6344
rect 11517 6307 11575 6313
rect 11517 6304 11529 6307
rect 11020 6276 11529 6304
rect 11020 6264 11026 6276
rect 11517 6273 11529 6276
rect 11563 6273 11575 6307
rect 12529 6307 12587 6313
rect 11517 6267 11575 6273
rect 12268 6276 12480 6304
rect 9355 6208 9628 6236
rect 9355 6205 9367 6208
rect 9309 6199 9367 6205
rect 9674 6196 9680 6248
rect 9732 6236 9738 6248
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 9732 6208 10425 6236
rect 9732 6196 9738 6208
rect 10413 6205 10425 6208
rect 10459 6236 10471 6239
rect 12158 6236 12164 6248
rect 10459 6208 12164 6236
rect 10459 6205 10471 6208
rect 10413 6199 10471 6205
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 12268 6245 12296 6276
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6205 12311 6239
rect 12253 6199 12311 6205
rect 5534 6168 5540 6180
rect 3988 6140 5540 6168
rect 3881 6131 3939 6137
rect 5534 6128 5540 6140
rect 5592 6168 5598 6180
rect 7193 6171 7251 6177
rect 5592 6140 6224 6168
rect 5592 6128 5598 6140
rect 2774 6060 2780 6112
rect 2832 6100 2838 6112
rect 3786 6100 3792 6112
rect 2832 6072 3792 6100
rect 2832 6060 2838 6072
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 4525 6103 4583 6109
rect 4525 6069 4537 6103
rect 4571 6100 4583 6103
rect 4798 6100 4804 6112
rect 4571 6072 4804 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 6196 6109 6224 6140
rect 7193 6137 7205 6171
rect 7239 6168 7251 6171
rect 10134 6168 10140 6180
rect 7239 6140 10140 6168
rect 7239 6137 7251 6140
rect 7193 6131 7251 6137
rect 10134 6128 10140 6140
rect 10192 6128 10198 6180
rect 10321 6171 10379 6177
rect 10321 6137 10333 6171
rect 10367 6168 10379 6171
rect 11606 6168 11612 6180
rect 10367 6140 11612 6168
rect 10367 6137 10379 6140
rect 10321 6131 10379 6137
rect 6181 6103 6239 6109
rect 6181 6069 6193 6103
rect 6227 6069 6239 6103
rect 6181 6063 6239 6069
rect 6270 6060 6276 6112
rect 6328 6100 6334 6112
rect 6825 6103 6883 6109
rect 6825 6100 6837 6103
rect 6328 6072 6837 6100
rect 6328 6060 6334 6072
rect 6825 6069 6837 6072
rect 6871 6069 6883 6103
rect 6825 6063 6883 6069
rect 7742 6060 7748 6112
rect 7800 6100 7806 6112
rect 7837 6103 7895 6109
rect 7837 6100 7849 6103
rect 7800 6072 7849 6100
rect 7800 6060 7806 6072
rect 7837 6069 7849 6072
rect 7883 6069 7895 6103
rect 7837 6063 7895 6069
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 8849 6103 8907 6109
rect 8849 6100 8861 6103
rect 8628 6072 8861 6100
rect 8628 6060 8634 6072
rect 8849 6069 8861 6072
rect 8895 6069 8907 6103
rect 8849 6063 8907 6069
rect 8938 6060 8944 6112
rect 8996 6100 9002 6112
rect 9217 6103 9275 6109
rect 9217 6100 9229 6103
rect 8996 6072 9229 6100
rect 8996 6060 9002 6072
rect 9217 6069 9229 6072
rect 9263 6069 9275 6103
rect 9217 6063 9275 6069
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 10336 6100 10364 6131
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 12452 6168 12480 6276
rect 12529 6273 12541 6307
rect 12575 6273 12587 6307
rect 14642 6304 14648 6316
rect 14603 6276 14648 6304
rect 12529 6267 12587 6273
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 14752 6313 14780 6344
rect 16577 6341 16589 6375
rect 16623 6372 16635 6375
rect 16623 6344 19104 6372
rect 16623 6341 16635 6344
rect 16577 6335 16635 6341
rect 14737 6307 14795 6313
rect 14737 6273 14749 6307
rect 14783 6273 14795 6307
rect 14737 6267 14795 6273
rect 14826 6264 14832 6316
rect 14884 6304 14890 6316
rect 15749 6307 15807 6313
rect 15749 6304 15761 6307
rect 14884 6276 15761 6304
rect 14884 6264 14890 6276
rect 15749 6273 15761 6276
rect 15795 6273 15807 6307
rect 15749 6267 15807 6273
rect 15838 6264 15844 6316
rect 15896 6304 15902 6316
rect 17497 6307 17555 6313
rect 17497 6304 17509 6307
rect 15896 6276 17509 6304
rect 15896 6264 15902 6276
rect 17497 6273 17509 6276
rect 17543 6304 17555 6307
rect 18414 6304 18420 6316
rect 17543 6276 18420 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 18414 6264 18420 6276
rect 18472 6264 18478 6316
rect 18782 6304 18788 6316
rect 18743 6276 18788 6304
rect 18782 6264 18788 6276
rect 18840 6264 18846 6316
rect 19076 6304 19104 6344
rect 19150 6332 19156 6384
rect 19208 6372 19214 6384
rect 19208 6344 19840 6372
rect 19208 6332 19214 6344
rect 19518 6304 19524 6316
rect 19076 6276 19524 6304
rect 19518 6264 19524 6276
rect 19576 6264 19582 6316
rect 19702 6304 19708 6316
rect 19663 6276 19708 6304
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 19812 6313 19840 6344
rect 19797 6307 19855 6313
rect 19797 6273 19809 6307
rect 19843 6273 19855 6307
rect 19797 6267 19855 6273
rect 20622 6264 20628 6316
rect 20680 6304 20686 6316
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 20680 6276 20821 6304
rect 20680 6264 20686 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 12802 6245 12808 6248
rect 12796 6236 12808 6245
rect 12763 6208 12808 6236
rect 12796 6199 12808 6208
rect 12802 6196 12808 6199
rect 12860 6196 12866 6248
rect 15470 6196 15476 6248
rect 15528 6236 15534 6248
rect 15657 6239 15715 6245
rect 15657 6236 15669 6239
rect 15528 6208 15669 6236
rect 15528 6196 15534 6208
rect 15657 6205 15669 6208
rect 15703 6205 15715 6239
rect 15657 6199 15715 6205
rect 16298 6196 16304 6248
rect 16356 6236 16362 6248
rect 16393 6239 16451 6245
rect 16393 6236 16405 6239
rect 16356 6208 16405 6236
rect 16356 6196 16362 6208
rect 16393 6205 16405 6208
rect 16439 6205 16451 6239
rect 16393 6199 16451 6205
rect 18601 6239 18659 6245
rect 18601 6205 18613 6239
rect 18647 6236 18659 6239
rect 19886 6236 19892 6248
rect 18647 6208 19892 6236
rect 18647 6205 18659 6208
rect 18601 6199 18659 6205
rect 19886 6196 19892 6208
rect 19944 6196 19950 6248
rect 14366 6168 14372 6180
rect 12452 6140 14372 6168
rect 14366 6128 14372 6140
rect 14424 6128 14430 6180
rect 14553 6171 14611 6177
rect 14553 6137 14565 6171
rect 14599 6168 14611 6171
rect 14599 6140 15240 6168
rect 14599 6137 14611 6140
rect 14553 6131 14611 6137
rect 9916 6072 10364 6100
rect 9916 6060 9922 6072
rect 10410 6060 10416 6112
rect 10468 6100 10474 6112
rect 11333 6103 11391 6109
rect 11333 6100 11345 6103
rect 10468 6072 11345 6100
rect 10468 6060 10474 6072
rect 11333 6069 11345 6072
rect 11379 6069 11391 6103
rect 11333 6063 11391 6069
rect 11425 6103 11483 6109
rect 11425 6069 11437 6103
rect 11471 6100 11483 6103
rect 11698 6100 11704 6112
rect 11471 6072 11704 6100
rect 11471 6069 11483 6072
rect 11425 6063 11483 6069
rect 11698 6060 11704 6072
rect 11756 6100 11762 6112
rect 13078 6100 13084 6112
rect 11756 6072 13084 6100
rect 11756 6060 11762 6072
rect 13078 6060 13084 6072
rect 13136 6060 13142 6112
rect 14185 6103 14243 6109
rect 14185 6069 14197 6103
rect 14231 6100 14243 6103
rect 14458 6100 14464 6112
rect 14231 6072 14464 6100
rect 14231 6069 14243 6072
rect 14185 6063 14243 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 15212 6109 15240 6140
rect 16666 6128 16672 6180
rect 16724 6168 16730 6180
rect 17405 6171 17463 6177
rect 17405 6168 17417 6171
rect 16724 6140 17417 6168
rect 16724 6128 16730 6140
rect 17405 6137 17417 6140
rect 17451 6137 17463 6171
rect 19613 6171 19671 6177
rect 19613 6168 19625 6171
rect 17405 6131 17463 6137
rect 18248 6140 19625 6168
rect 15197 6103 15255 6109
rect 15197 6069 15209 6103
rect 15243 6069 15255 6103
rect 15562 6100 15568 6112
rect 15523 6072 15568 6100
rect 15197 6063 15255 6069
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 17310 6100 17316 6112
rect 17271 6072 17316 6100
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 18248 6109 18276 6140
rect 19613 6137 19625 6140
rect 19659 6137 19671 6171
rect 19613 6131 19671 6137
rect 20530 6128 20536 6180
rect 20588 6168 20594 6180
rect 20625 6171 20683 6177
rect 20625 6168 20637 6171
rect 20588 6140 20637 6168
rect 20588 6128 20594 6140
rect 20625 6137 20637 6140
rect 20671 6137 20683 6171
rect 20625 6131 20683 6137
rect 18233 6103 18291 6109
rect 18233 6069 18245 6103
rect 18279 6069 18291 6103
rect 18233 6063 18291 6069
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 18782 6100 18788 6112
rect 18739 6072 18788 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 18782 6060 18788 6072
rect 18840 6060 18846 6112
rect 20346 6060 20352 6112
rect 20404 6100 20410 6112
rect 20717 6103 20775 6109
rect 20717 6100 20729 6103
rect 20404 6072 20729 6100
rect 20404 6060 20410 6072
rect 20717 6069 20729 6072
rect 20763 6100 20775 6103
rect 20898 6100 20904 6112
rect 20763 6072 20904 6100
rect 20763 6069 20775 6072
rect 20717 6063 20775 6069
rect 20898 6060 20904 6072
rect 20956 6060 20962 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3697 5899 3755 5905
rect 3697 5896 3709 5899
rect 2924 5868 3709 5896
rect 2924 5856 2930 5868
rect 3697 5865 3709 5868
rect 3743 5896 3755 5899
rect 3786 5896 3792 5908
rect 3743 5868 3792 5896
rect 3743 5865 3755 5868
rect 3697 5859 3755 5865
rect 3786 5856 3792 5868
rect 3844 5856 3850 5908
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 4985 5899 5043 5905
rect 4985 5896 4997 5899
rect 4764 5868 4997 5896
rect 4764 5856 4770 5868
rect 4985 5865 4997 5868
rect 5031 5865 5043 5899
rect 5442 5896 5448 5908
rect 5403 5868 5448 5896
rect 4985 5859 5043 5865
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 7800 5868 8677 5896
rect 7800 5856 7806 5868
rect 8665 5865 8677 5868
rect 8711 5865 8723 5899
rect 8665 5859 8723 5865
rect 8772 5868 10916 5896
rect 2584 5831 2642 5837
rect 2584 5797 2596 5831
rect 2630 5828 2642 5831
rect 2682 5828 2688 5840
rect 2630 5800 2688 5828
rect 2630 5797 2642 5800
rect 2584 5791 2642 5797
rect 2682 5788 2688 5800
rect 2740 5788 2746 5840
rect 5353 5831 5411 5837
rect 5353 5797 5365 5831
rect 5399 5828 5411 5831
rect 6270 5828 6276 5840
rect 5399 5800 6276 5828
rect 5399 5797 5411 5800
rect 5353 5791 5411 5797
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 6362 5788 6368 5840
rect 6420 5828 6426 5840
rect 6908 5831 6966 5837
rect 6420 5800 6776 5828
rect 6420 5788 6426 5800
rect 4798 5720 4804 5772
rect 4856 5760 4862 5772
rect 6641 5763 6699 5769
rect 6641 5760 6653 5763
rect 4856 5732 6653 5760
rect 4856 5720 4862 5732
rect 6641 5729 6653 5732
rect 6687 5729 6699 5763
rect 6748 5760 6776 5800
rect 6908 5797 6920 5831
rect 6954 5828 6966 5831
rect 8294 5828 8300 5840
rect 6954 5800 8300 5828
rect 6954 5797 6966 5800
rect 6908 5791 6966 5797
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 8772 5760 8800 5868
rect 10778 5828 10784 5840
rect 6748 5732 8800 5760
rect 8864 5800 10784 5828
rect 6641 5723 6699 5729
rect 1946 5652 1952 5704
rect 2004 5692 2010 5704
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 2004 5664 2329 5692
rect 2004 5652 2010 5664
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 5534 5692 5540 5704
rect 5495 5664 5540 5692
rect 2317 5655 2375 5661
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8757 5695 8815 5701
rect 8757 5692 8769 5695
rect 8352 5664 8769 5692
rect 8352 5652 8358 5664
rect 8757 5661 8769 5664
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 8864 5624 8892 5800
rect 10778 5788 10784 5800
rect 10836 5788 10842 5840
rect 10888 5828 10916 5868
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 11020 5868 11069 5896
rect 11020 5856 11026 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 13081 5899 13139 5905
rect 12492 5868 12537 5896
rect 12492 5856 12498 5868
rect 13081 5865 13093 5899
rect 13127 5896 13139 5899
rect 15562 5896 15568 5908
rect 13127 5868 15568 5896
rect 13127 5865 13139 5868
rect 13081 5859 13139 5865
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 18414 5856 18420 5908
rect 18472 5896 18478 5908
rect 19061 5899 19119 5905
rect 19061 5896 19073 5899
rect 18472 5868 19073 5896
rect 18472 5856 18478 5868
rect 19061 5865 19073 5868
rect 19107 5865 19119 5899
rect 19061 5859 19119 5865
rect 19797 5899 19855 5905
rect 19797 5865 19809 5899
rect 19843 5896 19855 5899
rect 20162 5896 20168 5908
rect 19843 5868 20168 5896
rect 19843 5865 19855 5868
rect 19797 5859 19855 5865
rect 20162 5856 20168 5868
rect 20220 5856 20226 5908
rect 12986 5828 12992 5840
rect 10888 5800 12992 5828
rect 12986 5788 12992 5800
rect 13044 5788 13050 5840
rect 13808 5831 13866 5837
rect 13808 5797 13820 5831
rect 13854 5828 13866 5831
rect 13906 5828 13912 5840
rect 13854 5800 13912 5828
rect 13854 5797 13866 5800
rect 13808 5791 13866 5797
rect 13906 5788 13912 5800
rect 13964 5788 13970 5840
rect 14642 5788 14648 5840
rect 14700 5828 14706 5840
rect 14700 5800 16620 5828
rect 14700 5788 14706 5800
rect 9933 5763 9991 5769
rect 9933 5760 9945 5763
rect 8956 5732 9945 5760
rect 8956 5704 8984 5732
rect 9933 5729 9945 5732
rect 9979 5729 9991 5763
rect 9933 5723 9991 5729
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 13538 5760 13544 5772
rect 12400 5732 13544 5760
rect 12400 5720 12406 5732
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 15470 5760 15476 5772
rect 15431 5732 15476 5760
rect 15470 5720 15476 5732
rect 15528 5760 15534 5772
rect 16040 5769 16068 5800
rect 16298 5769 16304 5772
rect 15841 5763 15899 5769
rect 15841 5760 15853 5763
rect 15528 5732 15853 5760
rect 15528 5720 15534 5732
rect 15841 5729 15853 5732
rect 15887 5729 15899 5763
rect 15841 5723 15899 5729
rect 16025 5763 16083 5769
rect 16025 5729 16037 5763
rect 16071 5729 16083 5763
rect 16292 5760 16304 5769
rect 16259 5732 16304 5760
rect 16025 5723 16083 5729
rect 16292 5723 16304 5732
rect 16298 5720 16304 5723
rect 16356 5720 16362 5772
rect 16592 5760 16620 5800
rect 17218 5788 17224 5840
rect 17276 5828 17282 5840
rect 18874 5828 18880 5840
rect 17276 5800 18880 5828
rect 17276 5788 17282 5800
rect 18874 5788 18880 5800
rect 18932 5788 18938 5840
rect 17126 5760 17132 5772
rect 16592 5732 17132 5760
rect 17126 5720 17132 5732
rect 17184 5760 17190 5772
rect 17589 5763 17647 5769
rect 17184 5732 17448 5760
rect 17184 5720 17190 5732
rect 17420 5704 17448 5732
rect 17589 5729 17601 5763
rect 17635 5760 17647 5763
rect 17937 5763 17995 5769
rect 17937 5760 17949 5763
rect 17635 5732 17949 5760
rect 17635 5729 17647 5732
rect 17589 5723 17647 5729
rect 17937 5729 17949 5732
rect 17983 5729 17995 5763
rect 20162 5760 20168 5772
rect 20123 5732 20168 5760
rect 17937 5723 17995 5729
rect 20162 5720 20168 5732
rect 20220 5720 20226 5772
rect 8938 5652 8944 5704
rect 8996 5692 9002 5704
rect 9677 5695 9735 5701
rect 8996 5664 9089 5692
rect 8996 5652 9002 5664
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 12526 5692 12532 5704
rect 12487 5664 12532 5692
rect 9677 5655 9735 5661
rect 7576 5596 8892 5624
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 7006 5556 7012 5568
rect 4120 5528 7012 5556
rect 4120 5516 4126 5528
rect 7006 5516 7012 5528
rect 7064 5556 7070 5568
rect 7576 5556 7604 5596
rect 9030 5584 9036 5636
rect 9088 5624 9094 5636
rect 9692 5624 9720 5655
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 12713 5695 12771 5701
rect 12713 5661 12725 5695
rect 12759 5692 12771 5695
rect 12802 5692 12808 5704
rect 12759 5664 12808 5692
rect 12759 5661 12771 5664
rect 12713 5655 12771 5661
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 17402 5652 17408 5704
rect 17460 5692 17466 5704
rect 17681 5695 17739 5701
rect 17681 5692 17693 5695
rect 17460 5664 17693 5692
rect 17460 5652 17466 5664
rect 17681 5661 17693 5664
rect 17727 5661 17739 5695
rect 17681 5655 17739 5661
rect 18782 5652 18788 5704
rect 18840 5692 18846 5704
rect 19337 5695 19395 5701
rect 19337 5692 19349 5695
rect 18840 5664 19349 5692
rect 18840 5652 18846 5664
rect 19337 5661 19349 5664
rect 19383 5661 19395 5695
rect 19337 5655 19395 5661
rect 19794 5652 19800 5704
rect 19852 5692 19858 5704
rect 20257 5695 20315 5701
rect 20257 5692 20269 5695
rect 19852 5664 20269 5692
rect 19852 5652 19858 5664
rect 20257 5661 20269 5664
rect 20303 5661 20315 5695
rect 20257 5655 20315 5661
rect 20441 5695 20499 5701
rect 20441 5661 20453 5695
rect 20487 5692 20499 5695
rect 20622 5692 20628 5704
rect 20487 5664 20628 5692
rect 20487 5661 20499 5664
rect 20441 5655 20499 5661
rect 20272 5624 20300 5655
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 20806 5624 20812 5636
rect 9088 5596 9720 5624
rect 17236 5596 17724 5624
rect 20272 5596 20812 5624
rect 9088 5584 9094 5596
rect 7064 5528 7604 5556
rect 8021 5559 8079 5565
rect 7064 5516 7070 5528
rect 8021 5525 8033 5559
rect 8067 5556 8079 5559
rect 8202 5556 8208 5568
rect 8067 5528 8208 5556
rect 8067 5525 8079 5528
rect 8021 5519 8079 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 8297 5559 8355 5565
rect 8297 5525 8309 5559
rect 8343 5556 8355 5559
rect 10870 5556 10876 5568
rect 8343 5528 10876 5556
rect 8343 5525 8355 5528
rect 8297 5519 8355 5525
rect 10870 5516 10876 5528
rect 10928 5516 10934 5568
rect 12069 5559 12127 5565
rect 12069 5525 12081 5559
rect 12115 5556 12127 5559
rect 13170 5556 13176 5568
rect 12115 5528 13176 5556
rect 12115 5525 12127 5528
rect 12069 5519 12127 5525
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 14550 5516 14556 5568
rect 14608 5556 14614 5568
rect 14921 5559 14979 5565
rect 14921 5556 14933 5559
rect 14608 5528 14933 5556
rect 14608 5516 14614 5528
rect 14921 5525 14933 5528
rect 14967 5525 14979 5559
rect 14921 5519 14979 5525
rect 15657 5559 15715 5565
rect 15657 5525 15669 5559
rect 15703 5556 15715 5559
rect 17236 5556 17264 5596
rect 15703 5528 17264 5556
rect 17405 5559 17463 5565
rect 15703 5525 15715 5528
rect 15657 5519 15715 5525
rect 17405 5525 17417 5559
rect 17451 5556 17463 5559
rect 17494 5556 17500 5568
rect 17451 5528 17500 5556
rect 17451 5525 17463 5528
rect 17405 5519 17463 5525
rect 17494 5516 17500 5528
rect 17552 5556 17558 5568
rect 17589 5559 17647 5565
rect 17589 5556 17601 5559
rect 17552 5528 17601 5556
rect 17552 5516 17558 5528
rect 17589 5525 17601 5528
rect 17635 5525 17647 5559
rect 17696 5556 17724 5596
rect 20806 5584 20812 5596
rect 20864 5584 20870 5636
rect 22462 5556 22468 5568
rect 17696 5528 22468 5556
rect 17589 5519 17647 5525
rect 22462 5516 22468 5528
rect 22520 5516 22526 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 1946 5312 1952 5364
rect 2004 5352 2010 5364
rect 2004 5324 3740 5352
rect 2004 5312 2010 5324
rect 3234 5244 3240 5296
rect 3292 5284 3298 5296
rect 3329 5287 3387 5293
rect 3329 5284 3341 5287
rect 3292 5256 3341 5284
rect 3292 5244 3298 5256
rect 3329 5253 3341 5256
rect 3375 5253 3387 5287
rect 3329 5247 3387 5253
rect 1394 5108 1400 5160
rect 1452 5148 1458 5160
rect 1946 5148 1952 5160
rect 1452 5120 1952 5148
rect 1452 5108 1458 5120
rect 1946 5108 1952 5120
rect 2004 5108 2010 5160
rect 3712 5157 3740 5324
rect 3970 5312 3976 5364
rect 4028 5352 4034 5364
rect 8938 5352 8944 5364
rect 4028 5324 8800 5352
rect 8899 5324 8944 5352
rect 4028 5312 4034 5324
rect 5077 5287 5135 5293
rect 5077 5253 5089 5287
rect 5123 5253 5135 5287
rect 8772 5284 8800 5324
rect 8938 5312 8944 5324
rect 8996 5312 9002 5364
rect 9030 5312 9036 5364
rect 9088 5352 9094 5364
rect 9217 5355 9275 5361
rect 9217 5352 9229 5355
rect 9088 5324 9229 5352
rect 9088 5312 9094 5324
rect 9217 5321 9229 5324
rect 9263 5321 9275 5355
rect 9217 5315 9275 5321
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 12526 5352 12532 5364
rect 12483 5324 12532 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 12526 5312 12532 5324
rect 12584 5312 12590 5364
rect 13446 5312 13452 5364
rect 13504 5352 13510 5364
rect 15838 5352 15844 5364
rect 13504 5324 15844 5352
rect 13504 5312 13510 5324
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 16022 5352 16028 5364
rect 15983 5324 16028 5352
rect 16022 5312 16028 5324
rect 16080 5312 16086 5364
rect 16945 5355 17003 5361
rect 16945 5321 16957 5355
rect 16991 5352 17003 5355
rect 17310 5352 17316 5364
rect 16991 5324 17316 5352
rect 16991 5321 17003 5324
rect 16945 5315 17003 5321
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 18601 5355 18659 5361
rect 18601 5321 18613 5355
rect 18647 5352 18659 5355
rect 18690 5352 18696 5364
rect 18647 5324 18696 5352
rect 18647 5321 18659 5324
rect 18601 5315 18659 5321
rect 18690 5312 18696 5324
rect 18748 5312 18754 5364
rect 20622 5312 20628 5364
rect 20680 5352 20686 5364
rect 20993 5355 21051 5361
rect 20993 5352 21005 5355
rect 20680 5324 21005 5352
rect 20680 5312 20686 5324
rect 20993 5321 21005 5324
rect 21039 5321 21051 5355
rect 20993 5315 21051 5321
rect 11057 5287 11115 5293
rect 11057 5284 11069 5287
rect 8772 5256 11069 5284
rect 5077 5247 5135 5253
rect 11057 5253 11069 5256
rect 11103 5253 11115 5287
rect 11057 5247 11115 5253
rect 11149 5287 11207 5293
rect 11149 5253 11161 5287
rect 11195 5284 11207 5287
rect 12894 5284 12900 5296
rect 11195 5256 12900 5284
rect 11195 5253 11207 5256
rect 11149 5247 11207 5253
rect 5092 5216 5120 5247
rect 12894 5244 12900 5256
rect 12952 5244 12958 5296
rect 14090 5284 14096 5296
rect 13004 5256 14096 5284
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5092 5188 6009 5216
rect 5997 5185 6009 5188
rect 6043 5216 6055 5219
rect 6178 5216 6184 5228
rect 6043 5188 6184 5216
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5216 7067 5219
rect 7098 5216 7104 5228
rect 7055 5188 7104 5216
rect 7055 5185 7067 5188
rect 7009 5179 7067 5185
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5216 10839 5219
rect 11330 5216 11336 5228
rect 10827 5188 11336 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 3697 5151 3755 5157
rect 3697 5117 3709 5151
rect 3743 5117 3755 5151
rect 3697 5111 3755 5117
rect 2216 5083 2274 5089
rect 2216 5049 2228 5083
rect 2262 5080 2274 5083
rect 2774 5080 2780 5092
rect 2262 5052 2780 5080
rect 2262 5049 2274 5052
rect 2216 5043 2274 5049
rect 2774 5040 2780 5052
rect 2832 5040 2838 5092
rect 3712 5012 3740 5111
rect 3786 5108 3792 5160
rect 3844 5148 3850 5160
rect 3953 5151 4011 5157
rect 3953 5148 3965 5151
rect 3844 5120 3965 5148
rect 3844 5108 3850 5120
rect 3953 5117 3965 5120
rect 3999 5117 4011 5151
rect 3953 5111 4011 5117
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 6730 5148 6736 5160
rect 5767 5120 6736 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 7558 5148 7564 5160
rect 7519 5120 7564 5148
rect 7558 5108 7564 5120
rect 7616 5108 7622 5160
rect 9401 5151 9459 5157
rect 9401 5148 9413 5151
rect 7668 5120 9413 5148
rect 4062 5040 4068 5092
rect 4120 5080 4126 5092
rect 4120 5052 5948 5080
rect 4120 5040 4126 5052
rect 4706 5012 4712 5024
rect 3712 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 5350 5012 5356 5024
rect 5311 4984 5356 5012
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5626 4972 5632 5024
rect 5684 5012 5690 5024
rect 5813 5015 5871 5021
rect 5813 5012 5825 5015
rect 5684 4984 5825 5012
rect 5684 4972 5690 4984
rect 5813 4981 5825 4984
rect 5859 4981 5871 5015
rect 5920 5012 5948 5052
rect 6454 5040 6460 5092
rect 6512 5080 6518 5092
rect 7668 5080 7696 5120
rect 9401 5117 9413 5120
rect 9447 5117 9459 5151
rect 9401 5111 9459 5117
rect 10318 5108 10324 5160
rect 10376 5148 10382 5160
rect 10796 5148 10824 5179
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 11882 5216 11888 5228
rect 11839 5188 11888 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 13004 5216 13032 5256
rect 14090 5244 14096 5256
rect 14148 5244 14154 5296
rect 16577 5287 16635 5293
rect 16577 5253 16589 5287
rect 16623 5284 16635 5287
rect 18046 5284 18052 5296
rect 16623 5256 18052 5284
rect 16623 5253 16635 5256
rect 16577 5247 16635 5253
rect 18046 5244 18052 5256
rect 18104 5244 18110 5296
rect 18233 5287 18291 5293
rect 18233 5253 18245 5287
rect 18279 5284 18291 5287
rect 19610 5284 19616 5296
rect 18279 5256 19616 5284
rect 18279 5253 18291 5256
rect 18233 5247 18291 5253
rect 19610 5244 19616 5256
rect 19668 5244 19674 5296
rect 11992 5188 13032 5216
rect 13081 5219 13139 5225
rect 10376 5120 10824 5148
rect 11057 5151 11115 5157
rect 10376 5108 10382 5120
rect 11057 5117 11069 5151
rect 11103 5148 11115 5151
rect 11609 5151 11667 5157
rect 11609 5148 11621 5151
rect 11103 5120 11621 5148
rect 11103 5117 11115 5120
rect 11057 5111 11115 5117
rect 11609 5117 11621 5120
rect 11655 5148 11667 5151
rect 11992 5148 12020 5188
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 13354 5216 13360 5228
rect 13127 5188 13360 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 14277 5219 14335 5225
rect 14277 5185 14289 5219
rect 14323 5185 14335 5219
rect 14277 5179 14335 5185
rect 11655 5120 12020 5148
rect 11655 5117 11667 5120
rect 11609 5111 11667 5117
rect 12802 5108 12808 5160
rect 12860 5148 12866 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12860 5120 12909 5148
rect 12860 5108 12866 5120
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 14292 5148 14320 5179
rect 14642 5176 14648 5228
rect 14700 5216 14706 5228
rect 14700 5188 14745 5216
rect 14700 5176 14706 5188
rect 16942 5176 16948 5228
rect 17000 5216 17006 5228
rect 17405 5219 17463 5225
rect 17405 5216 17417 5219
rect 17000 5188 17417 5216
rect 17000 5176 17006 5188
rect 17405 5185 17417 5188
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 17494 5176 17500 5228
rect 17552 5216 17558 5228
rect 18966 5216 18972 5228
rect 17552 5188 17597 5216
rect 17972 5188 18972 5216
rect 17552 5176 17558 5188
rect 16298 5148 16304 5160
rect 14292 5120 16304 5148
rect 12897 5111 12955 5117
rect 16298 5108 16304 5120
rect 16356 5108 16362 5160
rect 16393 5151 16451 5157
rect 16393 5117 16405 5151
rect 16439 5148 16451 5151
rect 17972 5148 18000 5188
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 19245 5219 19303 5225
rect 19245 5185 19257 5219
rect 19291 5185 19303 5219
rect 19245 5179 19303 5185
rect 16439 5120 18000 5148
rect 18049 5151 18107 5157
rect 16439 5117 16451 5120
rect 16393 5111 16451 5117
rect 18049 5117 18061 5151
rect 18095 5148 18107 5151
rect 18874 5148 18880 5160
rect 18095 5120 18880 5148
rect 18095 5117 18107 5120
rect 18049 5111 18107 5117
rect 18874 5108 18880 5120
rect 18932 5108 18938 5160
rect 6512 5052 7696 5080
rect 7828 5083 7886 5089
rect 6512 5040 6518 5052
rect 7828 5049 7840 5083
rect 7874 5080 7886 5083
rect 8202 5080 8208 5092
rect 7874 5052 8208 5080
rect 7874 5049 7886 5052
rect 7828 5043 7886 5049
rect 8202 5040 8208 5052
rect 8260 5040 8266 5092
rect 10505 5083 10563 5089
rect 10505 5080 10517 5083
rect 8312 5052 10517 5080
rect 8312 5012 8340 5052
rect 10505 5049 10517 5052
rect 10551 5049 10563 5083
rect 10505 5043 10563 5049
rect 10594 5040 10600 5092
rect 10652 5080 10658 5092
rect 10652 5052 10697 5080
rect 10652 5040 10658 5052
rect 11238 5040 11244 5092
rect 11296 5080 11302 5092
rect 14093 5083 14151 5089
rect 14093 5080 14105 5083
rect 11296 5052 14105 5080
rect 11296 5040 11302 5052
rect 14093 5049 14105 5052
rect 14139 5049 14151 5083
rect 14093 5043 14151 5049
rect 14912 5083 14970 5089
rect 14912 5049 14924 5083
rect 14958 5080 14970 5083
rect 15194 5080 15200 5092
rect 14958 5052 15200 5080
rect 14958 5049 14970 5052
rect 14912 5043 14970 5049
rect 15194 5040 15200 5052
rect 15252 5040 15258 5092
rect 17313 5083 17371 5089
rect 17313 5049 17325 5083
rect 17359 5080 17371 5083
rect 18782 5080 18788 5092
rect 17359 5052 18788 5080
rect 17359 5049 17371 5052
rect 17313 5043 17371 5049
rect 18782 5040 18788 5052
rect 18840 5040 18846 5092
rect 19260 5080 19288 5179
rect 19518 5108 19524 5160
rect 19576 5148 19582 5160
rect 19613 5151 19671 5157
rect 19613 5148 19625 5151
rect 19576 5120 19625 5148
rect 19576 5108 19582 5120
rect 19613 5117 19625 5120
rect 19659 5117 19671 5151
rect 19613 5111 19671 5117
rect 19880 5083 19938 5089
rect 19880 5080 19892 5083
rect 19260 5052 19892 5080
rect 19880 5049 19892 5052
rect 19926 5080 19938 5083
rect 20162 5080 20168 5092
rect 19926 5052 20168 5080
rect 19926 5049 19938 5052
rect 19880 5043 19938 5049
rect 20162 5040 20168 5052
rect 20220 5040 20226 5092
rect 5920 4984 8340 5012
rect 10137 5015 10195 5021
rect 5813 4975 5871 4981
rect 10137 4981 10149 5015
rect 10183 5012 10195 5015
rect 10778 5012 10784 5024
rect 10183 4984 10784 5012
rect 10183 4981 10195 4984
rect 10137 4975 10195 4981
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 11422 4972 11428 5024
rect 11480 5012 11486 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 11480 4984 11529 5012
rect 11480 4972 11486 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 12802 5012 12808 5024
rect 12763 4984 12808 5012
rect 11517 4975 11575 4981
rect 12802 4972 12808 4984
rect 12860 4972 12866 5024
rect 13630 5012 13636 5024
rect 13591 4984 13636 5012
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 13722 4972 13728 5024
rect 13780 5012 13786 5024
rect 14001 5015 14059 5021
rect 14001 5012 14013 5015
rect 13780 4984 14013 5012
rect 13780 4972 13786 4984
rect 14001 4981 14013 4984
rect 14047 4981 14059 5015
rect 14001 4975 14059 4981
rect 16758 4972 16764 5024
rect 16816 5012 16822 5024
rect 17494 5012 17500 5024
rect 16816 4984 17500 5012
rect 16816 4972 16822 4984
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 18690 4972 18696 5024
rect 18748 5012 18754 5024
rect 18969 5015 19027 5021
rect 18969 5012 18981 5015
rect 18748 4984 18981 5012
rect 18748 4972 18754 4984
rect 18969 4981 18981 4984
rect 19015 4981 19027 5015
rect 18969 4975 19027 4981
rect 19061 5015 19119 5021
rect 19061 4981 19073 5015
rect 19107 5012 19119 5015
rect 19978 5012 19984 5024
rect 19107 4984 19984 5012
rect 19107 4981 19119 4984
rect 19061 4975 19119 4981
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 2832 4780 2877 4808
rect 2832 4768 2838 4780
rect 3878 4768 3884 4820
rect 3936 4808 3942 4820
rect 6086 4808 6092 4820
rect 3936 4780 6092 4808
rect 3936 4768 3942 4780
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 7006 4808 7012 4820
rect 6967 4780 7012 4808
rect 7006 4768 7012 4780
rect 7064 4768 7070 4820
rect 7466 4768 7472 4820
rect 7524 4808 7530 4820
rect 7742 4808 7748 4820
rect 7524 4780 7748 4808
rect 7524 4768 7530 4780
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 8113 4811 8171 4817
rect 8113 4777 8125 4811
rect 8159 4808 8171 4811
rect 8294 4808 8300 4820
rect 8159 4780 8300 4808
rect 8159 4777 8171 4780
rect 8113 4771 8171 4777
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 8481 4811 8539 4817
rect 8481 4777 8493 4811
rect 8527 4808 8539 4811
rect 9677 4811 9735 4817
rect 9677 4808 9689 4811
rect 8527 4780 9689 4808
rect 8527 4777 8539 4780
rect 8481 4771 8539 4777
rect 9677 4777 9689 4780
rect 9723 4777 9735 4811
rect 9677 4771 9735 4777
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 13081 4811 13139 4817
rect 13081 4808 13093 4811
rect 11480 4780 13093 4808
rect 11480 4768 11486 4780
rect 13081 4777 13093 4780
rect 13127 4777 13139 4811
rect 13081 4771 13139 4777
rect 13630 4768 13636 4820
rect 13688 4808 13694 4820
rect 16025 4811 16083 4817
rect 16025 4808 16037 4811
rect 13688 4780 16037 4808
rect 13688 4768 13694 4780
rect 16025 4777 16037 4780
rect 16071 4777 16083 4811
rect 16025 4771 16083 4777
rect 16482 4768 16488 4820
rect 16540 4808 16546 4820
rect 17126 4808 17132 4820
rect 16540 4780 17132 4808
rect 16540 4768 16546 4780
rect 17126 4768 17132 4780
rect 17184 4808 17190 4820
rect 18509 4811 18567 4817
rect 17184 4780 17908 4808
rect 17184 4768 17190 4780
rect 4792 4743 4850 4749
rect 4792 4709 4804 4743
rect 4838 4740 4850 4743
rect 6178 4740 6184 4752
rect 4838 4712 6184 4740
rect 4838 4709 4850 4712
rect 4792 4703 4850 4709
rect 6178 4700 6184 4712
rect 6236 4700 6242 4752
rect 6822 4700 6828 4752
rect 6880 4740 6886 4752
rect 8570 4740 8576 4752
rect 6880 4712 7972 4740
rect 8531 4712 8576 4740
rect 6880 4700 6886 4712
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 1664 4675 1722 4681
rect 1664 4641 1676 4675
rect 1710 4672 1722 4675
rect 3142 4672 3148 4684
rect 1710 4644 3148 4672
rect 1710 4641 1722 4644
rect 1664 4635 1722 4641
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 4525 4675 4583 4681
rect 4525 4641 4537 4675
rect 4571 4672 4583 4675
rect 4614 4672 4620 4684
rect 4571 4644 4620 4672
rect 4571 4641 4583 4644
rect 4525 4635 4583 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 6914 4672 6920 4684
rect 6875 4644 6920 4672
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7944 4672 7972 4712
rect 8570 4700 8576 4712
rect 8628 4700 8634 4752
rect 11238 4740 11244 4752
rect 9876 4712 11244 4740
rect 9876 4672 9904 4712
rect 11238 4700 11244 4712
rect 11296 4700 11302 4752
rect 11330 4700 11336 4752
rect 11388 4740 11394 4752
rect 11882 4740 11888 4752
rect 11388 4712 11888 4740
rect 11388 4700 11394 4712
rect 11882 4700 11888 4712
rect 11940 4740 11946 4752
rect 12986 4740 12992 4752
rect 11940 4712 12992 4740
rect 11940 4700 11946 4712
rect 12986 4700 12992 4712
rect 13044 4700 13050 4752
rect 13808 4743 13866 4749
rect 13808 4709 13820 4743
rect 13854 4740 13866 4743
rect 14550 4740 14556 4752
rect 13854 4712 14556 4740
rect 13854 4709 13866 4712
rect 13808 4703 13866 4709
rect 14550 4700 14556 4712
rect 14608 4700 14614 4752
rect 16577 4743 16635 4749
rect 16577 4709 16589 4743
rect 16623 4740 16635 4743
rect 17770 4740 17776 4752
rect 16623 4712 17776 4740
rect 16623 4709 16635 4712
rect 16577 4703 16635 4709
rect 17770 4700 17776 4712
rect 17828 4700 17834 4752
rect 10042 4672 10048 4684
rect 7944 4644 9904 4672
rect 10003 4644 10048 4672
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 10873 4675 10931 4681
rect 10873 4641 10885 4675
rect 10919 4672 10931 4675
rect 11514 4672 11520 4684
rect 10919 4644 11520 4672
rect 10919 4641 10931 4644
rect 10873 4635 10931 4641
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 11692 4675 11750 4681
rect 11692 4641 11704 4675
rect 11738 4672 11750 4675
rect 13446 4672 13452 4684
rect 11738 4644 13452 4672
rect 11738 4641 11750 4644
rect 11692 4635 11750 4641
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 13538 4632 13544 4684
rect 13596 4672 13602 4684
rect 13596 4644 13641 4672
rect 13596 4632 13602 4644
rect 15102 4632 15108 4684
rect 15160 4672 15166 4684
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 15160 4644 15301 4672
rect 15160 4632 15166 4644
rect 15289 4641 15301 4644
rect 15335 4641 15347 4675
rect 15289 4635 15347 4641
rect 16025 4675 16083 4681
rect 16025 4641 16037 4675
rect 16071 4672 16083 4675
rect 16485 4675 16543 4681
rect 16485 4672 16497 4675
rect 16071 4644 16497 4672
rect 16071 4641 16083 4644
rect 16025 4635 16083 4641
rect 16485 4641 16497 4644
rect 16531 4641 16543 4675
rect 17126 4672 17132 4684
rect 17087 4644 17132 4672
rect 16485 4635 16543 4641
rect 17126 4632 17132 4644
rect 17184 4632 17190 4684
rect 17402 4681 17408 4684
rect 17396 4672 17408 4681
rect 17363 4644 17408 4672
rect 17396 4635 17408 4644
rect 17402 4632 17408 4635
rect 17460 4632 17466 4684
rect 17880 4672 17908 4780
rect 18509 4777 18521 4811
rect 18555 4777 18567 4811
rect 20162 4808 20168 4820
rect 20123 4780 20168 4808
rect 18509 4771 18567 4777
rect 18524 4740 18552 4771
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 19058 4749 19064 4752
rect 19030 4743 19064 4749
rect 19030 4740 19042 4743
rect 18524 4712 19042 4740
rect 19030 4709 19042 4712
rect 19116 4740 19122 4752
rect 19116 4712 19178 4740
rect 19030 4703 19064 4709
rect 19058 4700 19064 4703
rect 19116 4700 19122 4712
rect 18785 4675 18843 4681
rect 18785 4672 18797 4675
rect 17880 4644 18797 4672
rect 18785 4641 18797 4644
rect 18831 4672 18843 4675
rect 19518 4672 19524 4684
rect 18831 4644 19524 4672
rect 18831 4641 18843 4644
rect 18785 4635 18843 4641
rect 19518 4632 19524 4644
rect 19576 4632 19582 4684
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 7156 4576 7201 4604
rect 7156 4564 7162 4576
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 8665 4607 8723 4613
rect 8665 4604 8677 4607
rect 8260 4576 8677 4604
rect 8260 4564 8266 4576
rect 8665 4573 8677 4576
rect 8711 4573 8723 4607
rect 8665 4567 8723 4573
rect 9950 4564 9956 4616
rect 10008 4604 10014 4616
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 10008 4576 10149 4604
rect 10008 4564 10014 4576
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4573 11483 4607
rect 16758 4604 16764 4616
rect 16719 4576 16764 4604
rect 11425 4567 11483 4573
rect 5626 4496 5632 4548
rect 5684 4536 5690 4548
rect 5684 4508 9168 4536
rect 5684 4496 5690 4508
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 5905 4471 5963 4477
rect 5905 4468 5917 4471
rect 5316 4440 5917 4468
rect 5316 4428 5322 4440
rect 5905 4437 5917 4440
rect 5951 4437 5963 4471
rect 5905 4431 5963 4437
rect 6549 4471 6607 4477
rect 6549 4437 6561 4471
rect 6595 4468 6607 4471
rect 7190 4468 7196 4480
rect 6595 4440 7196 4468
rect 6595 4437 6607 4440
rect 6549 4431 6607 4437
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 9140 4468 9168 4508
rect 9214 4496 9220 4548
rect 9272 4536 9278 4548
rect 10244 4536 10272 4567
rect 9272 4508 10272 4536
rect 9272 4496 9278 4508
rect 10594 4468 10600 4480
rect 9140 4440 10600 4468
rect 10594 4428 10600 4440
rect 10652 4428 10658 4480
rect 11054 4468 11060 4480
rect 11015 4440 11060 4468
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 11440 4468 11468 4567
rect 16758 4564 16764 4576
rect 16816 4564 16822 4616
rect 16117 4539 16175 4545
rect 16117 4505 16129 4539
rect 16163 4536 16175 4539
rect 16666 4536 16672 4548
rect 16163 4508 16672 4536
rect 16163 4505 16175 4508
rect 16117 4499 16175 4505
rect 16666 4496 16672 4508
rect 16724 4496 16730 4548
rect 12342 4468 12348 4480
rect 11440 4440 12348 4468
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 12805 4471 12863 4477
rect 12805 4437 12817 4471
rect 12851 4468 12863 4471
rect 12986 4468 12992 4480
rect 12851 4440 12992 4468
rect 12851 4437 12863 4440
rect 12805 4431 12863 4437
rect 12986 4428 12992 4440
rect 13044 4428 13050 4480
rect 14918 4468 14924 4480
rect 14879 4440 14924 4468
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15473 4471 15531 4477
rect 15473 4437 15485 4471
rect 15519 4468 15531 4471
rect 15838 4468 15844 4480
rect 15519 4440 15844 4468
rect 15519 4437 15531 4440
rect 15473 4431 15531 4437
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 18782 4428 18788 4480
rect 18840 4468 18846 4480
rect 21082 4468 21088 4480
rect 18840 4440 21088 4468
rect 18840 4428 18846 4440
rect 21082 4428 21088 4440
rect 21140 4428 21146 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 4706 4264 4712 4276
rect 2976 4236 4712 4264
rect 2774 4196 2780 4208
rect 2608 4168 2780 4196
rect 2608 4137 2636 4168
rect 2774 4156 2780 4168
rect 2832 4156 2838 4208
rect 2976 4137 3004 4236
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 7374 4264 7380 4276
rect 6012 4236 7380 4264
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4097 2651 4131
rect 2593 4091 2651 4097
rect 2961 4131 3019 4137
rect 2961 4097 2973 4131
rect 3007 4097 3019 4131
rect 5258 4128 5264 4140
rect 2961 4091 3019 4097
rect 4724 4100 5264 4128
rect 3228 4063 3286 4069
rect 3228 4029 3240 4063
rect 3274 4060 3286 4063
rect 4724 4060 4752 4100
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 3274 4032 4752 4060
rect 5077 4063 5135 4069
rect 3274 4029 3286 4032
rect 3228 4023 3286 4029
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 5350 4060 5356 4072
rect 5123 4032 5356 4060
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 6012 4069 6040 4236
rect 6825 4199 6883 4205
rect 6825 4165 6837 4199
rect 6871 4165 6883 4199
rect 6825 4159 6883 4165
rect 6178 4128 6184 4140
rect 6139 4100 6184 4128
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4029 6055 4063
rect 5997 4023 6055 4029
rect 3142 3952 3148 4004
rect 3200 3992 3206 4004
rect 4985 3995 5043 4001
rect 3200 3964 4384 3992
rect 3200 3952 3206 3964
rect 1762 3884 1768 3936
rect 1820 3924 1826 3936
rect 1949 3927 2007 3933
rect 1949 3924 1961 3927
rect 1820 3896 1961 3924
rect 1820 3884 1826 3896
rect 1949 3893 1961 3896
rect 1995 3893 2007 3927
rect 2314 3924 2320 3936
rect 2275 3896 2320 3924
rect 1949 3887 2007 3893
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 2409 3927 2467 3933
rect 2409 3893 2421 3927
rect 2455 3924 2467 3927
rect 4062 3924 4068 3936
rect 2455 3896 4068 3924
rect 2455 3893 2467 3896
rect 2409 3887 2467 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4356 3933 4384 3964
rect 4985 3961 4997 3995
rect 5031 3992 5043 3995
rect 5031 3964 5672 3992
rect 5031 3961 5043 3964
rect 4985 3955 5043 3961
rect 4341 3927 4399 3933
rect 4341 3893 4353 3927
rect 4387 3893 4399 3927
rect 4341 3887 4399 3893
rect 4522 3884 4528 3936
rect 4580 3924 4586 3936
rect 5644 3933 5672 3964
rect 5718 3952 5724 4004
rect 5776 3992 5782 4004
rect 6089 3995 6147 4001
rect 6089 3992 6101 3995
rect 5776 3964 6101 3992
rect 5776 3952 5782 3964
rect 6089 3961 6101 3964
rect 6135 3992 6147 3995
rect 6638 3992 6644 4004
rect 6135 3964 6644 3992
rect 6135 3961 6147 3964
rect 6089 3955 6147 3961
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 6840 3992 6868 4159
rect 7300 4072 7328 4236
rect 7374 4224 7380 4236
rect 7432 4224 7438 4276
rect 9214 4264 9220 4276
rect 9175 4236 9220 4264
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 10226 4224 10232 4276
rect 10284 4264 10290 4276
rect 10284 4236 10999 4264
rect 10284 4224 10290 4236
rect 10971 4196 10999 4236
rect 11054 4224 11060 4276
rect 11112 4264 11118 4276
rect 19978 4264 19984 4276
rect 11112 4236 16804 4264
rect 19939 4236 19984 4264
rect 11112 4224 11118 4236
rect 13722 4196 13728 4208
rect 10971 4168 13728 4196
rect 13722 4156 13728 4168
rect 13780 4156 13786 4208
rect 14918 4156 14924 4208
rect 14976 4196 14982 4208
rect 16577 4199 16635 4205
rect 14976 4168 16068 4196
rect 14976 4156 14982 4168
rect 7466 4128 7472 4140
rect 7427 4100 7472 4128
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 7558 4088 7564 4140
rect 7616 4088 7622 4140
rect 12986 4128 12992 4140
rect 11072 4100 12848 4128
rect 12947 4100 12992 4128
rect 7190 4060 7196 4072
rect 7151 4032 7196 4060
rect 7190 4020 7196 4032
rect 7248 4020 7254 4072
rect 7282 4020 7288 4072
rect 7340 4020 7346 4072
rect 7576 4060 7604 4088
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 7576 4032 7849 4060
rect 7837 4029 7849 4032
rect 7883 4060 7895 4063
rect 8386 4060 8392 4072
rect 7883 4032 8392 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 8386 4020 8392 4032
rect 8444 4060 8450 4072
rect 9030 4060 9036 4072
rect 8444 4032 9036 4060
rect 8444 4020 8450 4032
rect 9030 4020 9036 4032
rect 9088 4060 9094 4072
rect 9582 4060 9588 4072
rect 9088 4032 9588 4060
rect 9088 4020 9094 4032
rect 9582 4020 9588 4032
rect 9640 4060 9646 4072
rect 10318 4069 10324 4072
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 9640 4032 10057 4060
rect 9640 4020 9646 4032
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 10312 4060 10324 4069
rect 10279 4032 10324 4060
rect 10045 4023 10103 4029
rect 10312 4023 10324 4032
rect 10318 4020 10324 4023
rect 10376 4020 10382 4072
rect 7558 3992 7564 4004
rect 6840 3964 7564 3992
rect 7558 3952 7564 3964
rect 7616 3952 7622 4004
rect 8104 3995 8162 4001
rect 8104 3961 8116 3995
rect 8150 3992 8162 3995
rect 8202 3992 8208 4004
rect 8150 3964 8208 3992
rect 8150 3961 8162 3964
rect 8104 3955 8162 3961
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 8846 3952 8852 4004
rect 8904 3992 8910 4004
rect 10686 3992 10692 4004
rect 8904 3964 10692 3992
rect 8904 3952 8910 3964
rect 10686 3952 10692 3964
rect 10744 3992 10750 4004
rect 11072 3992 11100 4100
rect 12820 4069 12848 4100
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 16040 4137 16068 4168
rect 16577 4165 16589 4199
rect 16623 4165 16635 4199
rect 16776 4196 16804 4236
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 18782 4196 18788 4208
rect 16776 4168 18788 4196
rect 16577 4159 16635 4165
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4097 16083 4131
rect 16592 4128 16620 4159
rect 18782 4156 18788 4168
rect 18840 4156 18846 4208
rect 19058 4156 19064 4208
rect 19116 4196 19122 4208
rect 19116 4168 20576 4196
rect 19116 4156 19122 4168
rect 17221 4131 17279 4137
rect 16592 4100 17172 4128
rect 16025 4091 16083 4097
rect 11793 4063 11851 4069
rect 11793 4029 11805 4063
rect 11839 4060 11851 4063
rect 12805 4063 12863 4069
rect 11839 4032 12756 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 12618 3992 12624 4004
rect 10744 3964 11100 3992
rect 11992 3964 12624 3992
rect 10744 3952 10750 3964
rect 4617 3927 4675 3933
rect 4617 3924 4629 3927
rect 4580 3896 4629 3924
rect 4580 3884 4586 3896
rect 4617 3893 4629 3896
rect 4663 3893 4675 3927
rect 4617 3887 4675 3893
rect 5629 3927 5687 3933
rect 5629 3893 5641 3927
rect 5675 3893 5687 3927
rect 5629 3887 5687 3893
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 7285 3927 7343 3933
rect 7285 3924 7297 3927
rect 6328 3896 7297 3924
rect 6328 3884 6334 3896
rect 7285 3893 7297 3896
rect 7331 3893 7343 3927
rect 11422 3924 11428 3936
rect 11383 3896 11428 3924
rect 7285 3887 7343 3893
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 11992 3933 12020 3964
rect 12618 3952 12624 3964
rect 12676 3952 12682 4004
rect 12728 3992 12756 4032
rect 12805 4029 12817 4063
rect 12851 4029 12863 4063
rect 12805 4023 12863 4029
rect 12897 4063 12955 4069
rect 12897 4029 12909 4063
rect 12943 4060 12955 4063
rect 13078 4060 13084 4072
rect 12943 4032 13084 4060
rect 12943 4029 12955 4032
rect 12897 4023 12955 4029
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 13538 4020 13544 4072
rect 13596 4060 13602 4072
rect 13817 4063 13875 4069
rect 13817 4060 13829 4063
rect 13596 4032 13829 4060
rect 13596 4020 13602 4032
rect 13817 4029 13829 4032
rect 13863 4029 13875 4063
rect 13817 4023 13875 4029
rect 14084 4063 14142 4069
rect 14084 4029 14096 4063
rect 14130 4060 14142 4063
rect 14918 4060 14924 4072
rect 14130 4032 14924 4060
rect 14130 4029 14142 4032
rect 14084 4023 14142 4029
rect 14918 4020 14924 4032
rect 14976 4020 14982 4072
rect 16850 4020 16856 4072
rect 16908 4060 16914 4072
rect 17037 4063 17095 4069
rect 17037 4060 17049 4063
rect 16908 4032 17049 4060
rect 16908 4020 16914 4032
rect 17037 4029 17049 4032
rect 17083 4029 17095 4063
rect 17144 4060 17172 4100
rect 17221 4097 17233 4131
rect 17267 4128 17279 4131
rect 17402 4128 17408 4140
rect 17267 4100 17408 4128
rect 17267 4097 17279 4100
rect 17221 4091 17279 4097
rect 17402 4088 17408 4100
rect 17460 4128 17466 4140
rect 18598 4128 18604 4140
rect 17460 4100 18604 4128
rect 17460 4088 17466 4100
rect 18598 4088 18604 4100
rect 18656 4128 18662 4140
rect 20548 4137 20576 4168
rect 19521 4131 19579 4137
rect 19521 4128 19533 4131
rect 18656 4100 19533 4128
rect 18656 4088 18662 4100
rect 19521 4097 19533 4100
rect 19567 4097 19579 4131
rect 19521 4091 19579 4097
rect 20533 4131 20591 4137
rect 20533 4097 20545 4131
rect 20579 4097 20591 4131
rect 20533 4091 20591 4097
rect 18322 4060 18328 4072
rect 17144 4032 18328 4060
rect 17037 4023 17095 4029
rect 18322 4020 18328 4032
rect 18380 4020 18386 4072
rect 18417 4063 18475 4069
rect 18417 4029 18429 4063
rect 18463 4060 18475 4063
rect 19334 4060 19340 4072
rect 18463 4032 19340 4060
rect 18463 4029 18475 4032
rect 18417 4023 18475 4029
rect 19334 4020 19340 4032
rect 19392 4020 19398 4072
rect 20438 4020 20444 4072
rect 20496 4060 20502 4072
rect 21542 4060 21548 4072
rect 20496 4032 21548 4060
rect 20496 4020 20502 4032
rect 21542 4020 21548 4032
rect 21600 4020 21606 4072
rect 13722 3992 13728 4004
rect 12728 3964 13728 3992
rect 13722 3952 13728 3964
rect 13780 3952 13786 4004
rect 15841 3995 15899 4001
rect 15841 3992 15853 3995
rect 14200 3964 15853 3992
rect 11977 3927 12035 3933
rect 11977 3893 11989 3927
rect 12023 3893 12035 3927
rect 11977 3887 12035 3893
rect 12158 3884 12164 3936
rect 12216 3924 12222 3936
rect 12437 3927 12495 3933
rect 12437 3924 12449 3927
rect 12216 3896 12449 3924
rect 12216 3884 12222 3896
rect 12437 3893 12449 3896
rect 12483 3893 12495 3927
rect 12437 3887 12495 3893
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 14200 3924 14228 3964
rect 15841 3961 15853 3964
rect 15887 3961 15899 3995
rect 15841 3955 15899 3961
rect 15933 3995 15991 4001
rect 15933 3961 15945 3995
rect 15979 3992 15991 3995
rect 16114 3992 16120 4004
rect 15979 3964 16120 3992
rect 15979 3961 15991 3964
rect 15933 3955 15991 3961
rect 16114 3952 16120 3964
rect 16172 3952 16178 4004
rect 16945 3995 17003 4001
rect 16945 3961 16957 3995
rect 16991 3992 17003 3995
rect 17218 3992 17224 4004
rect 16991 3964 17224 3992
rect 16991 3961 17003 3964
rect 16945 3955 17003 3961
rect 17218 3952 17224 3964
rect 17276 3952 17282 4004
rect 17954 3952 17960 4004
rect 18012 3992 18018 4004
rect 20530 3992 20536 4004
rect 18012 3964 20536 3992
rect 18012 3952 18018 3964
rect 20530 3952 20536 3964
rect 20588 3952 20594 4004
rect 15194 3924 15200 3936
rect 13136 3896 14228 3924
rect 15155 3896 15200 3924
rect 13136 3884 13142 3896
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 15473 3927 15531 3933
rect 15473 3893 15485 3927
rect 15519 3924 15531 3927
rect 15746 3924 15752 3936
rect 15519 3896 15752 3924
rect 15519 3893 15531 3896
rect 15473 3887 15531 3893
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 18230 3924 18236 3936
rect 17092 3896 18236 3924
rect 17092 3884 17098 3896
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 18601 3927 18659 3933
rect 18601 3893 18613 3927
rect 18647 3924 18659 3927
rect 18782 3924 18788 3936
rect 18647 3896 18788 3924
rect 18647 3893 18659 3896
rect 18601 3887 18659 3893
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 18966 3924 18972 3936
rect 18927 3896 18972 3924
rect 18966 3884 18972 3896
rect 19024 3884 19030 3936
rect 19334 3924 19340 3936
rect 19295 3896 19340 3924
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 19426 3884 19432 3936
rect 19484 3924 19490 3936
rect 20346 3924 20352 3936
rect 19484 3896 19529 3924
rect 20307 3896 20352 3924
rect 19484 3884 19490 3896
rect 20346 3884 20352 3896
rect 20404 3884 20410 3936
rect 20438 3884 20444 3936
rect 20496 3924 20502 3936
rect 20496 3896 20541 3924
rect 20496 3884 20502 3896
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 2314 3680 2320 3732
rect 2372 3720 2378 3732
rect 2593 3723 2651 3729
rect 2593 3720 2605 3723
rect 2372 3692 2605 3720
rect 2372 3680 2378 3692
rect 2593 3689 2605 3692
rect 2639 3689 2651 3723
rect 4062 3720 4068 3732
rect 4023 3692 4068 3720
rect 2593 3683 2651 3689
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 4522 3720 4528 3732
rect 4483 3692 4528 3720
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 5077 3723 5135 3729
rect 5077 3689 5089 3723
rect 5123 3689 5135 3723
rect 5077 3683 5135 3689
rect 6365 3723 6423 3729
rect 6365 3689 6377 3723
rect 6411 3720 6423 3723
rect 6914 3720 6920 3732
rect 6411 3692 6920 3720
rect 6411 3689 6423 3692
rect 6365 3683 6423 3689
rect 4433 3655 4491 3661
rect 4433 3621 4445 3655
rect 4479 3652 4491 3655
rect 5092 3652 5120 3683
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 8938 3680 8944 3732
rect 8996 3720 9002 3732
rect 9858 3720 9864 3732
rect 8996 3692 9864 3720
rect 8996 3680 9002 3692
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 13078 3720 13084 3732
rect 10060 3692 13084 3720
rect 10060 3664 10088 3692
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 14185 3723 14243 3729
rect 14185 3689 14197 3723
rect 14231 3689 14243 3723
rect 14185 3683 14243 3689
rect 4479 3624 5120 3652
rect 4479 3621 4491 3624
rect 4433 3615 4491 3621
rect 7190 3612 7196 3664
rect 7248 3652 7254 3664
rect 10042 3652 10048 3664
rect 7248 3624 10048 3652
rect 7248 3612 7254 3624
rect 10042 3612 10048 3624
rect 10100 3612 10106 3664
rect 10312 3655 10370 3661
rect 10312 3621 10324 3655
rect 10358 3652 10370 3655
rect 11422 3652 11428 3664
rect 10358 3624 11428 3652
rect 10358 3621 10370 3624
rect 10312 3615 10370 3621
rect 11422 3612 11428 3624
rect 11480 3652 11486 3664
rect 11882 3652 11888 3664
rect 11480 3624 11888 3652
rect 11480 3612 11486 3624
rect 11882 3612 11888 3624
rect 11940 3612 11946 3664
rect 12802 3652 12808 3664
rect 11992 3624 12808 3652
rect 2961 3587 3019 3593
rect 2961 3553 2973 3587
rect 3007 3584 3019 3587
rect 4154 3584 4160 3596
rect 3007 3556 4160 3584
rect 3007 3553 3019 3556
rect 2961 3547 3019 3553
rect 4154 3544 4160 3556
rect 4212 3544 4218 3596
rect 5442 3544 5448 3596
rect 5500 3584 5506 3596
rect 7092 3587 7150 3593
rect 5500 3556 5545 3584
rect 5500 3544 5506 3556
rect 7092 3553 7104 3587
rect 7138 3584 7150 3587
rect 7466 3584 7472 3596
rect 7138 3556 7472 3584
rect 7138 3553 7150 3556
rect 7092 3547 7150 3553
rect 7466 3544 7472 3556
rect 7524 3584 7530 3596
rect 7524 3556 8156 3584
rect 7524 3544 7530 3556
rect 8128 3528 8156 3556
rect 8570 3544 8576 3596
rect 8628 3584 8634 3596
rect 8849 3587 8907 3593
rect 8849 3584 8861 3587
rect 8628 3556 8861 3584
rect 8628 3544 8634 3556
rect 8849 3553 8861 3556
rect 8895 3553 8907 3587
rect 8849 3547 8907 3553
rect 8941 3587 8999 3593
rect 8941 3553 8953 3587
rect 8987 3584 8999 3587
rect 9858 3584 9864 3596
rect 8987 3556 9864 3584
rect 8987 3553 8999 3556
rect 8941 3547 8999 3553
rect 9858 3544 9864 3556
rect 9916 3544 9922 3596
rect 9950 3544 9956 3596
rect 10008 3584 10014 3596
rect 11992 3584 12020 3624
rect 12802 3612 12808 3624
rect 12860 3652 12866 3664
rect 13173 3655 13231 3661
rect 13173 3652 13185 3655
rect 12860 3624 13185 3652
rect 12860 3612 12866 3624
rect 13173 3621 13185 3624
rect 13219 3621 13231 3655
rect 14200 3652 14228 3683
rect 14274 3680 14280 3732
rect 14332 3720 14338 3732
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 14332 3692 14657 3720
rect 14332 3680 14338 3692
rect 14645 3689 14657 3692
rect 14691 3720 14703 3723
rect 15105 3723 15163 3729
rect 15105 3720 15117 3723
rect 14691 3692 15117 3720
rect 14691 3689 14703 3692
rect 14645 3683 14703 3689
rect 15105 3689 15117 3692
rect 15151 3689 15163 3723
rect 15746 3720 15752 3732
rect 15707 3692 15752 3720
rect 15105 3683 15163 3689
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 18414 3720 18420 3732
rect 16316 3692 18420 3720
rect 15657 3655 15715 3661
rect 15657 3652 15669 3655
rect 14200 3624 15669 3652
rect 13173 3615 13231 3621
rect 15657 3621 15669 3624
rect 15703 3621 15715 3655
rect 15657 3615 15715 3621
rect 10008 3556 12020 3584
rect 12069 3587 12127 3593
rect 10008 3544 10014 3556
rect 12069 3553 12081 3587
rect 12115 3584 12127 3587
rect 12250 3584 12256 3596
rect 12115 3556 12256 3584
rect 12115 3553 12127 3556
rect 12069 3547 12127 3553
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 12618 3544 12624 3596
rect 12676 3584 12682 3596
rect 13725 3587 13783 3593
rect 12676 3556 12756 3584
rect 12676 3544 12682 3556
rect 3050 3516 3056 3528
rect 3011 3488 3056 3516
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 3142 3476 3148 3528
rect 3200 3516 3206 3528
rect 4617 3519 4675 3525
rect 4617 3516 4629 3519
rect 3200 3488 4629 3516
rect 3200 3476 3206 3488
rect 4617 3485 4629 3488
rect 4663 3485 4675 3519
rect 5534 3516 5540 3528
rect 5495 3488 5540 3516
rect 4617 3479 4675 3485
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3485 5779 3519
rect 6822 3516 6828 3528
rect 6783 3488 6828 3516
rect 5721 3479 5779 3485
rect 198 3408 204 3460
rect 256 3448 262 3460
rect 3786 3448 3792 3460
rect 256 3420 3792 3448
rect 256 3408 262 3420
rect 3786 3408 3792 3420
rect 3844 3408 3850 3460
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 5736 3448 5764 3479
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 9033 3519 9091 3525
rect 9033 3516 9045 3519
rect 8168 3488 9045 3516
rect 8168 3476 8174 3488
rect 9033 3485 9045 3488
rect 9079 3485 9091 3519
rect 9033 3479 9091 3485
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 10045 3519 10103 3525
rect 10045 3516 10057 3519
rect 9640 3488 10057 3516
rect 9640 3476 9646 3488
rect 10045 3485 10057 3488
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 11606 3476 11612 3528
rect 11664 3516 11670 3528
rect 12161 3519 12219 3525
rect 12161 3516 12173 3519
rect 11664 3488 12173 3516
rect 11664 3476 11670 3488
rect 12161 3485 12173 3488
rect 12207 3485 12219 3519
rect 12161 3479 12219 3485
rect 12345 3519 12403 3525
rect 12345 3485 12357 3519
rect 12391 3516 12403 3519
rect 12529 3519 12587 3525
rect 12529 3516 12541 3519
rect 12391 3488 12541 3516
rect 12391 3485 12403 3488
rect 12345 3479 12403 3485
rect 12529 3485 12541 3488
rect 12575 3485 12587 3519
rect 12529 3479 12587 3485
rect 11701 3451 11759 3457
rect 5316 3420 5764 3448
rect 7760 3420 8616 3448
rect 5316 3408 5322 3420
rect 7760 3392 7788 3420
rect 3970 3340 3976 3392
rect 4028 3380 4034 3392
rect 5718 3380 5724 3392
rect 4028 3352 5724 3380
rect 4028 3340 4034 3352
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 5902 3340 5908 3392
rect 5960 3380 5966 3392
rect 7742 3380 7748 3392
rect 5960 3352 7748 3380
rect 5960 3340 5966 3352
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 8202 3380 8208 3392
rect 8163 3352 8208 3380
rect 8202 3340 8208 3352
rect 8260 3340 8266 3392
rect 8478 3380 8484 3392
rect 8439 3352 8484 3380
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 8588 3380 8616 3420
rect 11701 3417 11713 3451
rect 11747 3448 11759 3451
rect 12618 3448 12624 3460
rect 11747 3420 12624 3448
rect 11747 3417 11759 3420
rect 11701 3411 11759 3417
rect 12618 3408 12624 3420
rect 12676 3408 12682 3460
rect 12728 3448 12756 3556
rect 13725 3553 13737 3587
rect 13771 3584 13783 3587
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 13771 3556 14565 3584
rect 13771 3553 13783 3556
rect 13725 3547 13783 3553
rect 14553 3553 14565 3556
rect 14599 3553 14611 3587
rect 14553 3547 14611 3553
rect 15105 3587 15163 3593
rect 15105 3553 15117 3587
rect 15151 3584 15163 3587
rect 16316 3584 16344 3692
rect 18414 3680 18420 3692
rect 18472 3680 18478 3732
rect 18601 3723 18659 3729
rect 18601 3689 18613 3723
rect 18647 3720 18659 3723
rect 18690 3720 18696 3732
rect 18647 3692 18696 3720
rect 18647 3689 18659 3692
rect 18601 3683 18659 3689
rect 18690 3680 18696 3692
rect 18748 3680 18754 3732
rect 18966 3720 18972 3732
rect 18927 3692 18972 3720
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 19334 3680 19340 3732
rect 19392 3720 19398 3732
rect 20901 3723 20959 3729
rect 20901 3720 20913 3723
rect 19392 3692 20913 3720
rect 19392 3680 19398 3692
rect 20901 3689 20913 3692
rect 20947 3689 20959 3723
rect 20901 3683 20959 3689
rect 16752 3655 16810 3661
rect 16752 3621 16764 3655
rect 16798 3652 16810 3655
rect 17586 3652 17592 3664
rect 16798 3624 17592 3652
rect 16798 3621 16810 3624
rect 16752 3615 16810 3621
rect 17586 3612 17592 3624
rect 17644 3612 17650 3664
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 19886 3652 19892 3664
rect 19484 3624 19892 3652
rect 19484 3612 19490 3624
rect 19886 3612 19892 3624
rect 19944 3652 19950 3664
rect 20073 3655 20131 3661
rect 20073 3652 20085 3655
rect 19944 3624 20085 3652
rect 19944 3612 19950 3624
rect 20073 3621 20085 3624
rect 20119 3621 20131 3655
rect 20073 3615 20131 3621
rect 16482 3584 16488 3596
rect 15151 3556 16344 3584
rect 16443 3556 16488 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 18966 3584 18972 3596
rect 16592 3556 18972 3584
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 13044 3488 13277 3516
rect 13044 3476 13050 3488
rect 13265 3485 13277 3488
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 14829 3519 14887 3525
rect 14829 3485 14841 3519
rect 14875 3516 14887 3519
rect 15010 3516 15016 3528
rect 14875 3488 15016 3516
rect 14875 3485 14887 3488
rect 14829 3479 14887 3485
rect 15010 3476 15016 3488
rect 15068 3476 15074 3528
rect 15194 3476 15200 3528
rect 15252 3516 15258 3528
rect 15841 3519 15899 3525
rect 15841 3516 15853 3519
rect 15252 3488 15853 3516
rect 15252 3476 15258 3488
rect 15841 3485 15853 3488
rect 15887 3485 15899 3519
rect 15841 3479 15899 3485
rect 16298 3476 16304 3528
rect 16356 3516 16362 3528
rect 16592 3516 16620 3556
rect 18966 3544 18972 3556
rect 19024 3544 19030 3596
rect 19981 3587 20039 3593
rect 19981 3553 19993 3587
rect 20027 3584 20039 3587
rect 20254 3584 20260 3596
rect 20027 3556 20260 3584
rect 20027 3553 20039 3556
rect 19981 3547 20039 3553
rect 20254 3544 20260 3556
rect 20312 3544 20318 3596
rect 16356 3488 16620 3516
rect 16356 3476 16362 3488
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 19061 3519 19119 3525
rect 19061 3516 19073 3519
rect 18380 3488 19073 3516
rect 18380 3476 18386 3488
rect 19061 3485 19073 3488
rect 19107 3485 19119 3519
rect 19242 3516 19248 3528
rect 19203 3488 19248 3516
rect 19061 3479 19119 3485
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 20165 3519 20223 3525
rect 20165 3485 20177 3519
rect 20211 3485 20223 3519
rect 20165 3479 20223 3485
rect 16114 3448 16120 3460
rect 12728 3420 16120 3448
rect 16114 3408 16120 3420
rect 16172 3408 16178 3460
rect 17770 3408 17776 3460
rect 17828 3448 17834 3460
rect 19613 3451 19671 3457
rect 19613 3448 19625 3451
rect 17828 3420 19625 3448
rect 17828 3408 17834 3420
rect 19613 3417 19625 3420
rect 19659 3417 19671 3451
rect 19613 3411 19671 3417
rect 11054 3380 11060 3392
rect 8588 3352 11060 3380
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 11425 3383 11483 3389
rect 11425 3380 11437 3383
rect 11204 3352 11437 3380
rect 11204 3340 11210 3352
rect 11425 3349 11437 3352
rect 11471 3380 11483 3383
rect 12529 3383 12587 3389
rect 12529 3380 12541 3383
rect 11471 3352 12541 3380
rect 11471 3349 11483 3352
rect 11425 3343 11483 3349
rect 12529 3349 12541 3352
rect 12575 3349 12587 3383
rect 12710 3380 12716 3392
rect 12671 3352 12716 3380
rect 12529 3343 12587 3349
rect 12710 3340 12716 3352
rect 12768 3340 12774 3392
rect 15289 3383 15347 3389
rect 15289 3349 15301 3383
rect 15335 3380 15347 3383
rect 15470 3380 15476 3392
rect 15335 3352 15476 3380
rect 15335 3349 15347 3352
rect 15289 3343 15347 3349
rect 15470 3340 15476 3352
rect 15528 3340 15534 3392
rect 17865 3383 17923 3389
rect 17865 3349 17877 3383
rect 17911 3380 17923 3383
rect 18598 3380 18604 3392
rect 17911 3352 18604 3380
rect 17911 3349 17923 3352
rect 17865 3343 17923 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 18966 3340 18972 3392
rect 19024 3380 19030 3392
rect 20180 3380 20208 3479
rect 19024 3352 20208 3380
rect 19024 3340 19030 3352
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 3050 3136 3056 3188
rect 3108 3176 3114 3188
rect 3145 3179 3203 3185
rect 3145 3176 3157 3179
rect 3108 3148 3157 3176
rect 3108 3136 3114 3148
rect 3145 3145 3157 3148
rect 3191 3145 3203 3179
rect 3145 3139 3203 3145
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 5626 3176 5632 3188
rect 3936 3148 5632 3176
rect 3936 3136 3942 3148
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 5721 3179 5779 3185
rect 5721 3145 5733 3179
rect 5767 3176 5779 3179
rect 6270 3176 6276 3188
rect 5767 3148 6276 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 6840 3148 8064 3176
rect 1578 3068 1584 3120
rect 1636 3108 1642 3120
rect 6840 3108 6868 3148
rect 1636 3080 6868 3108
rect 1636 3068 1642 3080
rect 3234 3000 3240 3052
rect 3292 3040 3298 3052
rect 3602 3040 3608 3052
rect 3292 3012 3608 3040
rect 3292 3000 3298 3012
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 4801 3043 4859 3049
rect 4801 3040 4813 3043
rect 3835 3012 4813 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4801 3009 4813 3012
rect 4847 3040 4859 3043
rect 5258 3040 5264 3052
rect 4847 3012 5264 3040
rect 4847 3009 4859 3012
rect 4801 3003 4859 3009
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 5626 3000 5632 3052
rect 5684 3040 5690 3052
rect 6178 3040 6184 3052
rect 5684 3012 6184 3040
rect 5684 3000 5690 3012
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3040 6423 3043
rect 8036 3040 8064 3148
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 8168 3148 8217 3176
rect 8168 3136 8174 3148
rect 8205 3145 8217 3148
rect 8251 3145 8263 3179
rect 8570 3176 8576 3188
rect 8531 3148 8576 3176
rect 8205 3139 8263 3145
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 9122 3136 9128 3188
rect 9180 3176 9186 3188
rect 9306 3176 9312 3188
rect 9180 3148 9312 3176
rect 9180 3136 9186 3148
rect 9306 3136 9312 3148
rect 9364 3176 9370 3188
rect 15933 3179 15991 3185
rect 15933 3176 15945 3179
rect 9364 3148 15945 3176
rect 9364 3136 9370 3148
rect 15933 3145 15945 3148
rect 15979 3145 15991 3179
rect 15933 3139 15991 3145
rect 16117 3179 16175 3185
rect 16117 3145 16129 3179
rect 16163 3176 16175 3179
rect 20346 3176 20352 3188
rect 16163 3148 20352 3176
rect 16163 3145 16175 3148
rect 16117 3139 16175 3145
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 9674 3108 9680 3120
rect 9048 3080 9680 3108
rect 9048 3049 9076 3080
rect 9674 3068 9680 3080
rect 9732 3068 9738 3120
rect 11977 3111 12035 3117
rect 11977 3077 11989 3111
rect 12023 3108 12035 3111
rect 13446 3108 13452 3120
rect 12023 3080 13452 3108
rect 12023 3077 12035 3080
rect 11977 3071 12035 3077
rect 13446 3068 13452 3080
rect 13504 3068 13510 3120
rect 15378 3068 15384 3120
rect 15436 3108 15442 3120
rect 17313 3111 17371 3117
rect 17313 3108 17325 3111
rect 15436 3080 17325 3108
rect 15436 3068 15442 3080
rect 17313 3077 17325 3080
rect 17359 3077 17371 3111
rect 17313 3071 17371 3077
rect 18690 3068 18696 3120
rect 18748 3108 18754 3120
rect 20901 3111 20959 3117
rect 20901 3108 20913 3111
rect 18748 3080 20913 3108
rect 18748 3068 18754 3080
rect 20901 3077 20913 3080
rect 20947 3077 20959 3111
rect 20901 3071 20959 3077
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 6411 3012 6960 3040
rect 8036 3012 9045 3040
rect 6411 3009 6423 3012
rect 6365 3003 6423 3009
rect 3510 2972 3516 2984
rect 3471 2944 3516 2972
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 4062 2932 4068 2984
rect 4120 2972 4126 2984
rect 4617 2975 4675 2981
rect 4617 2972 4629 2975
rect 4120 2944 4629 2972
rect 4120 2932 4126 2944
rect 4617 2941 4629 2944
rect 4663 2972 4675 2975
rect 5810 2972 5816 2984
rect 4663 2944 5816 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 6086 2972 6092 2984
rect 6047 2944 6092 2972
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 6822 2972 6828 2984
rect 6735 2944 6828 2972
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 6932 2972 6960 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 9217 3003 9275 3009
rect 7098 2981 7104 2984
rect 7092 2972 7104 2981
rect 6932 2944 7104 2972
rect 7092 2935 7104 2944
rect 7156 2972 7162 2984
rect 9232 2972 9260 3003
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 9640 3012 10057 3040
rect 9640 3000 9646 3012
rect 10045 3009 10057 3012
rect 10091 3009 10103 3043
rect 10045 3003 10103 3009
rect 11882 3000 11888 3052
rect 11940 3040 11946 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 11940 3012 13001 3040
rect 11940 3000 11946 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 13078 3000 13084 3052
rect 13136 3040 13142 3052
rect 16577 3043 16635 3049
rect 16577 3040 16589 3043
rect 13136 3012 16589 3040
rect 13136 3000 13142 3012
rect 16577 3009 16589 3012
rect 16623 3009 16635 3043
rect 16577 3003 16635 3009
rect 16761 3043 16819 3049
rect 16761 3009 16773 3043
rect 16807 3040 16819 3043
rect 18598 3040 18604 3052
rect 16807 3012 18604 3040
rect 16807 3009 16819 3012
rect 16761 3003 16819 3009
rect 18598 3000 18604 3012
rect 18656 3040 18662 3052
rect 19245 3043 19303 3049
rect 19245 3040 19257 3043
rect 18656 3012 19257 3040
rect 18656 3000 18662 3012
rect 19245 3009 19257 3012
rect 19291 3009 19303 3043
rect 19245 3003 19303 3009
rect 19334 3000 19340 3052
rect 19392 3040 19398 3052
rect 20257 3043 20315 3049
rect 20257 3040 20269 3043
rect 19392 3012 20269 3040
rect 19392 3000 19398 3012
rect 20257 3009 20269 3012
rect 20303 3009 20315 3043
rect 20257 3003 20315 3009
rect 7156 2944 9260 2972
rect 7098 2932 7104 2935
rect 7156 2932 7162 2944
rect 1118 2864 1124 2916
rect 1176 2904 1182 2916
rect 6840 2904 6868 2932
rect 8386 2904 8392 2916
rect 1176 2876 6776 2904
rect 6840 2876 8392 2904
rect 1176 2864 1182 2876
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 3878 2836 3884 2848
rect 3568 2808 3884 2836
rect 3568 2796 3574 2808
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 4154 2836 4160 2848
rect 4115 2808 4160 2836
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 4338 2796 4344 2848
rect 4396 2836 4402 2848
rect 4525 2839 4583 2845
rect 4525 2836 4537 2839
rect 4396 2808 4537 2836
rect 4396 2796 4402 2808
rect 4525 2805 4537 2808
rect 4571 2805 4583 2839
rect 4525 2799 4583 2805
rect 5350 2796 5356 2848
rect 5408 2836 5414 2848
rect 5994 2836 6000 2848
rect 5408 2808 6000 2836
rect 5408 2796 5414 2808
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 6748 2836 6776 2876
rect 8386 2864 8392 2876
rect 8444 2864 8450 2916
rect 9232 2904 9260 2944
rect 10312 2975 10370 2981
rect 10312 2941 10324 2975
rect 10358 2972 10370 2975
rect 11146 2972 11152 2984
rect 10358 2944 11152 2972
rect 10358 2941 10370 2944
rect 10312 2935 10370 2941
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 11793 2975 11851 2981
rect 11793 2941 11805 2975
rect 11839 2972 11851 2975
rect 12250 2972 12256 2984
rect 11839 2944 12256 2972
rect 11839 2941 11851 2944
rect 11793 2935 11851 2941
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 12360 2944 12664 2972
rect 8864 2876 9168 2904
rect 9232 2876 10456 2904
rect 8864 2836 8892 2876
rect 6748 2808 8892 2836
rect 8938 2796 8944 2848
rect 8996 2836 9002 2848
rect 9140 2836 9168 2876
rect 10428 2848 10456 2876
rect 10778 2864 10784 2916
rect 10836 2904 10842 2916
rect 12360 2904 12388 2944
rect 10836 2876 12388 2904
rect 12636 2904 12664 2944
rect 12802 2932 12808 2984
rect 12860 2972 12866 2984
rect 12860 2944 12905 2972
rect 12860 2932 12866 2944
rect 13170 2932 13176 2984
rect 13228 2972 13234 2984
rect 13449 2975 13507 2981
rect 13449 2972 13461 2975
rect 13228 2944 13461 2972
rect 13228 2932 13234 2944
rect 13449 2941 13461 2944
rect 13495 2941 13507 2975
rect 13722 2972 13728 2984
rect 13683 2944 13728 2972
rect 13449 2935 13507 2941
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 14182 2972 14188 2984
rect 14143 2944 14188 2972
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 14458 2932 14464 2984
rect 14516 2972 14522 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14516 2944 14841 2972
rect 14516 2932 14522 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 15562 2972 15568 2984
rect 15523 2944 15568 2972
rect 14829 2935 14887 2941
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 15933 2975 15991 2981
rect 15933 2941 15945 2975
rect 15979 2972 15991 2975
rect 16485 2975 16543 2981
rect 16485 2972 16497 2975
rect 15979 2944 16497 2972
rect 15979 2941 15991 2944
rect 15933 2935 15991 2941
rect 16485 2941 16497 2944
rect 16531 2941 16543 2975
rect 16485 2935 16543 2941
rect 16666 2932 16672 2984
rect 16724 2972 16730 2984
rect 17129 2975 17187 2981
rect 17129 2972 17141 2975
rect 16724 2944 17141 2972
rect 16724 2932 16730 2944
rect 17129 2941 17141 2944
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 17310 2932 17316 2984
rect 17368 2972 17374 2984
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 17368 2944 18061 2972
rect 17368 2932 17374 2944
rect 18049 2941 18061 2944
rect 18095 2941 18107 2975
rect 20438 2972 20444 2984
rect 18049 2935 18107 2941
rect 18984 2944 20444 2972
rect 12897 2907 12955 2913
rect 12897 2904 12909 2907
rect 12636 2876 12909 2904
rect 10836 2864 10842 2876
rect 12897 2873 12909 2876
rect 12943 2873 12955 2907
rect 12897 2867 12955 2873
rect 15105 2907 15163 2913
rect 15105 2873 15117 2907
rect 15151 2904 15163 2907
rect 16298 2904 16304 2916
rect 15151 2876 16304 2904
rect 15151 2873 15163 2876
rect 15105 2867 15163 2873
rect 16298 2864 16304 2876
rect 16356 2864 16362 2916
rect 9950 2836 9956 2848
rect 8996 2808 9041 2836
rect 9140 2808 9956 2836
rect 8996 2796 9002 2808
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 10410 2796 10416 2848
rect 10468 2836 10474 2848
rect 11425 2839 11483 2845
rect 11425 2836 11437 2839
rect 10468 2808 11437 2836
rect 10468 2796 10474 2808
rect 11425 2805 11437 2808
rect 11471 2805 11483 2839
rect 11425 2799 11483 2805
rect 12437 2839 12495 2845
rect 12437 2805 12449 2839
rect 12483 2836 12495 2839
rect 12802 2836 12808 2848
rect 12483 2808 12808 2836
rect 12483 2805 12495 2808
rect 12437 2799 12495 2805
rect 12802 2796 12808 2808
rect 12860 2796 12866 2848
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 14369 2839 14427 2845
rect 14369 2836 14381 2839
rect 13964 2808 14381 2836
rect 13964 2796 13970 2808
rect 14369 2805 14381 2808
rect 14415 2805 14427 2839
rect 14369 2799 14427 2805
rect 15010 2796 15016 2848
rect 15068 2836 15074 2848
rect 15749 2839 15807 2845
rect 15749 2836 15761 2839
rect 15068 2808 15761 2836
rect 15068 2796 15074 2808
rect 15749 2805 15761 2808
rect 15795 2805 15807 2839
rect 15749 2799 15807 2805
rect 17402 2796 17408 2848
rect 17460 2836 17466 2848
rect 18233 2839 18291 2845
rect 18233 2836 18245 2839
rect 17460 2808 18245 2836
rect 17460 2796 17466 2808
rect 18233 2805 18245 2808
rect 18279 2805 18291 2839
rect 18233 2799 18291 2805
rect 18693 2839 18751 2845
rect 18693 2805 18705 2839
rect 18739 2836 18751 2839
rect 18984 2836 19012 2944
rect 20438 2932 20444 2944
rect 20496 2932 20502 2984
rect 20714 2972 20720 2984
rect 20675 2944 20720 2972
rect 20714 2932 20720 2944
rect 20772 2932 20778 2984
rect 19061 2907 19119 2913
rect 19061 2873 19073 2907
rect 19107 2904 19119 2907
rect 20073 2907 20131 2913
rect 19107 2876 19748 2904
rect 19107 2873 19119 2876
rect 19061 2867 19119 2873
rect 18739 2808 19012 2836
rect 18739 2805 18751 2808
rect 18693 2799 18751 2805
rect 19150 2796 19156 2848
rect 19208 2836 19214 2848
rect 19720 2845 19748 2876
rect 20073 2873 20085 2907
rect 20119 2904 20131 2907
rect 20254 2904 20260 2916
rect 20119 2876 20260 2904
rect 20119 2873 20131 2876
rect 20073 2867 20131 2873
rect 20254 2864 20260 2876
rect 20312 2864 20318 2916
rect 19705 2839 19763 2845
rect 19208 2808 19253 2836
rect 19208 2796 19214 2808
rect 19705 2805 19717 2839
rect 19751 2805 19763 2839
rect 20162 2836 20168 2848
rect 20075 2808 20168 2836
rect 19705 2799 19763 2805
rect 20162 2796 20168 2808
rect 20220 2836 20226 2848
rect 20622 2836 20628 2848
rect 20220 2808 20628 2836
rect 20220 2796 20226 2808
rect 20622 2796 20628 2808
rect 20680 2796 20686 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 4338 2632 4344 2644
rect 3559 2604 4344 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 7558 2592 7564 2644
rect 7616 2632 7622 2644
rect 8113 2635 8171 2641
rect 8113 2632 8125 2635
rect 7616 2604 8125 2632
rect 7616 2592 7622 2604
rect 8113 2601 8125 2604
rect 8159 2601 8171 2635
rect 8113 2595 8171 2601
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 9858 2632 9864 2644
rect 9815 2604 9864 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 10137 2635 10195 2641
rect 10137 2601 10149 2635
rect 10183 2632 10195 2635
rect 10318 2632 10324 2644
rect 10183 2604 10324 2632
rect 10183 2601 10195 2604
rect 10137 2595 10195 2601
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 11333 2635 11391 2641
rect 11333 2601 11345 2635
rect 11379 2632 11391 2635
rect 11606 2632 11612 2644
rect 11379 2604 11612 2632
rect 11379 2601 11391 2604
rect 11333 2595 11391 2601
rect 11606 2592 11612 2604
rect 11664 2592 11670 2644
rect 11701 2635 11759 2641
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 12710 2632 12716 2644
rect 11747 2604 12716 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 19061 2635 19119 2641
rect 19061 2601 19073 2635
rect 19107 2632 19119 2635
rect 19150 2632 19156 2644
rect 19107 2604 19156 2632
rect 19107 2601 19119 2604
rect 19061 2595 19119 2601
rect 19150 2592 19156 2604
rect 19208 2592 19214 2644
rect 8202 2524 8208 2576
rect 8260 2524 8266 2576
rect 10229 2567 10287 2573
rect 10229 2533 10241 2567
rect 10275 2564 10287 2567
rect 10594 2564 10600 2576
rect 10275 2536 10600 2564
rect 10275 2533 10287 2536
rect 10229 2527 10287 2533
rect 10594 2524 10600 2536
rect 10652 2524 10658 2576
rect 11793 2567 11851 2573
rect 11793 2533 11805 2567
rect 11839 2564 11851 2567
rect 12158 2564 12164 2576
rect 11839 2536 12164 2564
rect 11839 2533 11851 2536
rect 11793 2527 11851 2533
rect 12158 2524 12164 2536
rect 12216 2524 12222 2576
rect 12250 2524 12256 2576
rect 12308 2564 12314 2576
rect 12897 2567 12955 2573
rect 12897 2564 12909 2567
rect 12308 2536 12909 2564
rect 12308 2524 12314 2536
rect 12897 2533 12909 2536
rect 12943 2533 12955 2567
rect 12897 2527 12955 2533
rect 13633 2567 13691 2573
rect 13633 2533 13645 2567
rect 13679 2564 13691 2567
rect 15749 2567 15807 2573
rect 13679 2536 14872 2564
rect 13679 2533 13691 2536
rect 13633 2527 13691 2533
rect 8220 2496 8248 2524
rect 8849 2499 8907 2505
rect 8220 2468 8340 2496
rect 8312 2437 8340 2468
rect 8849 2465 8861 2499
rect 8895 2465 8907 2499
rect 8849 2459 8907 2465
rect 10781 2499 10839 2505
rect 10781 2465 10793 2499
rect 10827 2496 10839 2499
rect 12434 2496 12440 2508
rect 10827 2468 12440 2496
rect 10827 2465 10839 2468
rect 10781 2459 10839 2465
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 8220 2360 8248 2391
rect 8478 2360 8484 2372
rect 8220 2332 8484 2360
rect 8478 2320 8484 2332
rect 8536 2320 8542 2372
rect 7745 2295 7803 2301
rect 7745 2261 7757 2295
rect 7791 2292 7803 2295
rect 8864 2292 8892 2459
rect 12434 2456 12440 2468
rect 12492 2456 12498 2508
rect 12710 2505 12716 2508
rect 12652 2499 12716 2505
rect 12652 2465 12664 2499
rect 12698 2465 12716 2499
rect 12652 2459 12716 2465
rect 12710 2456 12716 2459
rect 12768 2456 12774 2508
rect 13265 2499 13323 2505
rect 13265 2465 13277 2499
rect 13311 2496 13323 2499
rect 13357 2499 13415 2505
rect 13357 2496 13369 2499
rect 13311 2468 13369 2496
rect 13311 2465 13323 2468
rect 13265 2459 13323 2465
rect 13357 2465 13369 2468
rect 13403 2465 13415 2499
rect 13357 2459 13415 2465
rect 13998 2456 14004 2508
rect 14056 2496 14062 2508
rect 14844 2505 14872 2536
rect 15749 2533 15761 2567
rect 15795 2564 15807 2567
rect 17310 2564 17316 2576
rect 15795 2536 17316 2564
rect 15795 2533 15807 2536
rect 15749 2527 15807 2533
rect 17310 2524 17316 2536
rect 17368 2524 17374 2576
rect 18874 2524 18880 2576
rect 18932 2564 18938 2576
rect 20441 2567 20499 2573
rect 20441 2564 20453 2567
rect 18932 2536 20453 2564
rect 18932 2524 18938 2536
rect 20441 2533 20453 2536
rect 20487 2533 20499 2567
rect 20441 2527 20499 2533
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 14056 2468 14105 2496
rect 14056 2456 14062 2468
rect 14093 2465 14105 2468
rect 14139 2465 14151 2499
rect 14093 2459 14151 2465
rect 14829 2499 14887 2505
rect 14829 2465 14841 2499
rect 14875 2465 14887 2499
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 14829 2459 14887 2465
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 16206 2496 16212 2508
rect 16167 2468 16212 2496
rect 16206 2456 16212 2468
rect 16264 2456 16270 2508
rect 16298 2456 16304 2508
rect 16356 2496 16362 2508
rect 16945 2499 17003 2505
rect 16945 2496 16957 2499
rect 16356 2468 16957 2496
rect 16356 2456 16362 2468
rect 16945 2465 16957 2468
rect 16991 2465 17003 2499
rect 16945 2459 17003 2465
rect 17497 2499 17555 2505
rect 17497 2465 17509 2499
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2496 18383 2499
rect 18506 2496 18512 2508
rect 18371 2468 18512 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 10410 2428 10416 2440
rect 10371 2400 10416 2428
rect 9125 2391 9183 2397
rect 9140 2360 9168 2391
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 10870 2388 10876 2440
rect 10928 2428 10934 2440
rect 11149 2431 11207 2437
rect 11149 2428 11161 2431
rect 10928 2400 11161 2428
rect 10928 2388 10934 2400
rect 11149 2397 11161 2400
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11756 2400 11897 2428
rect 11756 2388 11762 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2428 14427 2431
rect 15562 2428 15568 2440
rect 14415 2400 15568 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 16485 2431 16543 2437
rect 16485 2397 16497 2431
rect 16531 2428 16543 2431
rect 17512 2428 17540 2459
rect 18506 2456 18512 2468
rect 18564 2456 18570 2508
rect 19426 2496 19432 2508
rect 19387 2468 19432 2496
rect 19426 2456 19432 2468
rect 19484 2456 19490 2508
rect 20070 2456 20076 2508
rect 20128 2496 20134 2508
rect 20165 2499 20223 2505
rect 20165 2496 20177 2499
rect 20128 2468 20177 2496
rect 20128 2456 20134 2468
rect 20165 2465 20177 2468
rect 20211 2465 20223 2499
rect 20165 2459 20223 2465
rect 16531 2400 17540 2428
rect 16531 2397 16543 2400
rect 16485 2391 16543 2397
rect 17862 2388 17868 2440
rect 17920 2428 17926 2440
rect 19242 2428 19248 2440
rect 17920 2400 19248 2428
rect 17920 2388 17926 2400
rect 19242 2388 19248 2400
rect 19300 2428 19306 2440
rect 19521 2431 19579 2437
rect 19521 2428 19533 2431
rect 19300 2400 19533 2428
rect 19300 2388 19306 2400
rect 19521 2397 19533 2400
rect 19567 2397 19579 2431
rect 19521 2391 19579 2397
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 14182 2360 14188 2372
rect 9140 2332 14188 2360
rect 14182 2320 14188 2332
rect 14240 2320 14246 2372
rect 19334 2320 19340 2372
rect 19392 2360 19398 2372
rect 19628 2360 19656 2391
rect 19392 2332 19656 2360
rect 19392 2320 19398 2332
rect 10962 2292 10968 2304
rect 7791 2264 8892 2292
rect 10923 2264 10968 2292
rect 7791 2261 7803 2264
rect 7745 2255 7803 2261
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11149 2295 11207 2301
rect 11149 2261 11161 2295
rect 11195 2292 11207 2295
rect 13265 2295 13323 2301
rect 13265 2292 13277 2295
rect 11195 2264 13277 2292
rect 11195 2261 11207 2264
rect 11149 2255 11207 2261
rect 13265 2261 13277 2264
rect 13311 2261 13323 2295
rect 13265 2255 13323 2261
rect 14458 2252 14464 2304
rect 14516 2292 14522 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14516 2264 15025 2292
rect 14516 2252 14522 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17129 2295 17187 2301
rect 17129 2292 17141 2295
rect 16816 2264 17141 2292
rect 16816 2252 16822 2264
rect 17129 2261 17141 2264
rect 17175 2261 17187 2295
rect 17129 2255 17187 2261
rect 17681 2295 17739 2301
rect 17681 2261 17693 2295
rect 17727 2292 17739 2295
rect 17770 2292 17776 2304
rect 17727 2264 17776 2292
rect 17727 2261 17739 2264
rect 17681 2255 17739 2261
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 18506 2292 18512 2304
rect 18467 2264 18512 2292
rect 18506 2252 18512 2264
rect 18564 2252 18570 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 2498 2048 2504 2100
rect 2556 2088 2562 2100
rect 8938 2088 8944 2100
rect 2556 2060 8944 2088
rect 2556 2048 2562 2060
rect 8938 2048 8944 2060
rect 8996 2048 9002 2100
rect 10962 2048 10968 2100
rect 11020 2088 11026 2100
rect 22002 2088 22008 2100
rect 11020 2060 22008 2088
rect 11020 2048 11026 2060
rect 22002 2048 22008 2060
rect 22060 2048 22066 2100
rect 8202 1980 8208 2032
rect 8260 2020 8266 2032
rect 8662 2020 8668 2032
rect 8260 1992 8668 2020
rect 8260 1980 8266 1992
rect 8662 1980 8668 1992
rect 8720 1980 8726 2032
rect 11698 1980 11704 2032
rect 11756 2020 11762 2032
rect 11974 2020 11980 2032
rect 11756 1992 11980 2020
rect 11756 1980 11762 1992
rect 11974 1980 11980 1992
rect 12032 1980 12038 2032
rect 2038 1368 2044 1420
rect 2096 1408 2102 1420
rect 7190 1408 7196 1420
rect 2096 1380 7196 1408
rect 2096 1368 2102 1380
rect 7190 1368 7196 1380
rect 7248 1368 7254 1420
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 18696 19499 18748 19508
rect 18696 19465 18705 19499
rect 18705 19465 18739 19499
rect 18739 19465 18748 19499
rect 18696 19456 18748 19465
rect 20720 19499 20772 19508
rect 20720 19465 20729 19499
rect 20729 19465 20763 19499
rect 20763 19465 20772 19499
rect 20720 19456 20772 19465
rect 3424 19252 3476 19304
rect 17868 19252 17920 19304
rect 20536 19295 20588 19304
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 6736 19184 6788 19236
rect 2780 19116 2832 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1952 18955 2004 18964
rect 1952 18921 1961 18955
rect 1961 18921 1995 18955
rect 1995 18921 2004 18955
rect 1952 18912 2004 18921
rect 17868 18887 17920 18896
rect 17868 18853 17877 18887
rect 17877 18853 17911 18887
rect 17911 18853 17920 18887
rect 17868 18844 17920 18853
rect 6184 18776 6236 18828
rect 16672 18776 16724 18828
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 20720 18411 20772 18420
rect 20720 18377 20729 18411
rect 20729 18377 20763 18411
rect 20763 18377 20772 18411
rect 20720 18368 20772 18377
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 20536 18207 20588 18216
rect 20536 18173 20545 18207
rect 20545 18173 20579 18207
rect 20579 18173 20588 18207
rect 20536 18164 20588 18173
rect 16580 18096 16632 18148
rect 18972 18096 19024 18148
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1768 17756 1820 17808
rect 20536 17756 20588 17808
rect 6368 17688 6420 17740
rect 17132 17688 17184 17740
rect 7380 17620 7432 17672
rect 1676 17552 1728 17604
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 20168 17323 20220 17332
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 20720 17323 20772 17332
rect 20720 17289 20729 17323
rect 20729 17289 20763 17323
rect 20763 17289 20772 17323
rect 20720 17280 20772 17289
rect 7196 17076 7248 17128
rect 19340 17076 19392 17128
rect 20168 17076 20220 17128
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1860 16736 1912 16788
rect 20444 16779 20496 16788
rect 20444 16745 20453 16779
rect 20453 16745 20487 16779
rect 20487 16745 20496 16779
rect 20444 16736 20496 16745
rect 5816 16600 5868 16652
rect 20628 16600 20680 16652
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 3700 16235 3752 16244
rect 3700 16201 3709 16235
rect 3709 16201 3743 16235
rect 3743 16201 3752 16235
rect 3700 16192 3752 16201
rect 17960 16192 18012 16244
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 3240 15988 3292 16040
rect 3516 16031 3568 16040
rect 3516 15997 3525 16031
rect 3525 15997 3559 16031
rect 3559 15997 3568 16031
rect 3516 15988 3568 15997
rect 13728 15988 13780 16040
rect 20536 16031 20588 16040
rect 20536 15997 20545 16031
rect 20545 15997 20579 16031
rect 20579 15997 20588 16031
rect 20536 15988 20588 15997
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 2504 15691 2556 15700
rect 2504 15657 2513 15691
rect 2513 15657 2547 15691
rect 2547 15657 2556 15691
rect 2504 15648 2556 15657
rect 19892 15691 19944 15700
rect 19892 15657 19901 15691
rect 19901 15657 19935 15691
rect 19935 15657 19944 15691
rect 19892 15648 19944 15657
rect 20260 15648 20312 15700
rect 3516 15580 3568 15632
rect 13728 15623 13780 15632
rect 13728 15589 13737 15623
rect 13737 15589 13771 15623
rect 13771 15589 13780 15623
rect 13728 15580 13780 15589
rect 1860 15512 1912 15564
rect 3976 15512 4028 15564
rect 4252 15512 4304 15564
rect 13268 15512 13320 15564
rect 19432 15512 19484 15564
rect 19800 15512 19852 15564
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 2780 15104 2832 15156
rect 3056 15147 3108 15156
rect 3056 15113 3065 15147
rect 3065 15113 3099 15147
rect 3099 15113 3108 15147
rect 3056 15104 3108 15113
rect 3608 15147 3660 15156
rect 3608 15113 3617 15147
rect 3617 15113 3651 15147
rect 3651 15113 3660 15147
rect 3608 15104 3660 15113
rect 4068 15104 4120 15156
rect 20352 15104 20404 15156
rect 1952 15079 2004 15088
rect 1952 15045 1961 15079
rect 1961 15045 1995 15079
rect 1995 15045 2004 15079
rect 1952 15036 2004 15045
rect 17960 15036 18012 15088
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 5632 14968 5684 15020
rect 7564 14968 7616 15020
rect 14372 14968 14424 15020
rect 6000 14943 6052 14952
rect 6000 14909 6009 14943
rect 6009 14909 6043 14943
rect 6043 14909 6052 14943
rect 6000 14900 6052 14909
rect 11612 14943 11664 14952
rect 11612 14909 11621 14943
rect 11621 14909 11655 14943
rect 11655 14909 11664 14943
rect 11612 14900 11664 14909
rect 14464 14900 14516 14952
rect 19340 14900 19392 14952
rect 19708 14900 19760 14952
rect 20444 14900 20496 14952
rect 5356 14832 5408 14884
rect 17040 14832 17092 14884
rect 13636 14807 13688 14816
rect 13636 14773 13645 14807
rect 13645 14773 13679 14807
rect 13679 14773 13688 14807
rect 13636 14764 13688 14773
rect 14004 14807 14056 14816
rect 14004 14773 14013 14807
rect 14013 14773 14047 14807
rect 14047 14773 14056 14807
rect 14004 14764 14056 14773
rect 16948 14807 17000 14816
rect 16948 14773 16957 14807
rect 16957 14773 16991 14807
rect 16991 14773 17000 14807
rect 16948 14764 17000 14773
rect 19248 14764 19300 14816
rect 20260 14764 20312 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 7656 14560 7708 14612
rect 16580 14560 16632 14612
rect 19892 14603 19944 14612
rect 1768 14492 1820 14544
rect 3056 14492 3108 14544
rect 3148 14492 3200 14544
rect 6000 14492 6052 14544
rect 7748 14492 7800 14544
rect 11152 14492 11204 14544
rect 19892 14569 19901 14603
rect 19901 14569 19935 14603
rect 19935 14569 19944 14603
rect 19892 14560 19944 14569
rect 19984 14560 20036 14612
rect 20352 14560 20404 14612
rect 17592 14492 17644 14544
rect 2872 14424 2924 14476
rect 4896 14424 4948 14476
rect 7012 14424 7064 14476
rect 10692 14467 10744 14476
rect 10692 14433 10701 14467
rect 10701 14433 10735 14467
rect 10735 14433 10744 14467
rect 10692 14424 10744 14433
rect 12440 14424 12492 14476
rect 10784 14399 10836 14408
rect 2688 14288 2740 14340
rect 2228 14220 2280 14272
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 15108 14424 15160 14476
rect 16396 14467 16448 14476
rect 16396 14433 16430 14467
rect 16430 14433 16448 14467
rect 16396 14424 16448 14433
rect 19984 14424 20036 14476
rect 10048 14288 10100 14340
rect 15384 14356 15436 14408
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 18972 14356 19024 14408
rect 20352 14424 20404 14476
rect 19892 14288 19944 14340
rect 20168 14288 20220 14340
rect 8668 14220 8720 14272
rect 10324 14263 10376 14272
rect 10324 14229 10333 14263
rect 10333 14229 10367 14263
rect 10367 14229 10376 14263
rect 10324 14220 10376 14229
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 18512 14220 18564 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 2780 14016 2832 14068
rect 6276 14016 6328 14068
rect 7012 14059 7064 14068
rect 7012 14025 7021 14059
rect 7021 14025 7055 14059
rect 7055 14025 7064 14059
rect 7012 14016 7064 14025
rect 16396 14016 16448 14068
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 1768 13812 1820 13864
rect 4068 13880 4120 13932
rect 7656 13923 7708 13932
rect 7656 13889 7665 13923
rect 7665 13889 7699 13923
rect 7699 13889 7708 13923
rect 7656 13880 7708 13889
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 4160 13812 4212 13864
rect 7564 13812 7616 13864
rect 4068 13744 4120 13796
rect 5724 13744 5776 13796
rect 7012 13744 7064 13796
rect 10324 13812 10376 13864
rect 11244 13812 11296 13864
rect 11612 13923 11664 13932
rect 11612 13889 11621 13923
rect 11621 13889 11655 13923
rect 11655 13889 11664 13923
rect 11612 13880 11664 13889
rect 14004 13880 14056 13932
rect 17592 13923 17644 13932
rect 17592 13889 17601 13923
rect 17601 13889 17635 13923
rect 17635 13889 17644 13923
rect 17592 13880 17644 13889
rect 12440 13812 12492 13864
rect 14372 13812 14424 13864
rect 15384 13812 15436 13864
rect 15936 13812 15988 13864
rect 18788 13812 18840 13864
rect 20720 13948 20772 14000
rect 19708 13923 19760 13932
rect 19708 13889 19717 13923
rect 19717 13889 19751 13923
rect 19751 13889 19760 13923
rect 19708 13880 19760 13889
rect 20444 13923 20496 13932
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 19248 13812 19300 13864
rect 4344 13719 4396 13728
rect 4344 13685 4353 13719
rect 4353 13685 4387 13719
rect 4387 13685 4396 13719
rect 4344 13676 4396 13685
rect 4620 13719 4672 13728
rect 4620 13685 4629 13719
rect 4629 13685 4663 13719
rect 4663 13685 4672 13719
rect 4620 13676 4672 13685
rect 5080 13719 5132 13728
rect 5080 13685 5089 13719
rect 5089 13685 5123 13719
rect 5123 13685 5132 13719
rect 5080 13676 5132 13685
rect 6644 13676 6696 13728
rect 7472 13719 7524 13728
rect 7472 13685 7481 13719
rect 7481 13685 7515 13719
rect 7515 13685 7524 13719
rect 14188 13719 14240 13728
rect 7472 13676 7524 13685
rect 14188 13685 14197 13719
rect 14197 13685 14231 13719
rect 14231 13685 14240 13719
rect 14188 13676 14240 13685
rect 16764 13676 16816 13728
rect 17408 13719 17460 13728
rect 17408 13685 17417 13719
rect 17417 13685 17451 13719
rect 17451 13685 17460 13719
rect 17960 13744 18012 13796
rect 17408 13676 17460 13685
rect 18880 13676 18932 13728
rect 19156 13719 19208 13728
rect 19156 13685 19165 13719
rect 19165 13685 19199 13719
rect 19199 13685 19208 13719
rect 19156 13676 19208 13685
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 2872 13472 2924 13524
rect 4620 13472 4672 13524
rect 6644 13515 6696 13524
rect 6644 13481 6653 13515
rect 6653 13481 6687 13515
rect 6687 13481 6696 13515
rect 6644 13472 6696 13481
rect 7012 13515 7064 13524
rect 7012 13481 7021 13515
rect 7021 13481 7055 13515
rect 7055 13481 7064 13515
rect 7012 13472 7064 13481
rect 7472 13472 7524 13524
rect 10968 13472 11020 13524
rect 11244 13472 11296 13524
rect 13636 13472 13688 13524
rect 3516 13404 3568 13456
rect 4344 13404 4396 13456
rect 8208 13404 8260 13456
rect 8300 13404 8352 13456
rect 12808 13404 12860 13456
rect 12992 13447 13044 13456
rect 12992 13413 13001 13447
rect 13001 13413 13035 13447
rect 13035 13413 13044 13447
rect 12992 13404 13044 13413
rect 13452 13404 13504 13456
rect 14188 13404 14240 13456
rect 16764 13472 16816 13524
rect 16948 13515 17000 13524
rect 16948 13481 16957 13515
rect 16957 13481 16991 13515
rect 16991 13481 17000 13515
rect 16948 13472 17000 13481
rect 17040 13515 17092 13524
rect 17040 13481 17049 13515
rect 17049 13481 17083 13515
rect 17083 13481 17092 13515
rect 17040 13472 17092 13481
rect 18880 13472 18932 13524
rect 17408 13404 17460 13456
rect 18512 13404 18564 13456
rect 2044 13336 2096 13388
rect 2320 13268 2372 13320
rect 2596 13311 2648 13320
rect 2596 13277 2605 13311
rect 2605 13277 2639 13311
rect 2639 13277 2648 13311
rect 2596 13268 2648 13277
rect 8760 13336 8812 13388
rect 10048 13379 10100 13388
rect 10048 13345 10082 13379
rect 10082 13345 10100 13379
rect 11796 13379 11848 13388
rect 10048 13336 10100 13345
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4160 13268 4212 13277
rect 7748 13268 7800 13320
rect 8668 13268 8720 13320
rect 11796 13345 11805 13379
rect 11805 13345 11839 13379
rect 11839 13345 11848 13379
rect 11796 13336 11848 13345
rect 12900 13336 12952 13388
rect 12440 13268 12492 13320
rect 15292 13336 15344 13388
rect 16304 13336 16356 13388
rect 20168 13379 20220 13388
rect 20168 13345 20177 13379
rect 20177 13345 20211 13379
rect 20211 13345 20220 13379
rect 20168 13336 20220 13345
rect 3332 13200 3384 13252
rect 7012 13200 7064 13252
rect 16396 13268 16448 13320
rect 13452 13200 13504 13252
rect 17776 13268 17828 13320
rect 2136 13132 2188 13184
rect 5540 13175 5592 13184
rect 5540 13141 5549 13175
rect 5549 13141 5583 13175
rect 5583 13141 5592 13175
rect 5540 13132 5592 13141
rect 6092 13132 6144 13184
rect 11152 13132 11204 13184
rect 14280 13132 14332 13184
rect 14924 13175 14976 13184
rect 14924 13141 14933 13175
rect 14933 13141 14967 13175
rect 14967 13141 14976 13175
rect 14924 13132 14976 13141
rect 16764 13132 16816 13184
rect 17132 13132 17184 13184
rect 20352 13311 20404 13320
rect 20352 13277 20361 13311
rect 20361 13277 20395 13311
rect 20395 13277 20404 13311
rect 20352 13268 20404 13277
rect 18604 13132 18656 13184
rect 19156 13132 19208 13184
rect 19340 13132 19392 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 2044 12928 2096 12980
rect 2228 12835 2280 12844
rect 2228 12801 2237 12835
rect 2237 12801 2271 12835
rect 2271 12801 2280 12835
rect 2228 12792 2280 12801
rect 4068 12928 4120 12980
rect 5080 12928 5132 12980
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 7748 12928 7800 12980
rect 10048 12971 10100 12980
rect 10048 12937 10057 12971
rect 10057 12937 10091 12971
rect 10091 12937 10100 12971
rect 10048 12928 10100 12937
rect 17960 12928 18012 12980
rect 18880 12928 18932 12980
rect 6460 12792 6512 12844
rect 8668 12835 8720 12844
rect 8668 12801 8677 12835
rect 8677 12801 8711 12835
rect 8711 12801 8720 12835
rect 8668 12792 8720 12801
rect 10416 12792 10468 12844
rect 13452 12835 13504 12844
rect 13452 12801 13461 12835
rect 13461 12801 13495 12835
rect 13495 12801 13504 12835
rect 13452 12792 13504 12801
rect 16488 12860 16540 12912
rect 14924 12792 14976 12844
rect 2136 12767 2188 12776
rect 2136 12733 2145 12767
rect 2145 12733 2179 12767
rect 2179 12733 2188 12767
rect 2136 12724 2188 12733
rect 2872 12724 2924 12776
rect 4160 12724 4212 12776
rect 5264 12724 5316 12776
rect 6092 12767 6144 12776
rect 6092 12733 6101 12767
rect 6101 12733 6135 12767
rect 6135 12733 6144 12767
rect 6092 12724 6144 12733
rect 6644 12724 6696 12776
rect 10968 12767 11020 12776
rect 2596 12588 2648 12640
rect 4068 12656 4120 12708
rect 7288 12656 7340 12708
rect 10232 12656 10284 12708
rect 10968 12733 11002 12767
rect 11002 12733 11020 12767
rect 10968 12724 11020 12733
rect 13912 12724 13964 12776
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 12900 12656 12952 12708
rect 15384 12656 15436 12708
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 7748 12588 7800 12640
rect 8484 12588 8536 12640
rect 13176 12588 13228 12640
rect 13820 12588 13872 12640
rect 15108 12588 15160 12640
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 18604 12724 18656 12776
rect 19156 12767 19208 12776
rect 19156 12733 19190 12767
rect 19190 12733 19208 12767
rect 19156 12724 19208 12733
rect 20352 12928 20404 12980
rect 20720 12835 20772 12844
rect 20720 12801 20729 12835
rect 20729 12801 20763 12835
rect 20763 12801 20772 12835
rect 20720 12792 20772 12801
rect 20444 12724 20496 12776
rect 17592 12656 17644 12708
rect 17316 12631 17368 12640
rect 17316 12597 17325 12631
rect 17325 12597 17359 12631
rect 17359 12597 17368 12631
rect 17316 12588 17368 12597
rect 17408 12631 17460 12640
rect 17408 12597 17417 12631
rect 17417 12597 17451 12631
rect 17451 12597 17460 12631
rect 18696 12656 18748 12708
rect 17408 12588 17460 12597
rect 20720 12588 20772 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 1676 12427 1728 12436
rect 1676 12393 1685 12427
rect 1685 12393 1719 12427
rect 1719 12393 1728 12427
rect 1676 12384 1728 12393
rect 3056 12384 3108 12436
rect 3700 12384 3752 12436
rect 2504 12359 2556 12368
rect 2504 12325 2513 12359
rect 2513 12325 2547 12359
rect 2547 12325 2556 12359
rect 3332 12359 3384 12368
rect 2504 12316 2556 12325
rect 1860 12248 1912 12300
rect 3056 12291 3108 12300
rect 3056 12257 3065 12291
rect 3065 12257 3099 12291
rect 3099 12257 3108 12291
rect 3056 12248 3108 12257
rect 3332 12325 3341 12359
rect 3341 12325 3375 12359
rect 3375 12325 3384 12359
rect 3332 12316 3384 12325
rect 4160 12384 4212 12436
rect 4528 12384 4580 12436
rect 6460 12427 6512 12436
rect 4344 12248 4396 12300
rect 5172 12316 5224 12368
rect 6460 12393 6469 12427
rect 6469 12393 6503 12427
rect 6503 12393 6512 12427
rect 6460 12384 6512 12393
rect 7012 12384 7064 12436
rect 8208 12384 8260 12436
rect 8484 12384 8536 12436
rect 10784 12384 10836 12436
rect 13820 12384 13872 12436
rect 16488 12384 16540 12436
rect 18052 12384 18104 12436
rect 18144 12384 18196 12436
rect 19984 12384 20036 12436
rect 20628 12384 20680 12436
rect 9220 12316 9272 12368
rect 10600 12316 10652 12368
rect 14832 12316 14884 12368
rect 17132 12316 17184 12368
rect 6460 12248 6512 12300
rect 7380 12248 7432 12300
rect 8392 12291 8444 12300
rect 8392 12257 8401 12291
rect 8401 12257 8435 12291
rect 8435 12257 8444 12291
rect 8392 12248 8444 12257
rect 8484 12248 8536 12300
rect 8668 12248 8720 12300
rect 8944 12248 8996 12300
rect 3240 12180 3292 12232
rect 4712 12223 4764 12232
rect 2780 12112 2832 12164
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 5080 12223 5132 12232
rect 5080 12189 5089 12223
rect 5089 12189 5123 12223
rect 5123 12189 5132 12223
rect 5080 12180 5132 12189
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7288 12180 7340 12189
rect 8208 12180 8260 12232
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 4804 12112 4856 12164
rect 12072 12248 12124 12300
rect 12716 12248 12768 12300
rect 14372 12248 14424 12300
rect 9404 12180 9456 12232
rect 10048 12180 10100 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 11152 12223 11204 12232
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 12624 12180 12676 12232
rect 13176 12223 13228 12232
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 13452 12180 13504 12232
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14648 12180 14700 12189
rect 16028 12248 16080 12300
rect 16948 12248 17000 12300
rect 15292 12180 15344 12232
rect 3424 12044 3476 12096
rect 3608 12044 3660 12096
rect 3792 12044 3844 12096
rect 4988 12044 5040 12096
rect 5264 12044 5316 12096
rect 11796 12112 11848 12164
rect 16212 12180 16264 12232
rect 17408 12180 17460 12232
rect 18512 12316 18564 12368
rect 17960 12248 18012 12300
rect 19156 12248 19208 12300
rect 18880 12223 18932 12232
rect 8852 12087 8904 12096
rect 8852 12053 8861 12087
rect 8861 12053 8895 12087
rect 8895 12053 8904 12087
rect 8852 12044 8904 12053
rect 10232 12044 10284 12096
rect 11060 12044 11112 12096
rect 16488 12112 16540 12164
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 19800 12112 19852 12164
rect 12348 12044 12400 12096
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 13084 12044 13136 12096
rect 15752 12044 15804 12096
rect 17224 12044 17276 12096
rect 19432 12087 19484 12096
rect 19432 12053 19441 12087
rect 19441 12053 19475 12087
rect 19475 12053 19484 12087
rect 19432 12044 19484 12053
rect 19524 12044 19576 12096
rect 20536 12180 20588 12232
rect 20444 12112 20496 12164
rect 20904 12044 20956 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 3976 11840 4028 11892
rect 4712 11883 4764 11892
rect 3332 11772 3384 11824
rect 4712 11849 4721 11883
rect 4721 11849 4755 11883
rect 4755 11849 4764 11883
rect 4712 11840 4764 11849
rect 8208 11840 8260 11892
rect 8576 11840 8628 11892
rect 8760 11883 8812 11892
rect 8760 11849 8769 11883
rect 8769 11849 8803 11883
rect 8803 11849 8812 11883
rect 8760 11840 8812 11849
rect 9036 11840 9088 11892
rect 10508 11840 10560 11892
rect 10692 11883 10744 11892
rect 10692 11849 10701 11883
rect 10701 11849 10735 11883
rect 10735 11849 10744 11883
rect 10692 11840 10744 11849
rect 11152 11840 11204 11892
rect 11796 11840 11848 11892
rect 10600 11772 10652 11824
rect 11060 11772 11112 11824
rect 13360 11840 13412 11892
rect 15292 11883 15344 11892
rect 15292 11849 15301 11883
rect 15301 11849 15335 11883
rect 15335 11849 15344 11883
rect 15292 11840 15344 11849
rect 15660 11840 15712 11892
rect 16212 11840 16264 11892
rect 16488 11840 16540 11892
rect 17960 11840 18012 11892
rect 20536 11840 20588 11892
rect 2596 11747 2648 11756
rect 2596 11713 2605 11747
rect 2605 11713 2639 11747
rect 2639 11713 2648 11747
rect 2596 11704 2648 11713
rect 2780 11704 2832 11756
rect 5540 11704 5592 11756
rect 7104 11747 7156 11756
rect 7104 11713 7113 11747
rect 7113 11713 7147 11747
rect 7147 11713 7156 11747
rect 7104 11704 7156 11713
rect 8576 11704 8628 11756
rect 17408 11772 17460 11824
rect 18144 11772 18196 11824
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 13452 11704 13504 11756
rect 14372 11704 14424 11756
rect 14648 11704 14700 11756
rect 15200 11704 15252 11756
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 18512 11704 18564 11756
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 2964 11636 3016 11688
rect 3148 11636 3200 11688
rect 4068 11636 4120 11688
rect 9036 11636 9088 11688
rect 9956 11636 10008 11688
rect 10968 11636 11020 11688
rect 11704 11636 11756 11688
rect 2872 11568 2924 11620
rect 3240 11568 3292 11620
rect 5356 11568 5408 11620
rect 5816 11568 5868 11620
rect 3792 11500 3844 11552
rect 5264 11500 5316 11552
rect 7104 11500 7156 11552
rect 8392 11500 8444 11552
rect 10784 11500 10836 11552
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 12900 11500 12952 11552
rect 14096 11500 14148 11552
rect 15016 11500 15068 11552
rect 15660 11543 15712 11552
rect 15660 11509 15669 11543
rect 15669 11509 15703 11543
rect 15703 11509 15712 11543
rect 15660 11500 15712 11509
rect 16396 11636 16448 11688
rect 18880 11636 18932 11688
rect 19708 11636 19760 11688
rect 20260 11636 20312 11688
rect 16580 11611 16632 11620
rect 16580 11577 16614 11611
rect 16614 11577 16632 11611
rect 16580 11568 16632 11577
rect 16856 11568 16908 11620
rect 18972 11568 19024 11620
rect 16488 11500 16540 11552
rect 17040 11500 17092 11552
rect 19432 11500 19484 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 3056 11296 3108 11348
rect 5264 11339 5316 11348
rect 5264 11305 5273 11339
rect 5273 11305 5307 11339
rect 5307 11305 5316 11339
rect 5264 11296 5316 11305
rect 6368 11296 6420 11348
rect 7564 11296 7616 11348
rect 10968 11296 11020 11348
rect 1400 11228 1452 11280
rect 4160 11228 4212 11280
rect 9128 11228 9180 11280
rect 10876 11228 10928 11280
rect 11152 11228 11204 11280
rect 12992 11296 13044 11348
rect 13452 11296 13504 11348
rect 13912 11296 13964 11348
rect 1860 11160 1912 11212
rect 2872 11160 2924 11212
rect 3056 11203 3108 11212
rect 3056 11169 3065 11203
rect 3065 11169 3099 11203
rect 3099 11169 3108 11203
rect 3056 11160 3108 11169
rect 5540 11160 5592 11212
rect 6828 11203 6880 11212
rect 6828 11169 6837 11203
rect 6837 11169 6871 11203
rect 6871 11169 6880 11203
rect 6828 11160 6880 11169
rect 7288 11160 7340 11212
rect 8208 11160 8260 11212
rect 9680 11160 9732 11212
rect 3240 11092 3292 11144
rect 2504 11024 2556 11076
rect 2780 11024 2832 11076
rect 4804 11067 4856 11076
rect 4804 11033 4813 11067
rect 4813 11033 4847 11067
rect 4847 11033 4856 11067
rect 4804 11024 4856 11033
rect 5632 11092 5684 11144
rect 5816 11092 5868 11144
rect 6920 11135 6972 11144
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 7564 11092 7616 11144
rect 9772 11092 9824 11144
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 10508 11092 10560 11144
rect 12440 11160 12492 11212
rect 12716 11160 12768 11212
rect 16764 11296 16816 11348
rect 16856 11296 16908 11348
rect 19524 11339 19576 11348
rect 19524 11305 19533 11339
rect 19533 11305 19567 11339
rect 19567 11305 19576 11339
rect 19524 11296 19576 11305
rect 20352 11296 20404 11348
rect 20904 11339 20956 11348
rect 20904 11305 20913 11339
rect 20913 11305 20947 11339
rect 20947 11305 20956 11339
rect 20904 11296 20956 11305
rect 15016 11203 15068 11212
rect 15016 11169 15025 11203
rect 15025 11169 15059 11203
rect 15059 11169 15068 11203
rect 15016 11160 15068 11169
rect 16304 11228 16356 11280
rect 20628 11228 20680 11280
rect 16212 11203 16264 11212
rect 16212 11169 16221 11203
rect 16221 11169 16255 11203
rect 16255 11169 16264 11203
rect 16212 11160 16264 11169
rect 17868 11160 17920 11212
rect 20260 11203 20312 11212
rect 20260 11169 20269 11203
rect 20269 11169 20303 11203
rect 20303 11169 20312 11203
rect 20260 11160 20312 11169
rect 12624 11092 12676 11144
rect 13728 11092 13780 11144
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 15660 11092 15712 11144
rect 16856 11092 16908 11144
rect 17132 11135 17184 11144
rect 17132 11101 17141 11135
rect 17141 11101 17175 11135
rect 17175 11101 17184 11135
rect 17132 11092 17184 11101
rect 19432 11092 19484 11144
rect 19892 11092 19944 11144
rect 7380 11024 7432 11076
rect 8208 11024 8260 11076
rect 5632 10956 5684 11008
rect 6736 10956 6788 11008
rect 9496 10956 9548 11008
rect 11060 11024 11112 11076
rect 14188 11024 14240 11076
rect 15568 11067 15620 11076
rect 15568 11033 15577 11067
rect 15577 11033 15611 11067
rect 15611 11033 15620 11067
rect 15568 11024 15620 11033
rect 16580 11024 16632 11076
rect 18144 11024 18196 11076
rect 18880 11024 18932 11076
rect 19064 11024 19116 11076
rect 10416 10956 10468 11008
rect 16488 10956 16540 11008
rect 18604 10956 18656 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 3240 10795 3292 10804
rect 3240 10761 3249 10795
rect 3249 10761 3283 10795
rect 3283 10761 3292 10795
rect 3240 10752 3292 10761
rect 7104 10752 7156 10804
rect 10232 10795 10284 10804
rect 10232 10761 10241 10795
rect 10241 10761 10275 10795
rect 10275 10761 10284 10795
rect 10232 10752 10284 10761
rect 10416 10752 10468 10804
rect 6000 10684 6052 10736
rect 3516 10659 3568 10668
rect 3516 10625 3525 10659
rect 3525 10625 3559 10659
rect 3559 10625 3568 10659
rect 3516 10616 3568 10625
rect 6644 10616 6696 10668
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 11612 10752 11664 10804
rect 14280 10752 14332 10804
rect 16212 10752 16264 10804
rect 16304 10752 16356 10804
rect 19800 10752 19852 10804
rect 1676 10548 1728 10600
rect 3148 10548 3200 10600
rect 4160 10591 4212 10600
rect 4160 10557 4169 10591
rect 4169 10557 4203 10591
rect 4203 10557 4212 10591
rect 4160 10548 4212 10557
rect 5448 10548 5500 10600
rect 7656 10548 7708 10600
rect 8484 10548 8536 10600
rect 10508 10591 10560 10600
rect 10508 10557 10517 10591
rect 10517 10557 10551 10591
rect 10551 10557 10560 10591
rect 10508 10548 10560 10557
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 2504 10480 2556 10532
rect 3976 10480 4028 10532
rect 1952 10412 2004 10464
rect 3240 10412 3292 10464
rect 5632 10412 5684 10464
rect 7472 10480 7524 10532
rect 9772 10480 9824 10532
rect 14464 10616 14516 10668
rect 15108 10616 15160 10668
rect 15568 10659 15620 10668
rect 15568 10625 15577 10659
rect 15577 10625 15611 10659
rect 15611 10625 15620 10659
rect 15568 10616 15620 10625
rect 15752 10659 15804 10668
rect 15752 10625 15761 10659
rect 15761 10625 15795 10659
rect 15795 10625 15804 10659
rect 15752 10616 15804 10625
rect 16488 10616 16540 10668
rect 12716 10591 12768 10600
rect 12716 10557 12750 10591
rect 12750 10557 12768 10591
rect 12716 10548 12768 10557
rect 12992 10548 13044 10600
rect 10232 10412 10284 10464
rect 11244 10412 11296 10464
rect 13728 10412 13780 10464
rect 16028 10412 16080 10464
rect 19800 10616 19852 10668
rect 19984 10616 20036 10668
rect 20628 10659 20680 10668
rect 20628 10625 20637 10659
rect 20637 10625 20671 10659
rect 20671 10625 20680 10659
rect 20628 10616 20680 10625
rect 18512 10591 18564 10600
rect 18512 10557 18521 10591
rect 18521 10557 18555 10591
rect 18555 10557 18564 10591
rect 18512 10548 18564 10557
rect 19524 10548 19576 10600
rect 20444 10548 20496 10600
rect 20536 10548 20588 10600
rect 16580 10455 16632 10464
rect 16580 10421 16589 10455
rect 16589 10421 16623 10455
rect 16623 10421 16632 10455
rect 16580 10412 16632 10421
rect 18328 10412 18380 10464
rect 19156 10412 19208 10464
rect 19708 10412 19760 10464
rect 19892 10455 19944 10464
rect 19892 10421 19901 10455
rect 19901 10421 19935 10455
rect 19935 10421 19944 10455
rect 19892 10412 19944 10421
rect 20168 10455 20220 10464
rect 20168 10421 20177 10455
rect 20177 10421 20211 10455
rect 20211 10421 20220 10455
rect 20168 10412 20220 10421
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 2504 10208 2556 10260
rect 4068 10208 4120 10260
rect 5632 10140 5684 10192
rect 7564 10208 7616 10260
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 8944 10208 8996 10260
rect 9680 10251 9732 10260
rect 9680 10217 9689 10251
rect 9689 10217 9723 10251
rect 9723 10217 9732 10251
rect 9680 10208 9732 10217
rect 16856 10251 16908 10260
rect 16856 10217 16865 10251
rect 16865 10217 16899 10251
rect 16899 10217 16908 10251
rect 16856 10208 16908 10217
rect 2228 10072 2280 10124
rect 4160 10072 4212 10124
rect 5080 10072 5132 10124
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 5724 10072 5776 10124
rect 7748 10072 7800 10124
rect 9496 10072 9548 10124
rect 9680 10072 9732 10124
rect 9956 10072 10008 10124
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 7932 10047 7984 10056
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 3608 9868 3660 9920
rect 4068 9868 4120 9920
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 9956 9936 10008 9988
rect 9772 9868 9824 9920
rect 10232 9868 10284 9920
rect 10692 10140 10744 10192
rect 11152 10072 11204 10124
rect 11612 10072 11664 10124
rect 11980 10115 12032 10124
rect 11980 10081 11989 10115
rect 11989 10081 12023 10115
rect 12023 10081 12032 10115
rect 11980 10072 12032 10081
rect 12716 10140 12768 10192
rect 13728 10140 13780 10192
rect 13820 10140 13872 10192
rect 16304 10140 16356 10192
rect 19892 10140 19944 10192
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 11244 10004 11296 10013
rect 12440 10072 12492 10124
rect 14004 10072 14056 10124
rect 14188 10072 14240 10124
rect 15384 10072 15436 10124
rect 15752 10115 15804 10124
rect 15752 10081 15775 10115
rect 15775 10081 15804 10115
rect 15752 10072 15804 10081
rect 16028 10072 16080 10124
rect 16764 10072 16816 10124
rect 17132 10115 17184 10124
rect 17132 10081 17141 10115
rect 17141 10081 17175 10115
rect 17175 10081 17184 10115
rect 17132 10072 17184 10081
rect 15108 10004 15160 10056
rect 15476 10047 15528 10056
rect 15476 10013 15485 10047
rect 15485 10013 15519 10047
rect 15519 10013 15528 10047
rect 15476 10004 15528 10013
rect 19156 10047 19208 10056
rect 19156 10013 19165 10047
rect 19165 10013 19199 10047
rect 19199 10013 19208 10047
rect 19156 10004 19208 10013
rect 12624 9936 12676 9988
rect 12900 9868 12952 9920
rect 13360 9868 13412 9920
rect 18604 9868 18656 9920
rect 20536 9911 20588 9920
rect 20536 9877 20545 9911
rect 20545 9877 20579 9911
rect 20579 9877 20588 9911
rect 20536 9868 20588 9877
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 1860 9639 1912 9648
rect 1860 9605 1869 9639
rect 1869 9605 1903 9639
rect 1903 9605 1912 9639
rect 1860 9596 1912 9605
rect 2872 9639 2924 9648
rect 2872 9605 2881 9639
rect 2881 9605 2915 9639
rect 2915 9605 2924 9639
rect 2872 9596 2924 9605
rect 4252 9596 4304 9648
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 3884 9528 3936 9580
rect 5632 9596 5684 9648
rect 4804 9528 4856 9580
rect 5724 9528 5776 9580
rect 3516 9460 3568 9512
rect 3792 9460 3844 9512
rect 5172 9460 5224 9512
rect 5356 9460 5408 9512
rect 7932 9664 7984 9716
rect 8668 9664 8720 9716
rect 8760 9664 8812 9716
rect 9496 9664 9548 9716
rect 6920 9639 6972 9648
rect 6920 9605 6929 9639
rect 6929 9605 6963 9639
rect 6963 9605 6972 9639
rect 6920 9596 6972 9605
rect 9956 9664 10008 9716
rect 13820 9664 13872 9716
rect 15384 9707 15436 9716
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 7472 9571 7524 9580
rect 7472 9537 7481 9571
rect 7481 9537 7515 9571
rect 7515 9537 7524 9571
rect 7472 9528 7524 9537
rect 7840 9528 7892 9580
rect 8576 9528 8628 9580
rect 8668 9528 8720 9580
rect 11060 9596 11112 9648
rect 13268 9596 13320 9648
rect 13728 9596 13780 9648
rect 13912 9596 13964 9648
rect 15384 9673 15393 9707
rect 15393 9673 15427 9707
rect 15427 9673 15436 9707
rect 15384 9664 15436 9673
rect 15660 9639 15712 9648
rect 10600 9460 10652 9512
rect 10692 9460 10744 9512
rect 13820 9528 13872 9580
rect 14004 9571 14056 9580
rect 14004 9537 14013 9571
rect 14013 9537 14047 9571
rect 14047 9537 14056 9571
rect 14004 9528 14056 9537
rect 15660 9605 15669 9639
rect 15669 9605 15703 9639
rect 15703 9605 15712 9639
rect 15660 9596 15712 9605
rect 16304 9664 16356 9716
rect 17960 9664 18012 9716
rect 4712 9392 4764 9444
rect 1400 9367 1452 9376
rect 1400 9333 1409 9367
rect 1409 9333 1443 9367
rect 1443 9333 1452 9367
rect 1400 9324 1452 9333
rect 1952 9324 2004 9376
rect 2780 9324 2832 9376
rect 4068 9324 4120 9376
rect 6184 9392 6236 9444
rect 8300 9392 8352 9444
rect 9312 9392 9364 9444
rect 9404 9392 9456 9444
rect 16488 9528 16540 9580
rect 19432 9596 19484 9648
rect 19524 9596 19576 9648
rect 17960 9460 18012 9512
rect 19340 9460 19392 9512
rect 12900 9392 12952 9444
rect 13176 9435 13228 9444
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 13176 9392 13228 9401
rect 14004 9392 14056 9444
rect 5816 9367 5868 9376
rect 5816 9333 5825 9367
rect 5825 9333 5859 9367
rect 5859 9333 5868 9367
rect 5816 9324 5868 9333
rect 5908 9324 5960 9376
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 10416 9367 10468 9376
rect 10416 9333 10425 9367
rect 10425 9333 10459 9367
rect 10459 9333 10468 9367
rect 10416 9324 10468 9333
rect 10876 9367 10928 9376
rect 10876 9333 10885 9367
rect 10885 9333 10919 9367
rect 10919 9333 10928 9367
rect 10876 9324 10928 9333
rect 13084 9324 13136 9376
rect 13268 9367 13320 9376
rect 13268 9333 13277 9367
rect 13277 9333 13311 9367
rect 13311 9333 13320 9367
rect 13268 9324 13320 9333
rect 13728 9324 13780 9376
rect 19156 9392 19208 9444
rect 20536 9460 20588 9512
rect 17040 9367 17092 9376
rect 17040 9333 17049 9367
rect 17049 9333 17083 9367
rect 17083 9333 17092 9367
rect 17040 9324 17092 9333
rect 17684 9324 17736 9376
rect 18972 9324 19024 9376
rect 20352 9324 20404 9376
rect 20444 9324 20496 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 2780 9120 2832 9172
rect 3332 9163 3384 9172
rect 3332 9129 3341 9163
rect 3341 9129 3375 9163
rect 3375 9129 3384 9163
rect 3332 9120 3384 9129
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 4068 9163 4120 9172
rect 3424 9120 3476 9129
rect 4068 9129 4077 9163
rect 4077 9129 4111 9163
rect 4111 9129 4120 9163
rect 4068 9120 4120 9129
rect 4712 9120 4764 9172
rect 8484 9120 8536 9172
rect 14004 9120 14056 9172
rect 14556 9120 14608 9172
rect 15016 9120 15068 9172
rect 15568 9120 15620 9172
rect 16212 9120 16264 9172
rect 17684 9120 17736 9172
rect 17868 9120 17920 9172
rect 18880 9120 18932 9172
rect 1400 9052 1452 9104
rect 2228 8984 2280 9036
rect 2412 8959 2464 8968
rect 2412 8925 2421 8959
rect 2421 8925 2455 8959
rect 2455 8925 2464 8959
rect 2412 8916 2464 8925
rect 2688 8916 2740 8968
rect 4252 8984 4304 9036
rect 12624 9052 12676 9104
rect 13084 9052 13136 9104
rect 3608 8916 3660 8968
rect 4804 8916 4856 8968
rect 6000 8984 6052 9036
rect 7196 8984 7248 9036
rect 7564 8984 7616 9036
rect 8208 8984 8260 9036
rect 8576 9027 8628 9036
rect 8576 8993 8585 9027
rect 8585 8993 8619 9027
rect 8619 8993 8628 9027
rect 10600 9027 10652 9036
rect 8576 8984 8628 8993
rect 10600 8993 10609 9027
rect 10609 8993 10643 9027
rect 10643 8993 10652 9027
rect 10600 8984 10652 8993
rect 12348 8984 12400 9036
rect 13544 8984 13596 9036
rect 7656 8916 7708 8968
rect 3976 8848 4028 8900
rect 7472 8848 7524 8900
rect 8300 8916 8352 8968
rect 8760 8916 8812 8968
rect 12164 8916 12216 8968
rect 12440 8959 12492 8968
rect 12440 8925 12449 8959
rect 12449 8925 12483 8959
rect 12483 8925 12492 8959
rect 12440 8916 12492 8925
rect 12256 8848 12308 8900
rect 4068 8780 4120 8832
rect 9496 8780 9548 8832
rect 11888 8823 11940 8832
rect 11888 8789 11897 8823
rect 11897 8789 11931 8823
rect 11931 8789 11940 8823
rect 11888 8780 11940 8789
rect 13728 8780 13780 8832
rect 14464 9052 14516 9104
rect 14648 8984 14700 9036
rect 16580 8984 16632 9036
rect 15384 8916 15436 8968
rect 15844 8959 15896 8968
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 16488 8916 16540 8968
rect 17040 9052 17092 9104
rect 17316 9052 17368 9104
rect 19800 9052 19852 9104
rect 20168 9120 20220 9172
rect 20352 9052 20404 9104
rect 17960 8984 18012 9036
rect 19064 9027 19116 9036
rect 19064 8993 19073 9027
rect 19073 8993 19107 9027
rect 19107 8993 19116 9027
rect 19064 8984 19116 8993
rect 17408 8959 17460 8968
rect 15200 8848 15252 8900
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 19340 8959 19392 8968
rect 19340 8925 19349 8959
rect 19349 8925 19383 8959
rect 19383 8925 19392 8959
rect 19340 8916 19392 8925
rect 20444 8959 20496 8968
rect 20444 8925 20453 8959
rect 20453 8925 20487 8959
rect 20487 8925 20496 8959
rect 20444 8916 20496 8925
rect 16948 8848 17000 8900
rect 17224 8848 17276 8900
rect 19156 8780 19208 8832
rect 20076 8780 20128 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2688 8576 2740 8628
rect 3608 8619 3660 8628
rect 3608 8585 3617 8619
rect 3617 8585 3651 8619
rect 3651 8585 3660 8619
rect 3608 8576 3660 8585
rect 3240 8508 3292 8560
rect 5816 8576 5868 8628
rect 6828 8619 6880 8628
rect 6828 8585 6837 8619
rect 6837 8585 6871 8619
rect 6871 8585 6880 8619
rect 6828 8576 6880 8585
rect 3884 8508 3936 8560
rect 7656 8576 7708 8628
rect 9404 8576 9456 8628
rect 10140 8576 10192 8628
rect 10508 8576 10560 8628
rect 11152 8576 11204 8628
rect 12624 8576 12676 8628
rect 13820 8619 13872 8628
rect 13820 8585 13829 8619
rect 13829 8585 13863 8619
rect 13863 8585 13872 8619
rect 13820 8576 13872 8585
rect 14004 8576 14056 8628
rect 15844 8576 15896 8628
rect 7012 8508 7064 8560
rect 7748 8508 7800 8560
rect 10048 8508 10100 8560
rect 10232 8508 10284 8560
rect 1676 8440 1728 8492
rect 3792 8440 3844 8492
rect 5172 8440 5224 8492
rect 5448 8440 5500 8492
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 7564 8440 7616 8492
rect 8484 8483 8536 8492
rect 8484 8449 8493 8483
rect 8493 8449 8527 8483
rect 8527 8449 8536 8483
rect 8484 8440 8536 8449
rect 8944 8440 8996 8492
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 11152 8440 11204 8492
rect 12348 8440 12400 8492
rect 15200 8508 15252 8560
rect 16856 8576 16908 8628
rect 18880 8576 18932 8628
rect 17316 8508 17368 8560
rect 2320 8372 2372 8424
rect 2504 8372 2556 8424
rect 6828 8372 6880 8424
rect 11888 8372 11940 8424
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 12440 8372 12492 8381
rect 16764 8440 16816 8492
rect 17224 8440 17276 8492
rect 17868 8440 17920 8492
rect 19248 8576 19300 8628
rect 19984 8576 20036 8628
rect 17132 8372 17184 8424
rect 17500 8372 17552 8424
rect 18880 8372 18932 8424
rect 2412 8304 2464 8356
rect 2596 8236 2648 8288
rect 3240 8236 3292 8288
rect 3792 8236 3844 8288
rect 3976 8279 4028 8288
rect 3976 8245 3985 8279
rect 3985 8245 4019 8279
rect 4019 8245 4028 8279
rect 3976 8236 4028 8245
rect 4436 8279 4488 8288
rect 4436 8245 4445 8279
rect 4445 8245 4479 8279
rect 4479 8245 4488 8279
rect 4436 8236 4488 8245
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 5172 8236 5224 8288
rect 5816 8236 5868 8288
rect 6460 8304 6512 8356
rect 6552 8304 6604 8356
rect 7380 8304 7432 8356
rect 10692 8304 10744 8356
rect 11060 8304 11112 8356
rect 12808 8304 12860 8356
rect 12900 8304 12952 8356
rect 6644 8236 6696 8288
rect 10232 8236 10284 8288
rect 10324 8279 10376 8288
rect 10324 8245 10333 8279
rect 10333 8245 10367 8279
rect 10367 8245 10376 8279
rect 10324 8236 10376 8245
rect 13452 8236 13504 8288
rect 16580 8304 16632 8356
rect 16764 8347 16816 8356
rect 16764 8313 16773 8347
rect 16773 8313 16807 8347
rect 16807 8313 16816 8347
rect 16764 8304 16816 8313
rect 15752 8279 15804 8288
rect 15752 8245 15761 8279
rect 15761 8245 15795 8279
rect 15795 8245 15804 8279
rect 15752 8236 15804 8245
rect 15844 8236 15896 8288
rect 17040 8236 17092 8288
rect 17868 8236 17920 8288
rect 19064 8304 19116 8356
rect 19432 8372 19484 8424
rect 20444 8372 20496 8424
rect 18512 8279 18564 8288
rect 18512 8245 18521 8279
rect 18521 8245 18555 8279
rect 18555 8245 18564 8279
rect 18512 8236 18564 8245
rect 20444 8236 20496 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 4988 8032 5040 8084
rect 5356 8032 5408 8084
rect 6552 8075 6604 8084
rect 6552 8041 6561 8075
rect 6561 8041 6595 8075
rect 6595 8041 6604 8075
rect 6552 8032 6604 8041
rect 9312 8075 9364 8084
rect 9312 8041 9321 8075
rect 9321 8041 9355 8075
rect 9355 8041 9364 8075
rect 9312 8032 9364 8041
rect 10048 8075 10100 8084
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 10416 8032 10468 8084
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 11060 8075 11112 8084
rect 11060 8041 11069 8075
rect 11069 8041 11103 8075
rect 11103 8041 11112 8075
rect 11060 8032 11112 8041
rect 12532 8075 12584 8084
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 12624 8075 12676 8084
rect 12624 8041 12633 8075
rect 12633 8041 12667 8075
rect 12667 8041 12676 8075
rect 12624 8032 12676 8041
rect 13268 8032 13320 8084
rect 14464 8032 14516 8084
rect 15844 8032 15896 8084
rect 15936 8032 15988 8084
rect 16396 8032 16448 8084
rect 4896 7964 4948 8016
rect 5264 7964 5316 8016
rect 8944 7964 8996 8016
rect 2044 7896 2096 7948
rect 3424 7896 3476 7948
rect 4988 7896 5040 7948
rect 9036 7896 9088 7948
rect 9496 7964 9548 8016
rect 11888 7964 11940 8016
rect 15200 7964 15252 8016
rect 15568 8007 15620 8016
rect 15568 7973 15602 8007
rect 15602 7973 15620 8007
rect 15568 7964 15620 7973
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 3792 7828 3844 7880
rect 5172 7828 5224 7880
rect 5264 7828 5316 7880
rect 4804 7760 4856 7812
rect 5448 7760 5500 7812
rect 2596 7692 2648 7744
rect 2964 7692 3016 7744
rect 3792 7692 3844 7744
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 9128 7828 9180 7880
rect 10140 7828 10192 7880
rect 10968 7896 11020 7948
rect 11612 7896 11664 7948
rect 12624 7896 12676 7948
rect 12716 7896 12768 7948
rect 13268 7896 13320 7948
rect 13452 7896 13504 7948
rect 15016 7896 15068 7948
rect 17408 8032 17460 8084
rect 19432 8032 19484 8084
rect 19616 8032 19668 8084
rect 17224 8007 17276 8016
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 13728 7871 13780 7880
rect 12808 7828 12860 7837
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 14832 7871 14884 7880
rect 6920 7692 6972 7744
rect 10600 7692 10652 7744
rect 13176 7760 13228 7812
rect 13268 7760 13320 7812
rect 14464 7760 14516 7812
rect 14004 7692 14056 7744
rect 14832 7837 14841 7871
rect 14841 7837 14875 7871
rect 14875 7837 14884 7871
rect 14832 7828 14884 7837
rect 16856 7828 16908 7880
rect 17224 7973 17258 8007
rect 17258 7973 17276 8007
rect 17224 7964 17276 7973
rect 17868 7964 17920 8016
rect 17684 7692 17736 7744
rect 17868 7692 17920 7744
rect 19156 7896 19208 7948
rect 20904 7871 20956 7880
rect 20904 7837 20913 7871
rect 20913 7837 20947 7871
rect 20947 7837 20956 7871
rect 20904 7828 20956 7837
rect 19248 7692 19300 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 3056 7488 3108 7540
rect 4252 7488 4304 7540
rect 5540 7531 5592 7540
rect 5540 7497 5549 7531
rect 5549 7497 5583 7531
rect 5583 7497 5592 7531
rect 5540 7488 5592 7497
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 7288 7488 7340 7540
rect 8944 7488 8996 7540
rect 2872 7395 2924 7404
rect 2872 7361 2881 7395
rect 2881 7361 2915 7395
rect 2915 7361 2924 7395
rect 2872 7352 2924 7361
rect 2596 7327 2648 7336
rect 2596 7293 2605 7327
rect 2605 7293 2639 7327
rect 2639 7293 2648 7327
rect 2596 7284 2648 7293
rect 2688 7284 2740 7336
rect 5172 7352 5224 7404
rect 4252 7284 4304 7336
rect 5264 7284 5316 7336
rect 6920 7420 6972 7472
rect 5448 7352 5500 7404
rect 8760 7420 8812 7472
rect 10232 7488 10284 7540
rect 11060 7488 11112 7540
rect 12072 7488 12124 7540
rect 13268 7488 13320 7540
rect 13452 7531 13504 7540
rect 13452 7497 13461 7531
rect 13461 7497 13495 7531
rect 13495 7497 13504 7531
rect 13452 7488 13504 7497
rect 13544 7488 13596 7540
rect 10324 7420 10376 7472
rect 10600 7420 10652 7472
rect 7196 7352 7248 7404
rect 9036 7395 9088 7404
rect 9036 7361 9045 7395
rect 9045 7361 9079 7395
rect 9079 7361 9088 7395
rect 9036 7352 9088 7361
rect 10140 7352 10192 7404
rect 11152 7352 11204 7404
rect 11520 7420 11572 7472
rect 5448 7216 5500 7268
rect 8116 7284 8168 7336
rect 9128 7284 9180 7336
rect 10600 7284 10652 7336
rect 10968 7284 11020 7336
rect 13360 7352 13412 7404
rect 16304 7488 16356 7540
rect 18512 7488 18564 7540
rect 18972 7488 19024 7540
rect 15016 7420 15068 7472
rect 20536 7420 20588 7472
rect 14832 7352 14884 7404
rect 15568 7352 15620 7404
rect 16028 7352 16080 7404
rect 16396 7395 16448 7404
rect 16396 7361 16405 7395
rect 16405 7361 16439 7395
rect 16439 7361 16448 7395
rect 16396 7352 16448 7361
rect 17316 7395 17368 7404
rect 17316 7361 17325 7395
rect 17325 7361 17359 7395
rect 17359 7361 17368 7395
rect 17316 7352 17368 7361
rect 17868 7352 17920 7404
rect 17960 7352 18012 7404
rect 19248 7352 19300 7404
rect 14556 7284 14608 7336
rect 12624 7216 12676 7268
rect 13452 7216 13504 7268
rect 15292 7284 15344 7336
rect 16488 7284 16540 7336
rect 3608 7191 3660 7200
rect 3608 7157 3617 7191
rect 3617 7157 3651 7191
rect 3651 7157 3660 7191
rect 3608 7148 3660 7157
rect 4712 7148 4764 7200
rect 6000 7191 6052 7200
rect 6000 7157 6009 7191
rect 6009 7157 6043 7191
rect 6043 7157 6052 7191
rect 6000 7148 6052 7157
rect 7472 7148 7524 7200
rect 9680 7148 9732 7200
rect 10416 7148 10468 7200
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 11888 7148 11940 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12808 7191 12860 7200
rect 12440 7148 12492 7157
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 12808 7148 12860 7157
rect 13176 7148 13228 7200
rect 14372 7148 14424 7200
rect 16212 7148 16264 7200
rect 19432 7284 19484 7336
rect 20628 7352 20680 7404
rect 19892 7284 19944 7336
rect 20260 7216 20312 7268
rect 17224 7191 17276 7200
rect 17224 7157 17233 7191
rect 17233 7157 17267 7191
rect 17267 7157 17276 7191
rect 17224 7148 17276 7157
rect 18512 7191 18564 7200
rect 18512 7157 18521 7191
rect 18521 7157 18555 7191
rect 18555 7157 18564 7191
rect 18512 7148 18564 7157
rect 19524 7191 19576 7200
rect 19524 7157 19533 7191
rect 19533 7157 19567 7191
rect 19567 7157 19576 7191
rect 19524 7148 19576 7157
rect 19616 7191 19668 7200
rect 19616 7157 19625 7191
rect 19625 7157 19659 7191
rect 19659 7157 19668 7191
rect 19616 7148 19668 7157
rect 19892 7148 19944 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 2044 6987 2096 6996
rect 2044 6953 2053 6987
rect 2053 6953 2087 6987
rect 2087 6953 2096 6987
rect 2044 6944 2096 6953
rect 2964 6944 3016 6996
rect 3608 6944 3660 6996
rect 4896 6944 4948 6996
rect 5908 6944 5960 6996
rect 6920 6944 6972 6996
rect 7288 6944 7340 6996
rect 9680 6987 9732 6996
rect 9680 6953 9689 6987
rect 9689 6953 9723 6987
rect 9723 6953 9732 6987
rect 9680 6944 9732 6953
rect 12808 6944 12860 6996
rect 13268 6944 13320 6996
rect 15292 6987 15344 6996
rect 3976 6876 4028 6928
rect 7104 6919 7156 6928
rect 5448 6808 5500 6860
rect 6368 6808 6420 6860
rect 7104 6885 7113 6919
rect 7113 6885 7147 6919
rect 7147 6885 7156 6919
rect 7104 6876 7156 6885
rect 7564 6876 7616 6928
rect 11612 6876 11664 6928
rect 2504 6783 2556 6792
rect 2504 6749 2513 6783
rect 2513 6749 2547 6783
rect 2547 6749 2556 6783
rect 2504 6740 2556 6749
rect 2596 6783 2648 6792
rect 2596 6749 2605 6783
rect 2605 6749 2639 6783
rect 2639 6749 2648 6783
rect 2596 6740 2648 6749
rect 5908 6783 5960 6792
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 8024 6808 8076 6860
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 11060 6808 11112 6860
rect 11980 6876 12032 6928
rect 12164 6876 12216 6928
rect 15292 6953 15301 6987
rect 15301 6953 15335 6987
rect 15335 6953 15344 6987
rect 15292 6944 15344 6953
rect 15752 6944 15804 6996
rect 16396 6944 16448 6996
rect 16764 6919 16816 6928
rect 16764 6885 16773 6919
rect 16773 6885 16807 6919
rect 16807 6885 16816 6919
rect 17408 6944 17460 6996
rect 17684 6944 17736 6996
rect 17868 6944 17920 6996
rect 18512 6944 18564 6996
rect 16764 6876 16816 6885
rect 18604 6876 18656 6928
rect 13360 6808 13412 6860
rect 14464 6808 14516 6860
rect 18512 6808 18564 6860
rect 18788 6808 18840 6860
rect 7012 6740 7064 6792
rect 8300 6740 8352 6792
rect 9220 6740 9272 6792
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 4068 6604 4120 6656
rect 5448 6604 5500 6656
rect 5540 6604 5592 6656
rect 6460 6647 6512 6656
rect 6460 6613 6469 6647
rect 6469 6613 6503 6647
rect 6503 6613 6512 6647
rect 6460 6604 6512 6613
rect 8116 6672 8168 6724
rect 8760 6672 8812 6724
rect 11428 6672 11480 6724
rect 7564 6604 7616 6656
rect 7748 6647 7800 6656
rect 7748 6613 7757 6647
rect 7757 6613 7791 6647
rect 7791 6613 7800 6647
rect 7748 6604 7800 6613
rect 7840 6604 7892 6656
rect 11060 6604 11112 6656
rect 13912 6740 13964 6792
rect 14832 6740 14884 6792
rect 15660 6740 15712 6792
rect 16028 6740 16080 6792
rect 16856 6783 16908 6792
rect 16856 6749 16865 6783
rect 16865 6749 16899 6783
rect 16899 6749 16908 6783
rect 16856 6740 16908 6749
rect 16948 6740 17000 6792
rect 19432 6944 19484 6996
rect 19524 6944 19576 6996
rect 20904 6876 20956 6928
rect 19892 6808 19944 6860
rect 20168 6851 20220 6860
rect 20168 6817 20177 6851
rect 20177 6817 20211 6851
rect 20211 6817 20220 6851
rect 20168 6808 20220 6817
rect 12532 6672 12584 6724
rect 16764 6672 16816 6724
rect 19156 6740 19208 6792
rect 20260 6783 20312 6792
rect 18788 6672 18840 6724
rect 20260 6749 20269 6783
rect 20269 6749 20303 6783
rect 20303 6749 20312 6783
rect 20260 6740 20312 6749
rect 12256 6604 12308 6656
rect 12808 6604 12860 6656
rect 14648 6604 14700 6656
rect 17224 6604 17276 6656
rect 19708 6604 19760 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 2688 6400 2740 6452
rect 3424 6443 3476 6452
rect 3424 6409 3433 6443
rect 3433 6409 3467 6443
rect 3467 6409 3476 6443
rect 3424 6400 3476 6409
rect 2596 6196 2648 6248
rect 5540 6400 5592 6452
rect 5908 6400 5960 6452
rect 1952 6128 2004 6180
rect 3332 6128 3384 6180
rect 3700 6128 3752 6180
rect 4804 6239 4856 6248
rect 4804 6205 4813 6239
rect 4813 6205 4847 6239
rect 4847 6205 4856 6239
rect 4804 6196 4856 6205
rect 7196 6332 7248 6384
rect 8024 6332 8076 6384
rect 8208 6332 8260 6384
rect 10048 6400 10100 6452
rect 10140 6400 10192 6452
rect 11612 6400 11664 6452
rect 13452 6400 13504 6452
rect 13912 6443 13964 6452
rect 13912 6409 13921 6443
rect 13921 6409 13955 6443
rect 13955 6409 13964 6443
rect 13912 6400 13964 6409
rect 14832 6400 14884 6452
rect 15660 6400 15712 6452
rect 16488 6400 16540 6452
rect 16672 6400 16724 6452
rect 17500 6400 17552 6452
rect 18604 6400 18656 6452
rect 19616 6400 19668 6452
rect 20260 6443 20312 6452
rect 20260 6409 20269 6443
rect 20269 6409 20303 6443
rect 20303 6409 20312 6443
rect 20260 6400 20312 6409
rect 7748 6264 7800 6316
rect 10876 6332 10928 6384
rect 12348 6332 12400 6384
rect 9220 6264 9272 6316
rect 6828 6196 6880 6248
rect 8116 6196 8168 6248
rect 8484 6196 8536 6248
rect 10508 6264 10560 6316
rect 10600 6307 10652 6316
rect 10600 6273 10609 6307
rect 10609 6273 10643 6307
rect 10643 6273 10652 6307
rect 10600 6264 10652 6273
rect 10968 6264 11020 6316
rect 14556 6332 14608 6384
rect 9680 6196 9732 6248
rect 12164 6196 12216 6248
rect 5540 6128 5592 6180
rect 2780 6060 2832 6112
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 3792 6060 3844 6069
rect 4804 6060 4856 6112
rect 10140 6128 10192 6180
rect 6276 6060 6328 6112
rect 7748 6060 7800 6112
rect 8576 6060 8628 6112
rect 8944 6060 8996 6112
rect 9864 6060 9916 6112
rect 11612 6128 11664 6180
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 14832 6264 14884 6316
rect 15844 6264 15896 6316
rect 18420 6264 18472 6316
rect 18788 6307 18840 6316
rect 18788 6273 18797 6307
rect 18797 6273 18831 6307
rect 18831 6273 18840 6307
rect 18788 6264 18840 6273
rect 19156 6332 19208 6384
rect 19524 6264 19576 6316
rect 19708 6307 19760 6316
rect 19708 6273 19717 6307
rect 19717 6273 19751 6307
rect 19751 6273 19760 6307
rect 19708 6264 19760 6273
rect 20628 6264 20680 6316
rect 12808 6239 12860 6248
rect 12808 6205 12842 6239
rect 12842 6205 12860 6239
rect 12808 6196 12860 6205
rect 15476 6196 15528 6248
rect 16304 6196 16356 6248
rect 19892 6196 19944 6248
rect 14372 6128 14424 6180
rect 10416 6060 10468 6112
rect 11704 6060 11756 6112
rect 13084 6060 13136 6112
rect 14464 6060 14516 6112
rect 16672 6128 16724 6180
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 17316 6103 17368 6112
rect 17316 6069 17325 6103
rect 17325 6069 17359 6103
rect 17359 6069 17368 6103
rect 17316 6060 17368 6069
rect 20536 6128 20588 6180
rect 18788 6060 18840 6112
rect 20352 6060 20404 6112
rect 20904 6060 20956 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 2872 5856 2924 5908
rect 3792 5856 3844 5908
rect 4712 5856 4764 5908
rect 5448 5899 5500 5908
rect 5448 5865 5457 5899
rect 5457 5865 5491 5899
rect 5491 5865 5500 5899
rect 5448 5856 5500 5865
rect 7748 5856 7800 5908
rect 2688 5788 2740 5840
rect 6276 5788 6328 5840
rect 6368 5788 6420 5840
rect 4804 5720 4856 5772
rect 8300 5788 8352 5840
rect 1952 5652 2004 5704
rect 5540 5695 5592 5704
rect 5540 5661 5549 5695
rect 5549 5661 5583 5695
rect 5583 5661 5592 5695
rect 5540 5652 5592 5661
rect 8300 5652 8352 5704
rect 10784 5788 10836 5840
rect 10968 5856 11020 5908
rect 12440 5899 12492 5908
rect 12440 5865 12449 5899
rect 12449 5865 12483 5899
rect 12483 5865 12492 5899
rect 12440 5856 12492 5865
rect 15568 5856 15620 5908
rect 18420 5856 18472 5908
rect 20168 5856 20220 5908
rect 12992 5788 13044 5840
rect 13912 5788 13964 5840
rect 14648 5788 14700 5840
rect 12348 5720 12400 5772
rect 13544 5763 13596 5772
rect 13544 5729 13553 5763
rect 13553 5729 13587 5763
rect 13587 5729 13596 5763
rect 13544 5720 13596 5729
rect 15476 5763 15528 5772
rect 15476 5729 15485 5763
rect 15485 5729 15519 5763
rect 15519 5729 15528 5763
rect 15476 5720 15528 5729
rect 16304 5763 16356 5772
rect 16304 5729 16338 5763
rect 16338 5729 16356 5763
rect 16304 5720 16356 5729
rect 17224 5788 17276 5840
rect 18880 5788 18932 5840
rect 17132 5720 17184 5772
rect 20168 5763 20220 5772
rect 20168 5729 20177 5763
rect 20177 5729 20211 5763
rect 20211 5729 20220 5763
rect 20168 5720 20220 5729
rect 8944 5695 8996 5704
rect 8944 5661 8953 5695
rect 8953 5661 8987 5695
rect 8987 5661 8996 5695
rect 8944 5652 8996 5661
rect 12532 5695 12584 5704
rect 4068 5516 4120 5568
rect 7012 5516 7064 5568
rect 9036 5584 9088 5636
rect 12532 5661 12541 5695
rect 12541 5661 12575 5695
rect 12575 5661 12584 5695
rect 12532 5652 12584 5661
rect 12808 5652 12860 5704
rect 17408 5652 17460 5704
rect 18788 5652 18840 5704
rect 19800 5652 19852 5704
rect 20628 5652 20680 5704
rect 8208 5516 8260 5568
rect 10876 5516 10928 5568
rect 13176 5516 13228 5568
rect 14556 5516 14608 5568
rect 17500 5516 17552 5568
rect 20812 5584 20864 5636
rect 22468 5516 22520 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 1952 5312 2004 5364
rect 3240 5244 3292 5296
rect 1400 5108 1452 5160
rect 1952 5151 2004 5160
rect 1952 5117 1961 5151
rect 1961 5117 1995 5151
rect 1995 5117 2004 5151
rect 1952 5108 2004 5117
rect 3976 5312 4028 5364
rect 8944 5355 8996 5364
rect 8944 5321 8953 5355
rect 8953 5321 8987 5355
rect 8987 5321 8996 5355
rect 8944 5312 8996 5321
rect 9036 5312 9088 5364
rect 12532 5312 12584 5364
rect 13452 5312 13504 5364
rect 15844 5312 15896 5364
rect 16028 5355 16080 5364
rect 16028 5321 16037 5355
rect 16037 5321 16071 5355
rect 16071 5321 16080 5355
rect 16028 5312 16080 5321
rect 17316 5312 17368 5364
rect 18696 5312 18748 5364
rect 20628 5312 20680 5364
rect 12900 5244 12952 5296
rect 6184 5176 6236 5228
rect 7104 5176 7156 5228
rect 2780 5040 2832 5092
rect 3792 5108 3844 5160
rect 6736 5108 6788 5160
rect 7564 5151 7616 5160
rect 7564 5117 7573 5151
rect 7573 5117 7607 5151
rect 7607 5117 7616 5151
rect 7564 5108 7616 5117
rect 4068 5040 4120 5092
rect 4712 4972 4764 5024
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 5632 4972 5684 5024
rect 6460 5040 6512 5092
rect 10324 5108 10376 5160
rect 11336 5176 11388 5228
rect 11888 5176 11940 5228
rect 14096 5244 14148 5296
rect 18052 5244 18104 5296
rect 19616 5244 19668 5296
rect 13360 5176 13412 5228
rect 12808 5108 12860 5160
rect 14648 5219 14700 5228
rect 14648 5185 14657 5219
rect 14657 5185 14691 5219
rect 14691 5185 14700 5219
rect 14648 5176 14700 5185
rect 16948 5176 17000 5228
rect 17500 5219 17552 5228
rect 17500 5185 17509 5219
rect 17509 5185 17543 5219
rect 17543 5185 17552 5219
rect 17500 5176 17552 5185
rect 16304 5108 16356 5160
rect 18972 5176 19024 5228
rect 18880 5108 18932 5160
rect 8208 5040 8260 5092
rect 10600 5083 10652 5092
rect 10600 5049 10609 5083
rect 10609 5049 10643 5083
rect 10643 5049 10652 5083
rect 10600 5040 10652 5049
rect 11244 5040 11296 5092
rect 15200 5040 15252 5092
rect 18788 5040 18840 5092
rect 19524 5108 19576 5160
rect 20168 5040 20220 5092
rect 10784 4972 10836 5024
rect 11428 4972 11480 5024
rect 12808 5015 12860 5024
rect 12808 4981 12817 5015
rect 12817 4981 12851 5015
rect 12851 4981 12860 5015
rect 12808 4972 12860 4981
rect 13636 5015 13688 5024
rect 13636 4981 13645 5015
rect 13645 4981 13679 5015
rect 13679 4981 13688 5015
rect 13636 4972 13688 4981
rect 13728 4972 13780 5024
rect 16764 4972 16816 5024
rect 17500 4972 17552 5024
rect 18696 4972 18748 5024
rect 19984 4972 20036 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 2780 4811 2832 4820
rect 2780 4777 2789 4811
rect 2789 4777 2823 4811
rect 2823 4777 2832 4811
rect 2780 4768 2832 4777
rect 3884 4768 3936 4820
rect 6092 4768 6144 4820
rect 7012 4811 7064 4820
rect 7012 4777 7021 4811
rect 7021 4777 7055 4811
rect 7055 4777 7064 4811
rect 7012 4768 7064 4777
rect 7472 4768 7524 4820
rect 7748 4768 7800 4820
rect 8300 4768 8352 4820
rect 11428 4768 11480 4820
rect 13636 4768 13688 4820
rect 16488 4768 16540 4820
rect 17132 4768 17184 4820
rect 6184 4700 6236 4752
rect 6828 4700 6880 4752
rect 8576 4743 8628 4752
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 3148 4632 3200 4684
rect 4620 4632 4672 4684
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 8576 4709 8585 4743
rect 8585 4709 8619 4743
rect 8619 4709 8628 4743
rect 8576 4700 8628 4709
rect 11244 4700 11296 4752
rect 11336 4700 11388 4752
rect 11888 4700 11940 4752
rect 12992 4700 13044 4752
rect 14556 4700 14608 4752
rect 17776 4700 17828 4752
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 11520 4632 11572 4684
rect 13452 4632 13504 4684
rect 13544 4675 13596 4684
rect 13544 4641 13553 4675
rect 13553 4641 13587 4675
rect 13587 4641 13596 4675
rect 13544 4632 13596 4641
rect 15108 4632 15160 4684
rect 17132 4675 17184 4684
rect 17132 4641 17141 4675
rect 17141 4641 17175 4675
rect 17175 4641 17184 4675
rect 17132 4632 17184 4641
rect 17408 4675 17460 4684
rect 17408 4641 17442 4675
rect 17442 4641 17460 4675
rect 17408 4632 17460 4641
rect 20168 4811 20220 4820
rect 20168 4777 20177 4811
rect 20177 4777 20211 4811
rect 20211 4777 20220 4811
rect 20168 4768 20220 4777
rect 19064 4743 19116 4752
rect 19064 4709 19076 4743
rect 19076 4709 19116 4743
rect 19064 4700 19116 4709
rect 19524 4632 19576 4684
rect 7104 4607 7156 4616
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 7104 4564 7156 4573
rect 8208 4564 8260 4616
rect 9956 4564 10008 4616
rect 16764 4607 16816 4616
rect 5632 4496 5684 4548
rect 5264 4428 5316 4480
rect 7196 4428 7248 4480
rect 9220 4496 9272 4548
rect 10600 4428 10652 4480
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 16764 4573 16773 4607
rect 16773 4573 16807 4607
rect 16807 4573 16816 4607
rect 16764 4564 16816 4573
rect 16672 4496 16724 4548
rect 12348 4428 12400 4480
rect 12992 4428 13044 4480
rect 14924 4471 14976 4480
rect 14924 4437 14933 4471
rect 14933 4437 14967 4471
rect 14967 4437 14976 4471
rect 14924 4428 14976 4437
rect 15844 4428 15896 4480
rect 18788 4428 18840 4480
rect 21088 4428 21140 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 2780 4156 2832 4208
rect 4712 4224 4764 4276
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 5356 4020 5408 4072
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 3148 3952 3200 4004
rect 1768 3884 1820 3936
rect 2320 3927 2372 3936
rect 2320 3893 2329 3927
rect 2329 3893 2363 3927
rect 2363 3893 2372 3927
rect 2320 3884 2372 3893
rect 4068 3884 4120 3936
rect 4528 3884 4580 3936
rect 5724 3952 5776 4004
rect 6644 3952 6696 4004
rect 7380 4224 7432 4276
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 10232 4224 10284 4276
rect 11060 4224 11112 4276
rect 19984 4267 20036 4276
rect 13728 4156 13780 4208
rect 14924 4156 14976 4208
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 7564 4088 7616 4140
rect 12992 4131 13044 4140
rect 7196 4063 7248 4072
rect 7196 4029 7205 4063
rect 7205 4029 7239 4063
rect 7239 4029 7248 4063
rect 7196 4020 7248 4029
rect 7288 4020 7340 4072
rect 8392 4020 8444 4072
rect 9036 4020 9088 4072
rect 9588 4020 9640 4072
rect 10324 4063 10376 4072
rect 10324 4029 10358 4063
rect 10358 4029 10376 4063
rect 10324 4020 10376 4029
rect 7564 3952 7616 4004
rect 8208 3952 8260 4004
rect 8852 3952 8904 4004
rect 10692 3952 10744 4004
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 19984 4233 19993 4267
rect 19993 4233 20027 4267
rect 20027 4233 20036 4267
rect 19984 4224 20036 4233
rect 18788 4156 18840 4208
rect 19064 4156 19116 4208
rect 6276 3884 6328 3936
rect 11428 3927 11480 3936
rect 11428 3893 11437 3927
rect 11437 3893 11471 3927
rect 11471 3893 11480 3927
rect 11428 3884 11480 3893
rect 12624 3952 12676 4004
rect 13084 4020 13136 4072
rect 13544 4020 13596 4072
rect 14924 4020 14976 4072
rect 16856 4020 16908 4072
rect 17408 4088 17460 4140
rect 18604 4088 18656 4140
rect 18328 4020 18380 4072
rect 19340 4020 19392 4072
rect 20444 4020 20496 4072
rect 21548 4020 21600 4072
rect 13728 3952 13780 4004
rect 12164 3884 12216 3936
rect 13084 3884 13136 3936
rect 16120 3952 16172 4004
rect 17224 3952 17276 4004
rect 17960 3952 18012 4004
rect 20536 3952 20588 4004
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 15752 3884 15804 3936
rect 17040 3884 17092 3936
rect 18236 3884 18288 3936
rect 18788 3884 18840 3936
rect 18972 3927 19024 3936
rect 18972 3893 18981 3927
rect 18981 3893 19015 3927
rect 19015 3893 19024 3927
rect 18972 3884 19024 3893
rect 19340 3927 19392 3936
rect 19340 3893 19349 3927
rect 19349 3893 19383 3927
rect 19383 3893 19392 3927
rect 19340 3884 19392 3893
rect 19432 3927 19484 3936
rect 19432 3893 19441 3927
rect 19441 3893 19475 3927
rect 19475 3893 19484 3927
rect 20352 3927 20404 3936
rect 19432 3884 19484 3893
rect 20352 3893 20361 3927
rect 20361 3893 20395 3927
rect 20395 3893 20404 3927
rect 20352 3884 20404 3893
rect 20444 3927 20496 3936
rect 20444 3893 20453 3927
rect 20453 3893 20487 3927
rect 20487 3893 20496 3927
rect 20444 3884 20496 3893
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 2320 3680 2372 3732
rect 4068 3723 4120 3732
rect 4068 3689 4077 3723
rect 4077 3689 4111 3723
rect 4111 3689 4120 3723
rect 4068 3680 4120 3689
rect 4528 3723 4580 3732
rect 4528 3689 4537 3723
rect 4537 3689 4571 3723
rect 4571 3689 4580 3723
rect 4528 3680 4580 3689
rect 6920 3680 6972 3732
rect 8944 3680 8996 3732
rect 9864 3680 9916 3732
rect 13084 3723 13136 3732
rect 13084 3689 13093 3723
rect 13093 3689 13127 3723
rect 13127 3689 13136 3723
rect 13084 3680 13136 3689
rect 7196 3612 7248 3664
rect 10048 3612 10100 3664
rect 11428 3612 11480 3664
rect 11888 3612 11940 3664
rect 4160 3544 4212 3596
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 7472 3544 7524 3596
rect 8576 3544 8628 3596
rect 9864 3544 9916 3596
rect 9956 3544 10008 3596
rect 12808 3612 12860 3664
rect 14280 3680 14332 3732
rect 15752 3723 15804 3732
rect 15752 3689 15761 3723
rect 15761 3689 15795 3723
rect 15795 3689 15804 3723
rect 15752 3680 15804 3689
rect 12256 3544 12308 3596
rect 12624 3544 12676 3596
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 3148 3519 3200 3528
rect 3148 3485 3157 3519
rect 3157 3485 3191 3519
rect 3191 3485 3200 3519
rect 3148 3476 3200 3485
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 6828 3519 6880 3528
rect 204 3408 256 3460
rect 3792 3408 3844 3460
rect 5264 3408 5316 3460
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 8116 3476 8168 3528
rect 9588 3476 9640 3528
rect 11612 3476 11664 3528
rect 3976 3340 4028 3392
rect 5724 3340 5776 3392
rect 5908 3340 5960 3392
rect 7748 3340 7800 3392
rect 8208 3383 8260 3392
rect 8208 3349 8217 3383
rect 8217 3349 8251 3383
rect 8251 3349 8260 3383
rect 8208 3340 8260 3349
rect 8484 3383 8536 3392
rect 8484 3349 8493 3383
rect 8493 3349 8527 3383
rect 8527 3349 8536 3383
rect 8484 3340 8536 3349
rect 12624 3408 12676 3460
rect 18420 3680 18472 3732
rect 18696 3680 18748 3732
rect 18972 3723 19024 3732
rect 18972 3689 18981 3723
rect 18981 3689 19015 3723
rect 19015 3689 19024 3723
rect 18972 3680 19024 3689
rect 19340 3680 19392 3732
rect 17592 3612 17644 3664
rect 19432 3612 19484 3664
rect 19892 3612 19944 3664
rect 16488 3587 16540 3596
rect 16488 3553 16497 3587
rect 16497 3553 16531 3587
rect 16531 3553 16540 3587
rect 16488 3544 16540 3553
rect 12992 3476 13044 3528
rect 15016 3476 15068 3528
rect 15200 3476 15252 3528
rect 16304 3476 16356 3528
rect 18972 3544 19024 3596
rect 20260 3544 20312 3596
rect 18328 3476 18380 3528
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 16120 3408 16172 3460
rect 17776 3408 17828 3460
rect 11060 3340 11112 3392
rect 11152 3340 11204 3392
rect 12716 3383 12768 3392
rect 12716 3349 12725 3383
rect 12725 3349 12759 3383
rect 12759 3349 12768 3383
rect 12716 3340 12768 3349
rect 15476 3340 15528 3392
rect 18604 3340 18656 3392
rect 18972 3340 19024 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 3056 3136 3108 3188
rect 3884 3136 3936 3188
rect 5632 3136 5684 3188
rect 6276 3136 6328 3188
rect 1584 3068 1636 3120
rect 3240 3000 3292 3052
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 5264 3000 5316 3052
rect 5632 3000 5684 3052
rect 6184 3043 6236 3052
rect 6184 3009 6193 3043
rect 6193 3009 6227 3043
rect 6227 3009 6236 3043
rect 6184 3000 6236 3009
rect 8116 3136 8168 3188
rect 8576 3179 8628 3188
rect 8576 3145 8585 3179
rect 8585 3145 8619 3179
rect 8619 3145 8628 3179
rect 8576 3136 8628 3145
rect 9128 3136 9180 3188
rect 9312 3136 9364 3188
rect 20352 3136 20404 3188
rect 9680 3068 9732 3120
rect 13452 3068 13504 3120
rect 15384 3068 15436 3120
rect 18696 3068 18748 3120
rect 3516 2975 3568 2984
rect 3516 2941 3525 2975
rect 3525 2941 3559 2975
rect 3559 2941 3568 2975
rect 3516 2932 3568 2941
rect 4068 2932 4120 2984
rect 5816 2932 5868 2984
rect 6092 2975 6144 2984
rect 6092 2941 6101 2975
rect 6101 2941 6135 2975
rect 6135 2941 6144 2975
rect 6092 2932 6144 2941
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 7104 2975 7156 2984
rect 7104 2941 7138 2975
rect 7138 2941 7156 2975
rect 9588 3000 9640 3052
rect 11888 3000 11940 3052
rect 13084 3000 13136 3052
rect 18604 3000 18656 3052
rect 19340 3000 19392 3052
rect 7104 2932 7156 2941
rect 1124 2864 1176 2916
rect 3516 2796 3568 2848
rect 3884 2796 3936 2848
rect 4160 2839 4212 2848
rect 4160 2805 4169 2839
rect 4169 2805 4203 2839
rect 4203 2805 4212 2839
rect 4160 2796 4212 2805
rect 4344 2796 4396 2848
rect 5356 2796 5408 2848
rect 6000 2796 6052 2848
rect 8392 2864 8444 2916
rect 11152 2932 11204 2984
rect 12256 2932 12308 2984
rect 8944 2839 8996 2848
rect 8944 2805 8953 2839
rect 8953 2805 8987 2839
rect 8987 2805 8996 2839
rect 10784 2864 10836 2916
rect 12808 2975 12860 2984
rect 12808 2941 12817 2975
rect 12817 2941 12851 2975
rect 12851 2941 12860 2975
rect 12808 2932 12860 2941
rect 13176 2932 13228 2984
rect 13728 2975 13780 2984
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13728 2932 13780 2941
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 14464 2932 14516 2984
rect 15568 2975 15620 2984
rect 15568 2941 15577 2975
rect 15577 2941 15611 2975
rect 15611 2941 15620 2975
rect 15568 2932 15620 2941
rect 16672 2932 16724 2984
rect 17316 2932 17368 2984
rect 16304 2864 16356 2916
rect 8944 2796 8996 2805
rect 9956 2796 10008 2848
rect 10416 2796 10468 2848
rect 12808 2796 12860 2848
rect 13912 2796 13964 2848
rect 15016 2796 15068 2848
rect 17408 2796 17460 2848
rect 20444 2932 20496 2984
rect 20720 2975 20772 2984
rect 20720 2941 20729 2975
rect 20729 2941 20763 2975
rect 20763 2941 20772 2975
rect 20720 2932 20772 2941
rect 19156 2839 19208 2848
rect 19156 2805 19165 2839
rect 19165 2805 19199 2839
rect 19199 2805 19208 2839
rect 20260 2864 20312 2916
rect 19156 2796 19208 2805
rect 20168 2839 20220 2848
rect 20168 2805 20177 2839
rect 20177 2805 20211 2839
rect 20211 2805 20220 2839
rect 20168 2796 20220 2805
rect 20628 2796 20680 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 4344 2592 4396 2644
rect 7564 2592 7616 2644
rect 9864 2592 9916 2644
rect 10324 2592 10376 2644
rect 11612 2592 11664 2644
rect 12716 2592 12768 2644
rect 19156 2592 19208 2644
rect 8208 2524 8260 2576
rect 10600 2524 10652 2576
rect 12164 2524 12216 2576
rect 12256 2524 12308 2576
rect 8484 2320 8536 2372
rect 12440 2456 12492 2508
rect 12716 2456 12768 2508
rect 14004 2456 14056 2508
rect 17316 2524 17368 2576
rect 18880 2524 18932 2576
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 16212 2499 16264 2508
rect 16212 2465 16221 2499
rect 16221 2465 16255 2499
rect 16255 2465 16264 2499
rect 16212 2456 16264 2465
rect 16304 2456 16356 2508
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 10876 2388 10928 2440
rect 11704 2388 11756 2440
rect 15568 2388 15620 2440
rect 18512 2456 18564 2508
rect 19432 2499 19484 2508
rect 19432 2465 19441 2499
rect 19441 2465 19475 2499
rect 19475 2465 19484 2499
rect 19432 2456 19484 2465
rect 20076 2456 20128 2508
rect 17868 2388 17920 2440
rect 19248 2388 19300 2440
rect 14188 2320 14240 2372
rect 19340 2320 19392 2372
rect 10968 2295 11020 2304
rect 10968 2261 10977 2295
rect 10977 2261 11011 2295
rect 11011 2261 11020 2295
rect 10968 2252 11020 2261
rect 14464 2252 14516 2304
rect 16764 2252 16816 2304
rect 17776 2252 17828 2304
rect 18512 2295 18564 2304
rect 18512 2261 18521 2295
rect 18521 2261 18555 2295
rect 18555 2261 18564 2295
rect 18512 2252 18564 2261
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 2504 2048 2556 2100
rect 8944 2048 8996 2100
rect 10968 2048 11020 2100
rect 22008 2048 22060 2100
rect 8208 1980 8260 2032
rect 8668 1980 8720 2032
rect 11704 1980 11756 2032
rect 11980 1980 12032 2032
rect 2044 1368 2096 1420
rect 7196 1368 7248 1420
<< metal2 >>
rect 3146 22536 3202 22545
rect 3146 22471 3202 22480
rect 3054 21584 3110 21593
rect 3054 21519 3110 21528
rect 2502 21176 2558 21185
rect 2502 21111 2558 21120
rect 1950 19816 2006 19825
rect 1950 19751 2006 19760
rect 1964 19514 1992 19751
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1950 19272 2006 19281
rect 1950 19207 2006 19216
rect 1964 18970 1992 19207
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1950 18864 2006 18873
rect 1950 18799 2006 18808
rect 1964 18426 1992 18799
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1674 18320 1730 18329
rect 1674 18255 1730 18264
rect 1688 17610 1716 18255
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1780 17814 1808 18158
rect 1950 17912 2006 17921
rect 1950 17847 2006 17856
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 1676 17604 1728 17610
rect 1676 17546 1728 17552
rect 1858 17368 1914 17377
rect 1964 17338 1992 17847
rect 1858 17303 1914 17312
rect 1952 17332 2004 17338
rect 1872 16794 1900 17303
rect 1952 17274 2004 17280
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 1950 16552 2006 16561
rect 1950 16487 2006 16496
rect 1964 16250 1992 16487
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 1950 16008 2006 16017
rect 1950 15943 2006 15952
rect 1964 15706 1992 15943
rect 2516 15706 2544 21111
rect 2778 20224 2834 20233
rect 2778 20159 2834 20168
rect 2792 19174 2820 20159
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2778 15600 2834 15609
rect 1860 15564 1912 15570
rect 2778 15535 2834 15544
rect 1860 15506 1912 15512
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1780 14550 1808 14894
rect 1768 14544 1820 14550
rect 1768 14486 1820 14492
rect 1582 14104 1638 14113
rect 1582 14039 1638 14048
rect 1872 14056 1900 15506
rect 2792 15162 2820 15535
rect 3068 15162 3096 21519
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 1952 15088 2004 15094
rect 1950 15056 1952 15065
rect 2004 15056 2006 15065
rect 1950 14991 2006 15000
rect 2778 14648 2834 14657
rect 2778 14583 2834 14592
rect 2688 14340 2740 14346
rect 2688 14282 2740 14288
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 1596 13530 1624 14039
rect 1872 14028 1992 14056
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1674 13696 1730 13705
rect 1674 13631 1730 13640
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1582 13288 1638 13297
rect 1582 13223 1638 13232
rect 1596 11898 1624 13223
rect 1688 12442 1716 13631
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 11286 1440 11630
rect 1400 11280 1452 11286
rect 1400 11222 1452 11228
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1688 10062 1716 10542
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1412 9110 1440 9318
rect 1400 9104 1452 9110
rect 1400 9046 1452 9052
rect 1688 8498 1716 9998
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1412 4690 1440 5102
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 662 4040 718 4049
rect 662 3975 718 3984
rect 204 3460 256 3466
rect 204 3402 256 3408
rect 216 480 244 3402
rect 676 480 704 3975
rect 1780 3942 1808 13806
rect 1872 12306 1900 13874
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1872 9654 1900 11154
rect 1964 10470 1992 14028
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2056 12986 2084 13330
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 2148 12782 2176 13126
rect 2240 12850 2268 14214
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2596 13320 2648 13326
rect 2700 13308 2728 14282
rect 2792 14074 2820 14583
rect 3160 14550 3188 22471
rect 3790 22320 3846 22800
rect 11334 22320 11390 22800
rect 17222 22536 17278 22545
rect 17222 22471 17278 22480
rect 3606 22128 3662 22137
rect 3606 22063 3662 22072
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3056 14544 3108 14550
rect 3056 14486 3108 14492
rect 3148 14544 3200 14550
rect 3148 14486 3200 14492
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2884 13530 2912 14418
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2648 13280 2728 13308
rect 2596 13262 2648 13268
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 2228 10124 2280 10130
rect 2228 10066 2280 10072
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1964 9178 1992 9318
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2240 9042 2268 10066
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2332 8430 2360 13262
rect 2608 12646 2636 13262
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2884 12594 2912 12718
rect 2884 12566 3004 12594
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2516 11082 2544 12310
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2792 11762 2820 12106
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 2516 10266 2544 10474
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2516 9586 2544 10202
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2424 8362 2452 8910
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 2056 7002 2084 7890
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 2516 6798 2544 8366
rect 2608 8294 2636 11698
rect 2976 11694 3004 12566
rect 3068 12442 3096 14486
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2884 11336 2912 11562
rect 3068 11354 3096 12242
rect 3252 12238 3280 15982
rect 3436 15042 3464 19246
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3528 15638 3556 15982
rect 3516 15632 3568 15638
rect 3516 15574 3568 15580
rect 3620 15162 3648 22063
rect 3698 16960 3754 16969
rect 3698 16895 3754 16904
rect 3712 16250 3740 16895
rect 3700 16244 3752 16250
rect 3700 16186 3752 16192
rect 3804 15586 3832 22320
rect 4066 20632 4122 20641
rect 4066 20567 4122 20576
rect 3804 15558 3924 15586
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 3436 15014 3832 15042
rect 3516 13456 3568 13462
rect 3516 13398 3568 13404
rect 3332 13252 3384 13258
rect 3332 13194 3384 13200
rect 3344 12374 3372 13194
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3332 11824 3384 11830
rect 3332 11766 3384 11772
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3056 11348 3108 11354
rect 2884 11308 3004 11336
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2792 9466 2820 11018
rect 2884 9654 2912 11154
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2792 9438 2912 9466
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 9178 2820 9318
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2700 8634 2728 8910
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2608 7342 2636 7686
rect 2700 7342 2728 7822
rect 2884 7562 2912 9438
rect 2976 7750 3004 11308
rect 3056 11290 3108 11296
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2884 7534 3004 7562
rect 3068 7546 3096 11154
rect 3160 10606 3188 11630
rect 3240 11620 3292 11626
rect 3240 11562 3292 11568
rect 3252 11150 3280 11562
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3252 10810 3280 11086
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3252 8566 3280 10406
rect 3344 9178 3372 11766
rect 3436 9178 3464 12038
rect 3528 10674 3556 13398
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3620 9926 3648 12038
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 1952 6180 2004 6186
rect 1952 6122 2004 6128
rect 1964 5710 1992 6122
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1964 5370 1992 5646
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1964 5166 1992 5306
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2332 3738 2360 3878
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2516 3505 2544 6734
rect 2608 6254 2636 6734
rect 2700 6458 2728 7278
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2700 5846 2728 6394
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2792 5794 2820 6054
rect 2884 5914 2912 7346
rect 2976 7154 3004 7534
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2976 7126 3188 7154
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2792 5766 2912 5794
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2792 4826 2820 5034
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2792 4214 2820 4762
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2502 3496 2558 3505
rect 2502 3431 2558 3440
rect 1584 3120 1636 3126
rect 1584 3062 1636 3068
rect 1124 2916 1176 2922
rect 1124 2858 1176 2864
rect 1136 480 1164 2858
rect 1596 480 1624 3062
rect 2884 2553 2912 5766
rect 2870 2544 2926 2553
rect 2870 2479 2926 2488
rect 2504 2100 2556 2106
rect 2504 2042 2556 2048
rect 2044 1420 2096 1426
rect 2044 1362 2096 1368
rect 2056 480 2084 1362
rect 2516 480 2544 2042
rect 2976 649 3004 6938
rect 3160 4842 3188 7126
rect 3252 5302 3280 8230
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3436 6458 3464 7890
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 3160 4814 3280 4842
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3160 4010 3188 4626
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3160 3534 3188 3946
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 3068 3194 3096 3470
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 3252 3058 3280 4814
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3054 2816 3110 2825
rect 3054 2751 3110 2760
rect 2962 640 3018 649
rect 2962 575 3018 584
rect 3068 480 3096 2751
rect 3344 1601 3372 6122
rect 3528 2990 3556 9454
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3620 8634 3648 8910
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3620 7002 3648 7142
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3712 6186 3740 12378
rect 3804 12102 3832 15014
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3804 9518 3832 11494
rect 3896 9586 3924 15558
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3988 13433 4016 15506
rect 4080 15162 4108 20567
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 11348 19802 11376 22320
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 11164 19774 11376 19802
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 6736 19236 6788 19242
rect 6736 19178 6788 19184
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4080 13802 4108 13874
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 3974 13424 4030 13433
rect 3974 13359 4030 13368
rect 3988 12424 4016 13359
rect 4080 12986 4108 13738
rect 4172 13326 4200 13806
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4172 12782 4200 13262
rect 4160 12776 4212 12782
rect 4066 12744 4122 12753
rect 4160 12718 4212 12724
rect 4066 12679 4068 12688
rect 4120 12679 4122 12688
rect 4068 12650 4120 12656
rect 4160 12436 4212 12442
rect 3988 12396 4160 12424
rect 4160 12378 4212 12384
rect 3974 12336 4030 12345
rect 3974 12271 4030 12280
rect 3988 11898 4016 12271
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4080 11393 4108 11630
rect 4066 11384 4122 11393
rect 4066 11319 4122 11328
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 4066 10840 4122 10849
rect 4172 10826 4200 11222
rect 4122 10798 4200 10826
rect 4066 10775 4122 10784
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 3976 10532 4028 10538
rect 3976 10474 4028 10480
rect 3988 10033 4016 10474
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 4080 10266 4108 10367
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4172 10130 4200 10542
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 3974 10024 4030 10033
rect 3974 9959 4030 9968
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3792 9512 3844 9518
rect 4080 9489 4108 9862
rect 4264 9654 4292 15506
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4356 13462 4384 13670
rect 4632 13530 4660 13670
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4344 13456 4396 13462
rect 4344 13398 4396 13404
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4344 12300 4396 12306
rect 4540 12288 4568 12378
rect 4396 12260 4568 12288
rect 4344 12242 4396 12248
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4724 11898 4752 12174
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4816 11665 4844 12106
rect 4802 11656 4858 11665
rect 4802 11591 4858 11600
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4816 9586 4844 11018
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 3792 9454 3844 9460
rect 3882 9480 3938 9489
rect 3882 9415 3938 9424
rect 4066 9480 4122 9489
rect 4066 9415 4122 9424
rect 4712 9444 4764 9450
rect 3896 8566 3924 9415
rect 4712 9386 4764 9392
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4080 9178 4108 9318
rect 4724 9178 4752 9386
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4066 9072 4122 9081
rect 4066 9007 4122 9016
rect 4252 9036 4304 9042
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3884 8560 3936 8566
rect 3988 8537 4016 8842
rect 4080 8838 4108 9007
rect 4252 8978 4304 8984
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3884 8502 3936 8508
rect 3974 8528 4030 8537
rect 3792 8492 3844 8498
rect 3974 8463 4030 8472
rect 3792 8434 3844 8440
rect 3804 8294 3832 8434
rect 3974 8392 4030 8401
rect 3974 8327 4030 8336
rect 3988 8294 4016 8327
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3804 7886 3832 8230
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 3804 6118 3832 7686
rect 4264 7546 4292 8978
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4434 8392 4490 8401
rect 4434 8327 4490 8336
rect 4448 8294 4476 8327
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4816 7818 4844 8910
rect 4908 8022 4936 14418
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 5092 12986 5120 13670
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5184 12374 5212 12582
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5000 9636 5028 12038
rect 5092 10130 5120 12174
rect 5276 12102 5304 12718
rect 5264 12096 5316 12102
rect 5368 12073 5396 14826
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5264 12038 5316 12044
rect 5354 12064 5410 12073
rect 5354 11999 5410 12008
rect 5368 11626 5396 11999
rect 5552 11762 5580 13126
rect 5540 11756 5592 11762
rect 5460 11716 5540 11744
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5276 11354 5304 11494
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5460 10606 5488 11716
rect 5540 11698 5592 11704
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5000 9608 5111 9636
rect 5083 9602 5111 9608
rect 5083 9574 5120 9602
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 5000 8090 5028 8230
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 3974 7168 4030 7177
rect 3974 7103 4030 7112
rect 3988 6934 4016 7103
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6225 4108 6598
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3698 5672 3754 5681
rect 3698 5607 3754 5616
rect 3712 3913 3740 5607
rect 3804 5166 3832 5850
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 4080 5574 4108 5743
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3882 5264 3938 5273
rect 3882 5199 3938 5208
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3896 4826 3924 5199
rect 3988 4865 4016 5306
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3974 4856 4030 4865
rect 3884 4820 3936 4826
rect 3974 4791 4030 4800
rect 3884 4762 3936 4768
rect 3790 4720 3846 4729
rect 3790 4655 3846 4664
rect 3698 3904 3754 3913
rect 3698 3839 3754 3848
rect 3804 3466 3832 4655
rect 4080 4321 4108 5034
rect 4066 4312 4122 4321
rect 4066 4247 4122 4256
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3738 4108 3878
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3516 2984 3568 2990
rect 3436 2944 3516 2972
rect 3436 2009 3464 2944
rect 3516 2926 3568 2932
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3422 2000 3478 2009
rect 3422 1935 3478 1944
rect 3330 1592 3386 1601
rect 3330 1527 3386 1536
rect 3528 480 3556 2790
rect 3620 1057 3648 2994
rect 3896 2854 3924 3130
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3606 1048 3662 1057
rect 3606 983 3662 992
rect 3988 480 4016 3334
rect 4068 2984 4120 2990
rect 4066 2952 4068 2961
rect 4120 2952 4122 2961
rect 4066 2887 4122 2896
rect 4172 2854 4200 3538
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4264 1442 4292 7278
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4724 5914 4752 7142
rect 4908 7002 4936 7958
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 5000 7721 5028 7890
rect 4986 7712 5042 7721
rect 4986 7647 5042 7656
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4816 6118 4844 6190
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4816 5778 4844 6054
rect 4804 5772 4856 5778
rect 4724 5732 4804 5760
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4724 5030 4752 5732
rect 4804 5714 4856 5720
rect 4712 5024 4764 5030
rect 5092 4978 5120 9574
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5184 8498 5212 9454
rect 5262 8936 5318 8945
rect 5262 8871 5318 8880
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7886 5212 8230
rect 5276 8022 5304 8871
rect 5368 8090 5396 9454
rect 5460 8498 5488 10542
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5264 8016 5316 8022
rect 5316 7964 5396 7970
rect 5264 7958 5396 7964
rect 5276 7942 5396 7958
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5184 7410 5212 7822
rect 5276 7585 5304 7822
rect 5262 7576 5318 7585
rect 5262 7511 5318 7520
rect 5262 7440 5318 7449
rect 5172 7404 5224 7410
rect 5262 7375 5318 7384
rect 5172 7346 5224 7352
rect 5276 7342 5304 7375
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5368 5114 5396 7942
rect 5460 7818 5488 8434
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5460 7410 5488 7754
rect 5552 7546 5580 11154
rect 5644 11150 5672 14962
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5736 12986 5764 13738
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5828 11626 5856 16594
rect 6000 14952 6052 14958
rect 6000 14894 6052 14900
rect 6012 14550 6040 14894
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6104 12782 6132 13126
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6196 12628 6224 18770
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6104 12600 6224 12628
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5828 11257 5856 11562
rect 5814 11248 5870 11257
rect 5814 11183 5870 11192
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5644 10470 5672 10950
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5644 10198 5672 10406
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5644 9654 5672 10134
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5736 9926 5764 10066
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5736 9586 5764 9862
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5828 9466 5856 11086
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 6012 10062 6040 10678
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 5906 9616 5962 9625
rect 5906 9551 5962 9560
rect 5644 9438 5856 9466
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5460 6866 5488 7210
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5460 5914 5488 6598
rect 5552 6458 5580 6598
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5552 5710 5580 6122
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5368 5086 5488 5114
rect 4712 4966 4764 4972
rect 4724 4706 4752 4966
rect 4632 4690 4752 4706
rect 4620 4684 4752 4690
rect 4672 4678 4752 4684
rect 4620 4626 4672 4632
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4724 4282 4752 4678
rect 4908 4950 5120 4978
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4540 3738 4568 3878
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4356 2650 4384 2790
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4264 1414 4476 1442
rect 4448 480 4476 1414
rect 4908 480 4936 4950
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5276 4146 5304 4422
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5276 3466 5304 4082
rect 5368 4078 5396 4966
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5460 3602 5488 5086
rect 5644 5030 5672 9438
rect 5920 9382 5948 9551
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5828 8634 5856 9318
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4554 5672 4966
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 3058 5304 3402
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5368 480 5396 2790
rect 202 0 258 480
rect 662 0 718 480
rect 1122 0 1178 480
rect 1582 0 1638 480
rect 2042 0 2098 480
rect 2502 0 2558 480
rect 3054 0 3110 480
rect 3514 0 3570 480
rect 3974 0 4030 480
rect 4434 0 4490 480
rect 4894 0 4950 480
rect 5354 0 5410 480
rect 5460 241 5488 3538
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5552 3369 5580 3470
rect 5736 3398 5764 3946
rect 5724 3392 5776 3398
rect 5538 3360 5594 3369
rect 5724 3334 5776 3340
rect 5538 3295 5594 3304
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5644 3058 5672 3130
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5828 2990 5856 8230
rect 5920 7002 5948 9318
rect 6012 9042 6040 9998
rect 6104 9659 6132 12600
rect 6090 9650 6146 9659
rect 6090 9585 6146 9594
rect 6184 9444 6236 9450
rect 6184 9386 6236 9392
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 6196 8498 6224 9386
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6288 8344 6316 14010
rect 6380 11354 6408 17682
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 6656 13530 6684 13670
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6472 12442 6500 12786
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6472 8362 6500 12242
rect 6656 11801 6684 12718
rect 6642 11792 6698 11801
rect 6642 11727 6698 11736
rect 6656 10674 6684 11727
rect 6748 11014 6776 19178
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 7024 14074 7052 14418
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7012 13796 7064 13802
rect 7012 13738 7064 13744
rect 7024 13530 7052 13738
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 7024 12442 7052 13194
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7102 11792 7158 11801
rect 7102 11727 7104 11736
rect 7156 11727 7158 11736
rect 7208 11744 7236 17070
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 7300 12238 7328 12650
rect 7392 12306 7420 17614
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7576 13870 7604 14962
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7668 13938 7696 14554
rect 11164 14550 11192 19774
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 16580 18148 16632 18154
rect 16580 18090 16632 18096
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13740 15638 13768 15982
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7484 13530 7512 13670
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7208 11716 7328 11744
rect 7104 11698 7156 11704
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6460 8356 6512 8362
rect 6288 8316 6408 8344
rect 5998 7304 6054 7313
rect 5998 7239 6054 7248
rect 6012 7206 6040 7239
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5920 6458 5948 6734
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 5920 480 5948 3334
rect 6012 2854 6040 7142
rect 6380 6866 6408 8316
rect 6460 8298 6512 8304
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6564 8090 6592 8298
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6288 5846 6316 6054
rect 6380 5846 6408 6802
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6104 2990 6132 4762
rect 6196 4758 6224 5170
rect 6472 5098 6500 6598
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 6196 4146 6224 4694
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6656 4010 6684 8230
rect 6748 5166 6776 10950
rect 6840 8634 6868 11154
rect 7116 11150 7144 11494
rect 7300 11218 7328 11716
rect 7576 11354 7604 13806
rect 7760 13326 7788 14486
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 8208 13456 8260 13462
rect 8300 13456 8352 13462
rect 8208 13398 8260 13404
rect 8298 13424 8300 13433
rect 8352 13424 8354 13433
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7760 12986 7788 13262
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 6932 9654 6960 11086
rect 7116 10810 7144 11086
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 7392 9586 7420 11018
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7484 9586 7512 10474
rect 7576 10266 7604 11086
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7668 10266 7696 10542
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7656 10260 7708 10266
rect 7760 10248 7788 12582
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 8220 12442 8248 13398
rect 8298 13359 8354 13368
rect 8680 13326 8708 14214
rect 10060 13394 10088 14282
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10336 13870 10364 14214
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8680 12850 8708 13262
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8496 12442 8524 12582
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8680 12306 8708 12786
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8220 11898 8248 12174
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8404 11558 8432 12242
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8220 11082 8248 11154
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8496 10606 8524 12242
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8588 11898 8616 12174
rect 8772 11898 8800 13330
rect 10060 12986 10088 13330
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 9220 12368 9272 12374
rect 9220 12310 9272 12316
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8588 11762 8616 11834
rect 8864 11801 8892 12038
rect 8850 11792 8906 11801
rect 8576 11756 8628 11762
rect 8850 11727 8906 11736
rect 8576 11698 8628 11704
rect 8864 10674 8892 11727
rect 8852 10668 8904 10674
rect 8680 10628 8852 10656
rect 8484 10600 8536 10606
rect 8404 10560 8484 10588
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7760 10220 7880 10248
rect 7656 10202 7708 10208
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6840 7546 6868 8366
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6932 7478 6960 7686
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6932 7002 6960 7414
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7024 6798 7052 8502
rect 7208 7886 7236 8978
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7208 7410 7236 7822
rect 7300 7546 7328 9318
rect 7484 8906 7512 9522
rect 7576 9042 7604 10202
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7484 8514 7512 8842
rect 7668 8634 7696 8910
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7760 8566 7788 10066
rect 7852 9586 7880 10220
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7944 9722 7972 9998
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 7748 8560 7800 8566
rect 7484 8498 7604 8514
rect 7748 8502 7800 8508
rect 7484 8492 7616 8498
rect 7484 8486 7564 8492
rect 7564 8434 7616 8440
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6840 4758 6868 6190
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7024 4826 7052 5510
rect 7116 5234 7144 6870
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7208 5137 7236 6326
rect 7194 5128 7250 5137
rect 7194 5063 7250 5072
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6828 4752 6880 4758
rect 7208 4706 7236 5063
rect 6828 4694 6880 4700
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6182 3632 6238 3641
rect 6182 3567 6238 3576
rect 6196 3058 6224 3567
rect 6288 3194 6316 3878
rect 6840 3618 6868 4694
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 7024 4678 7236 4706
rect 6932 3738 6960 4626
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6840 3590 6960 3618
rect 6828 3528 6880 3534
rect 6366 3496 6422 3505
rect 6828 3470 6880 3476
rect 6366 3431 6422 3440
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6380 480 6408 3431
rect 6840 2990 6868 3470
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6932 2666 6960 3590
rect 7024 2825 7052 4678
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7116 2990 7144 4558
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7208 4078 7236 4422
rect 7300 4162 7328 6938
rect 7392 4282 7420 8298
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8116 7336 8168 7342
rect 8220 7324 8248 8978
rect 8312 8974 8340 9386
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8168 7296 8248 7324
rect 8116 7278 8168 7284
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7484 4826 7512 7142
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7576 6662 7604 6870
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 7838 6760 7894 6769
rect 7838 6695 7894 6704
rect 7852 6662 7880 6695
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7760 6322 7788 6598
rect 8036 6390 8064 6802
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8024 6384 8076 6390
rect 8024 6326 8076 6332
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 8128 6254 8156 6666
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7760 5914 7788 6054
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 8220 5574 8248 6326
rect 8312 5846 8340 6734
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7300 4134 7420 4162
rect 7576 4146 7604 5102
rect 8220 5098 8248 5510
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7010 2816 7066 2825
rect 7010 2751 7066 2760
rect 6840 2638 6960 2666
rect 6840 480 6868 2638
rect 7208 1426 7236 3606
rect 7196 1420 7248 1426
rect 7196 1362 7248 1368
rect 7300 480 7328 4014
rect 7392 1306 7420 4134
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7484 3602 7512 4082
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7576 2650 7604 3946
rect 7760 3398 7788 4762
rect 8220 4622 8248 5034
rect 8312 4826 8340 5646
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8404 4706 8432 10560
rect 8484 10542 8536 10548
rect 8680 9722 8708 10628
rect 8852 10610 8904 10616
rect 8956 10266 8984 12242
rect 9232 12073 9260 12310
rect 10244 12238 10272 12650
rect 9404 12232 9456 12238
rect 10048 12232 10100 12238
rect 9404 12174 9456 12180
rect 10046 12200 10048 12209
rect 10232 12232 10284 12238
rect 10100 12200 10102 12209
rect 9218 12064 9274 12073
rect 9218 11999 9274 12008
rect 9416 11937 9444 12174
rect 10232 12174 10284 12180
rect 10046 12135 10102 12144
rect 10244 12102 10272 12174
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 9402 11928 9458 11937
rect 9036 11892 9088 11898
rect 9402 11863 9458 11872
rect 9036 11834 9088 11840
rect 9048 11694 9076 11834
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9128 11280 9180 11286
rect 9126 11248 9128 11257
rect 9180 11248 9182 11257
rect 9126 11183 9182 11192
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9494 11112 9550 11121
rect 9494 11047 9550 11056
rect 9508 11014 9536 11047
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9692 10266 9720 11154
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9784 10538 9812 11086
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9508 9722 9536 10066
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 9496 9716 9548 9722
rect 9692 9704 9720 10066
rect 9784 9926 9812 10474
rect 9968 10130 9996 11630
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10232 11144 10284 11150
rect 10428 11132 10456 12786
rect 10600 12368 10652 12374
rect 10598 12336 10600 12345
rect 10652 12336 10654 12345
rect 10598 12271 10654 12280
rect 10704 11898 10732 14418
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10796 12442 10824 14350
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11624 13938 11652 14894
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 10980 13530 11008 13874
rect 12452 13870 12480 14418
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 11256 13530 11284 13806
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 10980 12782 11008 13466
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 11164 12238 11192 13126
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10520 11801 10548 11834
rect 11072 11830 11100 12038
rect 11164 11898 11192 12174
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 10600 11824 10652 11830
rect 10506 11792 10562 11801
rect 10600 11766 10652 11772
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 11150 11792 11206 11801
rect 10506 11727 10562 11736
rect 10508 11144 10560 11150
rect 10428 11104 10508 11132
rect 10232 11086 10284 11092
rect 10508 11086 10560 11092
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9968 9722 9996 9930
rect 9956 9716 10008 9722
rect 9692 9676 9812 9704
rect 9496 9658 9548 9664
rect 8680 9586 8708 9658
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8484 9172 8536 9178
rect 8588 9160 8616 9522
rect 8588 9132 8708 9160
rect 8484 9114 8536 9120
rect 8496 8498 8524 9114
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8588 8945 8616 8978
rect 8574 8936 8630 8945
rect 8574 8871 8630 8880
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8482 8392 8538 8401
rect 8482 8327 8538 8336
rect 8496 6254 8524 8327
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8588 4758 8616 6054
rect 8312 4678 8432 4706
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 8128 3194 8156 3470
rect 8220 3398 8248 3946
rect 8312 3505 8340 4678
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8298 3496 8354 3505
rect 8298 3431 8354 3440
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 8220 2582 8248 3334
rect 8404 2922 8432 4014
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 8496 2378 8524 3334
rect 8588 3194 8616 3538
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 8680 2038 8708 9132
rect 8772 8974 8800 9658
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 8022 8984 8434
rect 9324 8090 9352 9386
rect 9416 8634 9444 9386
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9508 8022 9536 8774
rect 8944 8016 8996 8022
rect 8944 7958 8996 7964
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 8956 7546 8984 7958
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 8772 6730 8800 7414
rect 9048 7410 9076 7890
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 7721 9168 7822
rect 9126 7712 9182 7721
rect 9126 7647 9182 7656
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8208 2032 8260 2038
rect 8208 1974 8260 1980
rect 8668 2032 8720 2038
rect 8668 1974 8720 1980
rect 7392 1278 7788 1306
rect 7760 480 7788 1278
rect 8220 480 8248 1974
rect 8772 480 8800 6666
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8956 5930 8984 6054
rect 8864 5902 8984 5930
rect 8864 4729 8892 5902
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8956 5370 8984 5646
rect 9048 5642 9076 7346
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 9048 5370 9076 5578
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8850 4720 8906 4729
rect 8850 4655 8906 4664
rect 8864 4010 8892 4655
rect 9048 4078 9076 5306
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 8956 2854 8984 3674
rect 9140 3194 9168 7278
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 7002 9720 7142
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9232 6322 9260 6734
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9232 4554 9260 6258
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9232 4282 9260 4490
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9600 3534 9628 4014
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 8956 2106 8984 2790
rect 9324 2666 9352 3130
rect 9600 3058 9628 3470
rect 9692 3126 9720 6190
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9784 2972 9812 9676
rect 9956 9658 10008 9664
rect 10152 8634 10180 11086
rect 10244 10810 10272 11086
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10428 10810 10456 10950
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10230 10568 10286 10577
rect 10230 10503 10286 10512
rect 10244 10470 10272 10503
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10428 10180 10456 10746
rect 10520 10606 10548 11086
rect 10612 10713 10640 11766
rect 11150 11727 11206 11736
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10598 10704 10654 10713
rect 10598 10639 10654 10648
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10692 10192 10744 10198
rect 10428 10152 10692 10180
rect 10692 10134 10744 10140
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10244 8566 10272 9862
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10060 8090 10088 8502
rect 10428 8498 10456 9318
rect 10612 9042 10640 9454
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10704 8922 10732 9454
rect 10612 8894 10732 8922
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10152 7410 10180 7822
rect 10244 7546 10272 8230
rect 10336 7857 10364 8230
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10322 7848 10378 7857
rect 10322 7783 10378 7792
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 6458 10088 6802
rect 10336 6798 10364 7414
rect 10428 7206 10456 8026
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10152 6458 10180 6734
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10140 6452 10192 6458
rect 10520 6440 10548 8570
rect 10612 7970 10640 8894
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10704 8090 10732 8298
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10612 7942 10732 7970
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10612 7478 10640 7686
rect 10600 7472 10652 7478
rect 10600 7414 10652 7420
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10140 6394 10192 6400
rect 10428 6412 10548 6440
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9876 3738 9904 6054
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9968 3602 9996 4558
rect 10060 3670 10088 4626
rect 10152 4298 10180 6122
rect 10428 6118 10456 6412
rect 10612 6322 10640 7278
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10520 6225 10548 6258
rect 10506 6216 10562 6225
rect 10506 6151 10562 6160
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10152 4282 10272 4298
rect 10152 4276 10284 4282
rect 10152 4270 10232 4276
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9232 2638 9352 2666
rect 9692 2944 9812 2972
rect 8944 2100 8996 2106
rect 8944 2042 8996 2048
rect 9232 480 9260 2638
rect 9692 480 9720 2944
rect 9876 2650 9904 3538
rect 9968 2854 9996 3538
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 10152 480 10180 4270
rect 10232 4218 10284 4224
rect 10336 4078 10364 5102
rect 10324 4072 10376 4078
rect 10428 4049 10456 6054
rect 10598 5128 10654 5137
rect 10598 5063 10600 5072
rect 10652 5063 10654 5072
rect 10600 5034 10652 5040
rect 10598 4720 10654 4729
rect 10598 4655 10654 4664
rect 10612 4486 10640 4655
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 10324 4014 10376 4020
rect 10414 4040 10470 4049
rect 10414 3975 10470 3984
rect 10428 3210 10456 3975
rect 10336 3182 10456 3210
rect 10336 2650 10364 3182
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10428 2446 10456 2790
rect 10612 2582 10640 4422
rect 10704 4010 10732 7942
rect 10796 7177 10824 11494
rect 10980 11354 11008 11630
rect 11164 11558 11192 11727
rect 11716 11694 11744 12174
rect 11808 12170 11836 13330
rect 12452 13326 12480 13806
rect 12912 13518 13124 13546
rect 12808 13456 12860 13462
rect 12806 13424 12808 13433
rect 12860 13424 12862 13433
rect 12912 13394 12940 13518
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 12806 13359 12862 13368
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11704 11688 11756 11694
rect 11610 11656 11666 11665
rect 11704 11630 11756 11636
rect 11610 11591 11666 11600
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11624 11506 11652 11591
rect 11624 11478 11744 11506
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 10888 9382 10916 11222
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11072 9654 11100 11018
rect 11164 10690 11192 11222
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11164 10662 11284 10690
rect 11256 10470 11284 10662
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 11164 8634 11192 10066
rect 11256 10062 11284 10406
rect 11624 10130 11652 10746
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 10874 8528 10930 8537
rect 10874 8463 10930 8472
rect 11152 8492 11204 8498
rect 10782 7168 10838 7177
rect 10782 7103 10838 7112
rect 10888 6390 10916 8463
rect 11152 8434 11204 8440
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 11072 8090 11100 8298
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10980 7342 11008 7890
rect 11058 7576 11114 7585
rect 11058 7511 11060 7520
rect 11112 7511 11114 7520
rect 11060 7482 11112 7488
rect 11164 7410 11192 8434
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11520 7472 11572 7478
rect 11518 7440 11520 7449
rect 11572 7440 11574 7449
rect 11152 7404 11204 7410
rect 11518 7375 11574 7384
rect 11152 7346 11204 7352
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 6866 11100 7142
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11072 6662 11100 6802
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10980 5914 11008 6258
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10784 5840 10836 5846
rect 10782 5808 10784 5817
rect 10836 5808 10838 5817
rect 11164 5760 11192 7346
rect 11624 6934 11652 7890
rect 11612 6928 11664 6934
rect 11612 6870 11664 6876
rect 11426 6760 11482 6769
rect 11426 6695 11428 6704
rect 11480 6695 11482 6704
rect 11428 6666 11480 6672
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11624 6186 11652 6394
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11716 6118 11744 11478
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 10782 5743 10838 5752
rect 10980 5732 11192 5760
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10690 3360 10746 3369
rect 10690 3295 10746 3304
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 10416 2440 10468 2446
rect 10704 2428 10732 3295
rect 10796 2922 10824 4966
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10888 2446 10916 5510
rect 10980 2972 11008 5732
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11256 4758 11284 5034
rect 11348 4758 11376 5170
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11518 4992 11574 5001
rect 11440 4826 11468 4966
rect 11518 4927 11574 4936
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11532 4690 11560 4927
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4282 11100 4422
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3670 11468 3878
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11072 3097 11100 3334
rect 11058 3088 11114 3097
rect 11058 3023 11114 3032
rect 11164 2990 11192 3334
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11152 2984 11204 2990
rect 10980 2944 11100 2972
rect 10416 2382 10468 2388
rect 10612 2400 10732 2428
rect 10876 2440 10928 2446
rect 10612 480 10640 2400
rect 10876 2382 10928 2388
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 2106 11008 2246
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 11072 480 11100 2944
rect 11152 2926 11204 2932
rect 11624 2650 11652 3470
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11716 2038 11744 2382
rect 11704 2032 11756 2038
rect 11704 1974 11756 1980
rect 11808 1850 11836 11834
rect 12084 11257 12112 12242
rect 12348 12096 12400 12102
rect 12452 12084 12480 13262
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12624 12232 12676 12238
rect 12622 12200 12624 12209
rect 12676 12200 12678 12209
rect 12622 12135 12678 12144
rect 12400 12056 12480 12084
rect 12348 12038 12400 12044
rect 12070 11248 12126 11257
rect 12452 11218 12480 12056
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12070 11183 12126 11192
rect 12440 11212 12492 11218
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11992 9761 12020 10066
rect 11978 9752 12034 9761
rect 11978 9687 12034 9696
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11900 8430 11928 8774
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11888 8016 11940 8022
rect 11992 7993 12020 9687
rect 11888 7958 11940 7964
rect 11978 7984 12034 7993
rect 11900 7206 11928 7958
rect 11978 7919 12034 7928
rect 12084 7868 12112 11183
rect 12440 11154 12492 11160
rect 12452 10606 12480 11154
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12452 10130 12480 10542
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12164 8968 12216 8974
rect 12162 8936 12164 8945
rect 12216 8936 12218 8945
rect 12162 8871 12218 8880
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 11992 7840 12112 7868
rect 12268 7857 12296 8842
rect 12360 8498 12388 8978
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12452 8430 12480 8910
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12254 7848 12310 7857
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11900 5352 11928 7142
rect 11992 6934 12020 7840
rect 12254 7783 12310 7792
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 11900 5324 12020 5352
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11900 4758 11928 5170
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11888 3664 11940 3670
rect 11992 3641 12020 5324
rect 11888 3606 11940 3612
rect 11978 3632 12034 3641
rect 11900 3346 11928 3606
rect 11978 3567 12034 3576
rect 11900 3318 12020 3346
rect 11900 3058 11928 3318
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 11992 2038 12020 3318
rect 11980 2032 12032 2038
rect 11980 1974 12032 1980
rect 11624 1822 11836 1850
rect 11624 480 11652 1822
rect 12084 480 12112 7482
rect 12452 7290 12480 8366
rect 12544 8090 12572 12038
rect 12728 11218 12756 12242
rect 12912 11762 12940 12650
rect 13004 11937 13032 13398
rect 13096 12102 13124 13518
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 13188 12238 13216 12582
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12990 11928 13046 11937
rect 12990 11863 13046 11872
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12636 9994 12664 11086
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12728 10198 12756 10542
rect 12912 10452 12940 11494
rect 13004 11354 13032 11698
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13004 10606 13032 11290
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 12912 10424 13032 10452
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12900 9920 12952 9926
rect 12898 9888 12900 9897
rect 12952 9888 12954 9897
rect 12898 9823 12954 9832
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12624 9104 12676 9110
rect 12912 9081 12940 9386
rect 12624 9046 12676 9052
rect 12898 9072 12954 9081
rect 12636 8786 12664 9046
rect 12898 9007 12954 9016
rect 12636 8758 12756 8786
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12636 8090 12664 8570
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12622 7984 12678 7993
rect 12728 7954 12756 8758
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12622 7919 12624 7928
rect 12676 7919 12678 7928
rect 12716 7948 12768 7954
rect 12624 7890 12676 7896
rect 12716 7890 12768 7896
rect 12820 7886 12848 8298
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12360 7262 12480 7290
rect 12624 7268 12676 7274
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12176 6254 12204 6870
rect 12256 6656 12308 6662
rect 12360 6644 12388 7262
rect 12624 7210 12676 7216
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12308 6616 12388 6644
rect 12256 6598 12308 6604
rect 12360 6390 12388 6616
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12360 5778 12388 6326
rect 12452 5914 12480 7142
rect 12530 6760 12586 6769
rect 12530 6695 12532 6704
rect 12584 6695 12586 6704
rect 12532 6666 12584 6672
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12360 4486 12388 5714
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12544 5370 12572 5646
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12636 4185 12664 7210
rect 12808 7200 12860 7206
rect 12912 7177 12940 8298
rect 12808 7142 12860 7148
rect 12898 7168 12954 7177
rect 12820 7002 12848 7142
rect 12898 7103 12954 7112
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12820 6254 12848 6598
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12820 5710 12848 6190
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12912 5386 12940 7103
rect 13004 6848 13032 10424
rect 13280 9654 13308 15506
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13648 13530 13676 14758
rect 14016 13938 14044 14758
rect 14384 14278 14412 14962
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 14384 13870 14412 14214
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 14200 13462 14228 13670
rect 13452 13456 13504 13462
rect 13452 13398 13504 13404
rect 14188 13456 14240 13462
rect 14188 13398 14240 13404
rect 13464 13258 13492 13398
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13464 12850 13492 13194
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 14292 12782 14320 13126
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13832 12442 13860 12582
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13452 12232 13504 12238
rect 13504 12180 13584 12186
rect 13452 12174 13584 12180
rect 13464 12158 13584 12174
rect 13358 11928 13414 11937
rect 13358 11863 13360 11872
rect 13412 11863 13414 11872
rect 13360 11834 13412 11840
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13464 11354 13492 11698
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13096 9110 13124 9318
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 13188 7818 13216 9386
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13280 8090 13308 9318
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13280 7818 13308 7890
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13280 7698 13308 7754
rect 13188 7670 13308 7698
rect 13188 7206 13216 7670
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13280 7002 13308 7482
rect 13372 7410 13400 9862
rect 13450 9480 13506 9489
rect 13450 9415 13506 9424
rect 13464 8294 13492 9415
rect 13556 9042 13584 12158
rect 13924 11354 13952 12718
rect 14384 12306 14412 13806
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14384 11762 14412 12242
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13740 10470 13768 11086
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10198 13768 10406
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13832 9722 13860 10134
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13740 9382 13768 9590
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13464 7546 13492 7890
rect 13556 7546 13584 8978
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13740 7886 13768 8774
rect 13832 8634 13860 9522
rect 13924 8945 13952 9590
rect 14016 9586 14044 10066
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 14016 9178 14044 9386
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 13910 8936 13966 8945
rect 13910 8871 13966 8880
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13372 6866 13400 7346
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13360 6860 13412 6866
rect 13004 6820 13308 6848
rect 13082 6760 13138 6769
rect 13082 6695 13138 6704
rect 13096 6118 13124 6695
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 12992 5840 13044 5846
rect 13044 5800 13124 5828
rect 12992 5782 13044 5788
rect 12820 5358 12940 5386
rect 12820 5166 12848 5358
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12622 4176 12678 4185
rect 12544 4120 12622 4128
rect 12544 4111 12678 4120
rect 12544 4100 12664 4111
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12176 2582 12204 3878
rect 12438 3632 12494 3641
rect 12256 3596 12308 3602
rect 12308 3556 12388 3584
rect 12438 3567 12494 3576
rect 12256 3538 12308 3544
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 12268 2582 12296 2926
rect 12360 2825 12388 3556
rect 12346 2816 12402 2825
rect 12346 2751 12402 2760
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 12452 2514 12480 3567
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12544 480 12572 4100
rect 12636 4051 12664 4100
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12636 3602 12664 3946
rect 12820 3670 12848 4966
rect 12808 3664 12860 3670
rect 12808 3606 12860 3612
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12636 2496 12664 3402
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12728 2650 12756 3334
rect 12808 2984 12860 2990
rect 12912 2972 12940 5238
rect 12992 4752 13044 4758
rect 12992 4694 13044 4700
rect 13004 4486 13032 4694
rect 13096 4593 13124 5800
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13082 4584 13138 4593
rect 13082 4519 13138 4528
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 13004 4146 13032 4422
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13004 3534 13032 4082
rect 13096 4078 13124 4519
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13096 3738 13124 3878
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13082 3088 13138 3097
rect 13082 3023 13084 3032
rect 13136 3023 13138 3032
rect 13084 2994 13136 3000
rect 13188 2990 13216 5510
rect 12860 2944 12940 2972
rect 13176 2984 13228 2990
rect 12808 2926 12860 2932
rect 13176 2926 13228 2932
rect 12808 2848 12860 2854
rect 12806 2816 12808 2825
rect 13280 2836 13308 6820
rect 13360 6802 13412 6808
rect 13372 5234 13400 6802
rect 13464 6458 13492 7210
rect 13924 6798 13952 8871
rect 14016 8634 14044 9114
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13924 5846 13952 6394
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13464 4690 13492 5306
rect 13556 4690 13584 5714
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13648 4826 13676 4966
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13556 4078 13584 4626
rect 13740 4214 13768 4966
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 12860 2816 12862 2825
rect 12806 2751 12862 2760
rect 13004 2808 13308 2836
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12716 2508 12768 2514
rect 12636 2468 12716 2496
rect 12716 2450 12768 2456
rect 13004 480 13032 2808
rect 13464 480 13492 3062
rect 13740 2990 13768 3946
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13924 480 13952 2790
rect 14016 2514 14044 7686
rect 14108 5302 14136 11494
rect 14384 11150 14412 11698
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14200 10130 14228 11018
rect 14292 10810 14320 11086
rect 14476 10826 14504 14894
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 16592 14618 16620 18090
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14936 12850 14964 13126
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 15120 12646 15148 14418
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15396 13870 15424 14350
rect 16408 14074 16436 14418
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14832 12368 14884 12374
rect 14830 12336 14832 12345
rect 14884 12336 14886 12345
rect 14830 12271 14886 12280
rect 15014 12336 15070 12345
rect 15014 12271 15070 12280
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14660 11762 14688 12174
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 15028 11558 15056 12271
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14384 10798 14504 10826
rect 14278 10568 14334 10577
rect 14278 10503 14334 10512
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 14292 3738 14320 10503
rect 14384 7857 14412 10798
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14476 9110 14504 10610
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 15028 9178 15056 11154
rect 15120 10674 15148 12582
rect 15304 12322 15332 13330
rect 15396 12714 15424 13806
rect 15384 12708 15436 12714
rect 15436 12668 15516 12696
rect 15384 12650 15436 12656
rect 15304 12294 15424 12322
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15304 11898 15332 12174
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14370 7848 14426 7857
rect 14476 7818 14504 8026
rect 14370 7783 14426 7792
rect 14464 7812 14516 7818
rect 14464 7754 14516 7760
rect 14568 7342 14596 9114
rect 14646 9072 14702 9081
rect 14646 9007 14648 9016
rect 14700 9007 14702 9016
rect 14648 8978 14700 8984
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14844 7410 14872 7822
rect 15028 7478 15056 7890
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14384 6848 14412 7142
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14464 6860 14516 6866
rect 14384 6820 14464 6848
rect 14384 6186 14412 6820
rect 14464 6802 14516 6808
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14556 6384 14608 6390
rect 14556 6326 14608 6332
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14476 2990 14504 6054
rect 14568 5574 14596 6326
rect 14660 6322 14688 6598
rect 14844 6458 14872 6734
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14844 6322 14872 6394
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14648 5840 14700 5846
rect 14648 5782 14700 5788
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14568 4758 14596 5510
rect 14660 5234 14688 5782
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 15120 4690 15148 9998
rect 15212 8906 15240 11698
rect 15396 11540 15424 12294
rect 15304 11512 15424 11540
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15212 8022 15240 8502
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 15304 7426 15332 11512
rect 15488 11064 15516 12668
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15672 11558 15700 11834
rect 15764 11762 15792 12038
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15568 11076 15620 11082
rect 15488 11036 15568 11064
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15396 9722 15424 10066
rect 15488 10062 15516 11036
rect 15568 11018 15620 11024
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15474 9888 15530 9897
rect 15474 9823 15530 9832
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15212 7398 15332 7426
rect 15212 5273 15240 7398
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15304 7002 15332 7278
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15198 5264 15254 5273
rect 15198 5199 15254 5208
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14936 4214 14964 4422
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14936 4078 14964 4150
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14936 3924 14964 4014
rect 15212 3942 15240 5034
rect 15200 3936 15252 3942
rect 14936 3896 15056 3924
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 15028 3534 15056 3896
rect 15200 3878 15252 3884
rect 15212 3534 15240 3878
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15200 3528 15252 3534
rect 15396 3505 15424 8910
rect 15488 8106 15516 9823
rect 15580 9178 15608 10610
rect 15672 9654 15700 11086
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15764 10130 15792 10610
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8634 15884 8910
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15488 8078 15700 8106
rect 15568 8016 15620 8022
rect 15568 7958 15620 7964
rect 15474 7848 15530 7857
rect 15474 7783 15530 7792
rect 15488 6254 15516 7783
rect 15580 7410 15608 7958
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15672 6798 15700 8078
rect 15764 7002 15792 8230
rect 15856 8090 15884 8230
rect 15948 8090 15976 13806
rect 16302 13424 16358 13433
rect 16302 13359 16304 13368
rect 16356 13359 16358 13368
rect 16304 13330 16356 13336
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 16040 10470 16068 12242
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16224 11898 16252 12174
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16316 11393 16344 13330
rect 16408 13326 16436 14010
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16500 12442 16528 12854
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11898 16528 12106
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16396 11688 16448 11694
rect 16448 11636 16620 11642
rect 16396 11630 16620 11636
rect 16408 11626 16620 11630
rect 16408 11620 16632 11626
rect 16408 11614 16580 11620
rect 16580 11562 16632 11568
rect 16488 11552 16540 11558
rect 16540 11500 16620 11506
rect 16488 11494 16620 11500
rect 16500 11478 16620 11494
rect 16302 11384 16358 11393
rect 16302 11319 16358 11328
rect 16304 11280 16356 11286
rect 16302 11248 16304 11257
rect 16356 11248 16358 11257
rect 16212 11212 16264 11218
rect 16302 11183 16358 11192
rect 16212 11154 16264 11160
rect 16118 10976 16174 10985
rect 16118 10911 16174 10920
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 16040 10130 16068 10406
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 16040 6798 16068 7346
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 15672 6458 15700 6734
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5914 15608 6054
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15488 5681 15516 5714
rect 15474 5672 15530 5681
rect 15474 5607 15530 5616
rect 15856 5370 15884 6258
rect 16040 5370 16068 6734
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15764 3738 15792 3878
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15200 3470 15252 3476
rect 15382 3496 15438 3505
rect 15382 3431 15438 3440
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15384 3120 15436 3126
rect 15384 3062 15436 3068
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 14200 2378 14228 2926
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14476 480 14504 2246
rect 15028 1442 15056 2790
rect 14936 1414 15056 1442
rect 14936 480 14964 1414
rect 15396 480 15424 3062
rect 15488 2514 15516 3334
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15580 2446 15608 2926
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15856 480 15884 4422
rect 16132 4010 16160 10911
rect 16224 10810 16252 11154
rect 16486 11112 16542 11121
rect 16592 11082 16620 11478
rect 16486 11047 16542 11056
rect 16580 11076 16632 11082
rect 16500 11014 16528 11047
rect 16580 11018 16632 11024
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16316 10282 16344 10746
rect 16578 10704 16634 10713
rect 16488 10668 16540 10674
rect 16578 10639 16634 10648
rect 16488 10610 16540 10616
rect 16224 10254 16344 10282
rect 16224 9761 16252 10254
rect 16304 10192 16356 10198
rect 16304 10134 16356 10140
rect 16210 9752 16266 9761
rect 16316 9722 16344 10134
rect 16210 9687 16266 9696
rect 16304 9716 16356 9722
rect 16224 9178 16252 9687
rect 16304 9658 16356 9664
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16210 9072 16266 9081
rect 16210 9007 16266 9016
rect 16224 7426 16252 9007
rect 16316 7546 16344 9658
rect 16500 9586 16528 10610
rect 16592 10470 16620 10639
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16500 8974 16528 9522
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16592 8480 16620 8978
rect 16500 8452 16620 8480
rect 16500 8242 16528 8452
rect 16578 8392 16634 8401
rect 16578 8327 16580 8336
rect 16632 8327 16634 8336
rect 16580 8298 16632 8304
rect 16500 8214 16620 8242
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16224 7398 16344 7426
rect 16408 7410 16436 8026
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 16132 1986 16160 3402
rect 16224 2514 16252 7142
rect 16316 6254 16344 7398
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16304 5772 16356 5778
rect 16408 5760 16436 6938
rect 16500 6458 16528 7278
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16356 5732 16436 5760
rect 16304 5714 16356 5720
rect 16316 5166 16344 5714
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16316 3534 16344 5102
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16500 3602 16528 4762
rect 16592 4434 16620 8214
rect 16684 6458 16712 18770
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17040 14884 17092 14890
rect 17040 14826 17092 14832
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16776 13530 16804 13670
rect 16960 13530 16988 14758
rect 17052 13530 17080 14826
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16776 11354 16804 13126
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16868 11354 16896 11562
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16868 10266 16896 11086
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16776 8498 16804 10066
rect 16960 9024 16988 12242
rect 17052 11937 17080 13466
rect 17144 13190 17172 17682
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17132 12368 17184 12374
rect 17132 12310 17184 12316
rect 17038 11928 17094 11937
rect 17038 11863 17094 11872
rect 17144 11801 17172 12310
rect 17236 12102 17264 22471
rect 18970 22320 19026 22800
rect 18694 20632 18750 20641
rect 18694 20567 18750 20576
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18708 19514 18736 20567
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17880 18902 17908 19246
rect 17868 18896 17920 18902
rect 17868 18838 17920 18844
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18984 18154 19012 22320
rect 20258 22128 20314 22137
rect 20258 22063 20314 22072
rect 19982 20224 20038 20233
rect 19982 20159 20038 20168
rect 18972 18148 19024 18154
rect 18972 18090 19024 18096
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 17958 16960 18014 16969
rect 17958 16895 18014 16904
rect 17972 16250 18000 16895
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 17960 15088 18012 15094
rect 17958 15056 17960 15065
rect 18012 15056 18014 15065
rect 17958 14991 18014 15000
rect 19352 14958 19380 17070
rect 19890 16008 19946 16017
rect 19890 15943 19946 15952
rect 19904 15706 19932 15943
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17604 13938 17632 14486
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17420 13462 17448 13670
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17788 13326 17816 14350
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17972 12986 18000 13738
rect 18524 13462 18552 14214
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 17592 12708 17644 12714
rect 17592 12650 17644 12656
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17130 11792 17186 11801
rect 17130 11727 17186 11736
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17052 10713 17080 11494
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17038 10704 17094 10713
rect 17038 10639 17094 10648
rect 17144 10130 17172 11086
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17052 9110 17080 9318
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 16868 8996 16988 9024
rect 16868 8634 16896 8996
rect 17236 8906 17264 12038
rect 17328 9110 17356 12582
rect 17420 12238 17448 12582
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17420 11830 17448 12174
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 17224 8900 17276 8906
rect 17224 8842 17276 8848
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16776 7313 16804 8298
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16762 7304 16818 7313
rect 16762 7239 16818 7248
rect 16764 6928 16816 6934
rect 16764 6870 16816 6876
rect 16776 6730 16804 6870
rect 16868 6798 16896 7822
rect 16960 6798 16988 8842
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 17052 6610 17080 8230
rect 16960 6582 17080 6610
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16684 4554 16712 6122
rect 16960 5234 16988 6582
rect 17144 5930 17172 8366
rect 17236 8022 17264 8434
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17328 7410 17356 8502
rect 17420 8090 17448 8910
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17236 6662 17264 7142
rect 17420 7002 17448 8026
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17052 5902 17172 5930
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16776 4622 16804 4966
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16592 4406 16712 4434
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16684 2990 16712 4406
rect 16854 4176 16910 4185
rect 16854 4111 16910 4120
rect 16868 4078 16896 4111
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 17052 3942 17080 5902
rect 17224 5840 17276 5846
rect 17222 5808 17224 5817
rect 17276 5808 17278 5817
rect 17132 5772 17184 5778
rect 17222 5743 17278 5752
rect 17132 5714 17184 5720
rect 17144 4826 17172 5714
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17144 4690 17172 4762
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 17236 4010 17264 5743
rect 17328 5370 17356 6054
rect 17420 5710 17448 6938
rect 17512 6458 17540 8366
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17512 5234 17540 5510
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17512 5030 17540 5170
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17420 4146 17448 4626
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17224 4004 17276 4010
rect 17224 3946 17276 3952
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17604 3670 17632 12650
rect 18064 12442 18092 12718
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18156 12345 18184 12378
rect 18524 12374 18552 13398
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18616 12782 18644 13126
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18512 12368 18564 12374
rect 18142 12336 18198 12345
rect 17960 12300 18012 12306
rect 18512 12310 18564 12316
rect 18142 12271 18198 12280
rect 17960 12242 18012 12248
rect 17972 11898 18000 12242
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 18144 11824 18196 11830
rect 18144 11766 18196 11772
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 9178 17724 9318
rect 17880 9178 17908 11154
rect 18156 11082 18184 11766
rect 18524 11762 18552 12310
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18616 11642 18644 12718
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18524 11614 18644 11642
rect 18144 11076 18196 11082
rect 18144 11018 18196 11024
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18524 10606 18552 11614
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18328 10464 18380 10470
rect 17958 10432 18014 10441
rect 18380 10424 18552 10452
rect 18328 10406 18380 10412
rect 17958 10367 18014 10376
rect 17972 9722 18000 10367
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17960 9512 18012 9518
rect 17958 9480 17960 9489
rect 18012 9480 18014 9489
rect 17958 9415 18014 9424
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17696 8514 17724 9114
rect 17696 8486 17816 8514
rect 17880 8498 17908 9114
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17696 7002 17724 7686
rect 17684 6996 17736 7002
rect 17684 6938 17736 6944
rect 17788 6089 17816 8486
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17880 8022 17908 8230
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17880 7410 17908 7686
rect 17972 7410 18000 8978
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18524 8548 18552 10424
rect 18616 10033 18644 10950
rect 18602 10024 18658 10033
rect 18602 9959 18658 9968
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 18432 8520 18552 8548
rect 18432 8129 18460 8520
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18418 8120 18474 8129
rect 18418 8055 18474 8064
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18524 7546 18552 8230
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18524 7002 18552 7142
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 17774 6080 17830 6089
rect 17774 6015 17830 6024
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 17316 2984 17368 2990
rect 17604 2961 17632 3606
rect 17788 3466 17816 4694
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17316 2926 17368 2932
rect 17590 2952 17646 2961
rect 16304 2916 16356 2922
rect 16304 2858 16356 2864
rect 16316 2514 16344 2858
rect 17328 2582 17356 2926
rect 17590 2887 17646 2896
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17316 2576 17368 2582
rect 17316 2518 17368 2524
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 16304 2508 16356 2514
rect 16304 2450 16356 2456
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16132 1958 16344 1986
rect 16316 480 16344 1958
rect 16776 480 16804 2246
rect 17420 1442 17448 2790
rect 17880 2446 17908 6938
rect 18616 6934 18644 9862
rect 18604 6928 18656 6934
rect 18604 6870 18656 6876
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18432 5914 18460 6258
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 17958 5808 18014 5817
rect 17958 5743 18014 5752
rect 17972 4729 18000 5743
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 18052 5296 18104 5302
rect 18052 5238 18104 5244
rect 17958 4720 18014 4729
rect 17958 4655 18014 4664
rect 18064 4570 18092 5238
rect 17972 4542 18092 4570
rect 17972 4010 18000 4542
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18248 3505 18276 3878
rect 18340 3534 18368 4014
rect 18418 3768 18474 3777
rect 18418 3703 18420 3712
rect 18472 3703 18474 3712
rect 18420 3674 18472 3680
rect 18328 3528 18380 3534
rect 18234 3496 18290 3505
rect 18328 3470 18380 3476
rect 18234 3431 18290 3440
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18524 2514 18552 6802
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18616 4457 18644 6394
rect 18708 5370 18736 12650
rect 18800 6866 18828 13806
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18892 13530 18920 13670
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18892 12986 18920 13466
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18880 12232 18932 12238
rect 18984 12209 19012 14350
rect 19260 14113 19288 14758
rect 19246 14104 19302 14113
rect 19246 14039 19302 14048
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 19156 13728 19208 13734
rect 19154 13696 19156 13705
rect 19208 13696 19210 13705
rect 19154 13631 19210 13640
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 19168 12782 19196 13126
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19168 12306 19196 12718
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 18880 12174 18932 12180
rect 18970 12200 19026 12209
rect 18892 11694 18920 12174
rect 18970 12135 19026 12144
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18984 11626 19012 12135
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 18892 9178 18920 11018
rect 18972 9376 19024 9382
rect 18970 9344 18972 9353
rect 19024 9344 19026 9353
rect 18970 9279 19026 9288
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 19076 9042 19104 11018
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 19168 10062 19196 10406
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19168 9450 19196 9998
rect 19156 9444 19208 9450
rect 19156 9386 19208 9392
rect 19064 9036 19116 9042
rect 19260 9024 19288 13806
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19352 9518 19380 13126
rect 19444 12209 19472 15506
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19720 13938 19748 14894
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19430 12200 19486 12209
rect 19812 12170 19840 15506
rect 19890 14648 19946 14657
rect 19996 14618 20024 20159
rect 20166 19272 20222 19281
rect 20166 19207 20222 19216
rect 20180 17338 20208 19207
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 20074 15600 20130 15609
rect 20074 15535 20130 15544
rect 19890 14583 19892 14592
rect 19944 14583 19946 14592
rect 19984 14612 20036 14618
rect 19892 14554 19944 14560
rect 19984 14554 20036 14560
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 19892 14340 19944 14346
rect 19892 14282 19944 14288
rect 19430 12135 19486 12144
rect 19800 12164 19852 12170
rect 19800 12106 19852 12112
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19444 11558 19472 12038
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19536 11354 19564 12038
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 9654 19472 11086
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19536 9654 19564 10542
rect 19720 10470 19748 11630
rect 19904 11234 19932 14282
rect 19996 12442 20024 14418
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19982 12200 20038 12209
rect 19982 12135 20038 12144
rect 19812 11206 19932 11234
rect 19812 10810 19840 11206
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19812 10044 19840 10610
rect 19904 10470 19932 11086
rect 19996 10674 20024 12135
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 10198 19932 10406
rect 19892 10192 19944 10198
rect 19892 10134 19944 10140
rect 19812 10016 19932 10044
rect 19614 9752 19670 9761
rect 19614 9687 19670 9696
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19064 8978 19116 8984
rect 19168 8996 19288 9024
rect 19168 8922 19196 8996
rect 19340 8968 19392 8974
rect 19076 8894 19196 8922
rect 19246 8936 19302 8945
rect 18880 8628 18932 8634
rect 18932 8588 19012 8616
rect 18880 8570 18932 8576
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 18788 6724 18840 6730
rect 18788 6666 18840 6672
rect 18800 6322 18828 6666
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18788 6112 18840 6118
rect 18786 6080 18788 6089
rect 18840 6080 18842 6089
rect 18786 6015 18842 6024
rect 18892 5846 18920 8366
rect 18984 7546 19012 8588
rect 19076 8362 19104 8894
rect 19340 8910 19392 8916
rect 19246 8871 19302 8880
rect 19156 8832 19208 8838
rect 19156 8774 19208 8780
rect 19168 8514 19196 8774
rect 19260 8634 19288 8871
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19168 8486 19288 8514
rect 19064 8356 19116 8362
rect 19064 8298 19116 8304
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 18970 7168 19026 7177
rect 18970 7103 19026 7112
rect 18880 5840 18932 5846
rect 18880 5782 18932 5788
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18800 5098 18828 5646
rect 18984 5234 19012 7103
rect 19168 6798 19196 7890
rect 19260 7857 19288 8486
rect 19246 7848 19302 7857
rect 19246 7783 19302 7792
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 7410 19288 7686
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19168 6390 19196 6734
rect 19156 6384 19208 6390
rect 19156 6326 19208 6332
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18880 5160 18932 5166
rect 18880 5102 18932 5108
rect 18788 5092 18840 5098
rect 18788 5034 18840 5040
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18602 4448 18658 4457
rect 18602 4383 18658 4392
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18616 3398 18644 4082
rect 18708 3738 18736 4966
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18800 4214 18828 4422
rect 18788 4208 18840 4214
rect 18788 4150 18840 4156
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 3058 18644 3334
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18512 2508 18564 2514
rect 18512 2450 18564 2456
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 17328 1414 17448 1442
rect 17328 480 17356 1414
rect 17788 480 17816 2246
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 18524 1170 18552 2246
rect 18248 1142 18552 1170
rect 18248 480 18276 1142
rect 18708 480 18736 3062
rect 18800 1986 18828 3878
rect 18892 2582 18920 5102
rect 19064 4752 19116 4758
rect 19064 4694 19116 4700
rect 19076 4214 19104 4694
rect 19064 4208 19116 4214
rect 19116 4168 19196 4196
rect 19064 4150 19116 4156
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 18984 3738 19012 3878
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 18984 3398 19012 3538
rect 19168 3516 19196 4168
rect 19352 4078 19380 8910
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19444 8090 19472 8366
rect 19628 8090 19656 9687
rect 19800 9104 19852 9110
rect 19800 9046 19852 9052
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19444 7002 19472 7278
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19616 7200 19668 7206
rect 19616 7142 19668 7148
rect 19536 7002 19564 7142
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19628 6458 19656 7142
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19720 6322 19748 6598
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19536 5386 19564 6258
rect 19812 5710 19840 9046
rect 19904 7993 19932 10016
rect 20088 8922 20116 15535
rect 20180 14346 20208 17070
rect 20272 15706 20300 22063
rect 20626 21584 20682 21593
rect 20626 21519 20682 21528
rect 20350 21176 20406 21185
rect 20350 21111 20406 21120
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20364 15162 20392 21111
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20548 18329 20576 19246
rect 20534 18320 20590 18329
rect 20534 18255 20590 18264
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20548 17814 20576 18158
rect 20536 17808 20588 17814
rect 20536 17750 20588 17756
rect 20442 17368 20498 17377
rect 20442 17303 20498 17312
rect 20456 16794 20484 17303
rect 20640 16810 20668 21519
rect 20718 19816 20774 19825
rect 20718 19751 20774 19760
rect 20732 19514 20760 19751
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20718 18864 20774 18873
rect 20718 18799 20774 18808
rect 20732 18426 20760 18799
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20810 18320 20866 18329
rect 20810 18255 20866 18264
rect 20718 17912 20774 17921
rect 20718 17847 20774 17856
rect 20732 17338 20760 17847
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20548 16782 20668 16810
rect 20548 16674 20576 16782
rect 20456 16646 20576 16674
rect 20628 16652 20680 16658
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20456 15042 20484 16646
rect 20628 16594 20680 16600
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20364 15014 20484 15042
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20168 14340 20220 14346
rect 20168 14282 20220 14288
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 20180 12753 20208 13330
rect 20272 13297 20300 14758
rect 20364 14618 20392 15014
rect 20444 14952 20496 14958
rect 20444 14894 20496 14900
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20352 14476 20404 14482
rect 20352 14418 20404 14424
rect 20364 13410 20392 14418
rect 20456 13938 20484 14894
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20364 13382 20484 13410
rect 20352 13320 20404 13326
rect 20258 13288 20314 13297
rect 20352 13262 20404 13268
rect 20258 13223 20314 13232
rect 20364 12986 20392 13262
rect 20352 12980 20404 12986
rect 20272 12940 20352 12968
rect 20166 12744 20222 12753
rect 20166 12679 20222 12688
rect 20272 11694 20300 12940
rect 20352 12922 20404 12928
rect 20456 12866 20484 13382
rect 20364 12838 20484 12866
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20364 11354 20392 12838
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20456 12345 20484 12718
rect 20442 12336 20498 12345
rect 20548 12322 20576 15982
rect 20640 12442 20668 16594
rect 20718 16552 20774 16561
rect 20718 16487 20774 16496
rect 20732 16250 20760 16487
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 20732 12850 20760 13942
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20548 12294 20668 12322
rect 20442 12271 20498 12280
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 20180 9178 20208 10406
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 19996 8894 20116 8922
rect 19996 8634 20024 8894
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19890 7984 19946 7993
rect 19890 7919 19946 7928
rect 19904 7342 19932 7919
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19904 6866 19932 7142
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 19536 5358 19840 5386
rect 19616 5296 19668 5302
rect 19616 5238 19668 5244
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19536 4690 19564 5102
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19352 3738 19380 3878
rect 19444 3777 19472 3878
rect 19430 3768 19486 3777
rect 19340 3732 19392 3738
rect 19430 3703 19486 3712
rect 19340 3674 19392 3680
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19248 3528 19300 3534
rect 19168 3488 19248 3516
rect 19248 3470 19300 3476
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19246 2952 19302 2961
rect 19352 2938 19380 2994
rect 19302 2910 19380 2938
rect 19246 2887 19302 2896
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 19168 2650 19196 2790
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 18800 1958 19196 1986
rect 19168 480 19196 1958
rect 5446 232 5502 241
rect 5446 167 5502 176
rect 5906 0 5962 480
rect 6366 0 6422 480
rect 6826 0 6882 480
rect 7286 0 7342 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8758 0 8814 480
rect 9218 0 9274 480
rect 9678 0 9734 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 11058 0 11114 480
rect 11610 0 11666 480
rect 12070 0 12126 480
rect 12530 0 12586 480
rect 12990 0 13046 480
rect 13450 0 13506 480
rect 13910 0 13966 480
rect 14462 0 14518 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15842 0 15898 480
rect 16302 0 16358 480
rect 16762 0 16818 480
rect 17314 0 17370 480
rect 17774 0 17830 480
rect 18234 0 18290 480
rect 18694 0 18750 480
rect 19154 0 19210 480
rect 19260 241 19288 2382
rect 19352 2378 19380 2910
rect 19444 2514 19472 3606
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19340 2372 19392 2378
rect 19340 2314 19392 2320
rect 19444 1057 19472 2450
rect 19430 1048 19486 1057
rect 19430 983 19486 992
rect 19628 480 19656 5238
rect 19812 1850 19840 5358
rect 19904 3670 19932 6190
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19996 4282 20024 4966
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19892 3664 19944 3670
rect 19892 3606 19944 3612
rect 20088 2514 20116 8774
rect 20272 7274 20300 11154
rect 20456 10962 20484 12106
rect 20548 11898 20576 12174
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20364 10934 20484 10962
rect 20364 9382 20392 10934
rect 20548 10826 20576 11834
rect 20640 11286 20668 12294
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20456 10798 20576 10826
rect 20626 10840 20682 10849
rect 20456 10606 20484 10798
rect 20626 10775 20682 10784
rect 20640 10674 20668 10775
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20548 9926 20576 10542
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20548 9518 20576 9862
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20352 9104 20404 9110
rect 20352 9046 20404 9052
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 20180 5914 20208 6802
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20272 6458 20300 6734
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20364 6118 20392 9046
rect 20456 8974 20484 9318
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20456 8430 20484 8910
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 20180 5250 20208 5714
rect 20180 5222 20300 5250
rect 20168 5092 20220 5098
rect 20168 5034 20220 5040
rect 20180 4826 20208 5034
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20272 3602 20300 5222
rect 20456 4078 20484 8230
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20548 6186 20576 7414
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20640 6322 20668 7346
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20548 4162 20576 6122
rect 20640 5710 20668 6258
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20640 5370 20668 5646
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20548 4134 20668 4162
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20536 4004 20588 4010
rect 20536 3946 20588 3952
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 20272 2961 20300 3538
rect 20364 3194 20392 3878
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20456 2990 20484 3878
rect 20444 2984 20496 2990
rect 20258 2952 20314 2961
rect 20444 2926 20496 2932
rect 20258 2887 20260 2896
rect 20312 2887 20314 2896
rect 20260 2858 20312 2864
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 20180 2009 20208 2790
rect 20548 2530 20576 3946
rect 20640 2854 20668 4134
rect 20732 2990 20760 12582
rect 20824 9897 20852 18255
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 20916 11354 20944 12038
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20810 9888 20866 9897
rect 20810 9823 20866 9832
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20916 6934 20944 7822
rect 20904 6928 20956 6934
rect 20904 6870 20956 6876
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20812 5636 20864 5642
rect 20812 5578 20864 5584
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20824 2553 20852 5578
rect 20810 2544 20866 2553
rect 20548 2502 20668 2530
rect 20166 2000 20222 2009
rect 20166 1935 20222 1944
rect 19812 1822 20208 1850
rect 20180 480 20208 1822
rect 20640 480 20668 2502
rect 20810 2479 20866 2488
rect 20916 1601 20944 6054
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 20902 1592 20958 1601
rect 20902 1527 20958 1536
rect 21100 480 21128 4422
rect 21548 4072 21600 4078
rect 21548 4014 21600 4020
rect 21560 480 21588 4014
rect 22008 2100 22060 2106
rect 22008 2042 22060 2048
rect 22020 480 22048 2042
rect 22480 480 22508 5510
rect 19246 232 19302 241
rect 19246 167 19302 176
rect 19614 0 19670 480
rect 20166 0 20222 480
rect 20626 0 20682 480
rect 21086 0 21142 480
rect 21546 0 21602 480
rect 22006 0 22062 480
rect 22466 0 22522 480
<< via2 >>
rect 3146 22480 3202 22536
rect 3054 21528 3110 21584
rect 2502 21120 2558 21176
rect 1950 19760 2006 19816
rect 1950 19216 2006 19272
rect 1950 18808 2006 18864
rect 1674 18264 1730 18320
rect 1950 17856 2006 17912
rect 1858 17312 1914 17368
rect 1950 16496 2006 16552
rect 1950 15952 2006 16008
rect 2778 20168 2834 20224
rect 2778 15544 2834 15600
rect 1582 14048 1638 14104
rect 1950 15036 1952 15056
rect 1952 15036 2004 15056
rect 2004 15036 2006 15056
rect 1950 15000 2006 15036
rect 2778 14592 2834 14648
rect 1674 13640 1730 13696
rect 1582 13232 1638 13288
rect 662 3984 718 4040
rect 17222 22480 17278 22536
rect 3606 22072 3662 22128
rect 3698 16904 3754 16960
rect 4066 20576 4122 20632
rect 2502 3440 2558 3496
rect 2870 2488 2926 2544
rect 3054 2760 3110 2816
rect 2962 584 3018 640
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 3974 13368 4030 13424
rect 4066 12708 4122 12744
rect 4066 12688 4068 12708
rect 4068 12688 4120 12708
rect 4120 12688 4122 12708
rect 3974 12280 4030 12336
rect 4066 11328 4122 11384
rect 4066 10784 4122 10840
rect 4066 10376 4122 10432
rect 3974 9968 4030 10024
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4802 11600 4858 11656
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 3882 9424 3938 9480
rect 4066 9424 4122 9480
rect 4066 9016 4122 9072
rect 3974 8472 4030 8528
rect 3974 8336 4030 8392
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4434 8336 4490 8392
rect 5354 12008 5410 12064
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 3974 7112 4030 7168
rect 4066 6160 4122 6216
rect 3698 5616 3754 5672
rect 4066 5752 4122 5808
rect 3882 5208 3938 5264
rect 3974 4800 4030 4856
rect 3790 4664 3846 4720
rect 3698 3848 3754 3904
rect 4066 4256 4122 4312
rect 3422 1944 3478 2000
rect 3330 1536 3386 1592
rect 3606 992 3662 1048
rect 4066 2932 4068 2952
rect 4068 2932 4120 2952
rect 4120 2932 4122 2952
rect 4066 2896 4122 2932
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4986 7656 5042 7712
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 5262 8880 5318 8936
rect 5262 7520 5318 7576
rect 5262 7384 5318 7440
rect 5814 11192 5870 11248
rect 5906 9560 5962 9616
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 5538 3304 5594 3360
rect 6090 9594 6146 9650
rect 6642 11736 6698 11792
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7102 11756 7158 11792
rect 7102 11736 7104 11756
rect 7104 11736 7156 11756
rect 7156 11736 7158 11756
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 5998 7248 6054 7304
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 8298 13404 8300 13424
rect 8300 13404 8352 13424
rect 8352 13404 8354 13424
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 8298 13368 8354 13404
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 8850 11736 8906 11792
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7194 5072 7250 5128
rect 6182 3576 6238 3632
rect 6366 3440 6422 3496
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7838 6704 7894 6760
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7010 2760 7066 2816
rect 10046 12180 10048 12200
rect 10048 12180 10100 12200
rect 10100 12180 10102 12200
rect 9218 12008 9274 12064
rect 10046 12144 10102 12180
rect 9402 11872 9458 11928
rect 9126 11228 9128 11248
rect 9128 11228 9180 11248
rect 9180 11228 9182 11248
rect 9126 11192 9182 11228
rect 9494 11056 9550 11112
rect 10598 12316 10600 12336
rect 10600 12316 10652 12336
rect 10652 12316 10654 12336
rect 10598 12280 10654 12316
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 10506 11736 10562 11792
rect 8574 8880 8630 8936
rect 8482 8336 8538 8392
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 8298 3440 8354 3496
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 9126 7656 9182 7712
rect 8850 4664 8906 4720
rect 10230 10512 10286 10568
rect 11150 11736 11206 11792
rect 10598 10648 10654 10704
rect 10322 7792 10378 7848
rect 10506 6160 10562 6216
rect 10598 5092 10654 5128
rect 10598 5072 10600 5092
rect 10600 5072 10652 5092
rect 10652 5072 10654 5092
rect 10598 4664 10654 4720
rect 10414 3984 10470 4040
rect 12806 13404 12808 13424
rect 12808 13404 12860 13424
rect 12860 13404 12862 13424
rect 12806 13368 12862 13404
rect 11610 11600 11666 11656
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 10874 8472 10930 8528
rect 10782 7112 10838 7168
rect 11058 7540 11114 7576
rect 11058 7520 11060 7540
rect 11060 7520 11112 7540
rect 11112 7520 11114 7540
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11518 7420 11520 7440
rect 11520 7420 11572 7440
rect 11572 7420 11574 7440
rect 11518 7384 11574 7420
rect 10782 5788 10784 5808
rect 10784 5788 10836 5808
rect 10836 5788 10838 5808
rect 10782 5752 10838 5788
rect 11426 6724 11482 6760
rect 11426 6704 11428 6724
rect 11428 6704 11480 6724
rect 11480 6704 11482 6724
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 10690 3304 10746 3360
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11518 4936 11574 4992
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11058 3032 11114 3088
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 12622 12180 12624 12200
rect 12624 12180 12676 12200
rect 12676 12180 12678 12200
rect 12622 12144 12678 12180
rect 12070 11192 12126 11248
rect 11978 9696 12034 9752
rect 11978 7928 12034 7984
rect 12162 8916 12164 8936
rect 12164 8916 12216 8936
rect 12216 8916 12218 8936
rect 12162 8880 12218 8916
rect 12254 7792 12310 7848
rect 11978 3576 12034 3632
rect 12990 11872 13046 11928
rect 12898 9868 12900 9888
rect 12900 9868 12952 9888
rect 12952 9868 12954 9888
rect 12898 9832 12954 9868
rect 12898 9016 12954 9072
rect 12622 7948 12678 7984
rect 12622 7928 12624 7948
rect 12624 7928 12676 7948
rect 12676 7928 12678 7948
rect 12530 6724 12586 6760
rect 12530 6704 12532 6724
rect 12532 6704 12584 6724
rect 12584 6704 12586 6724
rect 12898 7112 12954 7168
rect 13358 11892 13414 11928
rect 13358 11872 13360 11892
rect 13360 11872 13412 11892
rect 13412 11872 13414 11892
rect 13450 9424 13506 9480
rect 13910 8880 13966 8936
rect 13082 6704 13138 6760
rect 12622 4120 12678 4176
rect 12438 3576 12494 3632
rect 12346 2760 12402 2816
rect 13082 4528 13138 4584
rect 13082 3052 13138 3088
rect 13082 3032 13084 3052
rect 13084 3032 13136 3052
rect 13136 3032 13138 3052
rect 12806 2796 12808 2816
rect 12808 2796 12860 2816
rect 12860 2796 12862 2816
rect 12806 2760 12862 2796
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14830 12316 14832 12336
rect 14832 12316 14884 12336
rect 14884 12316 14886 12336
rect 14830 12280 14886 12316
rect 15014 12280 15070 12336
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14278 10512 14334 10568
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14370 7792 14426 7848
rect 14646 9036 14702 9072
rect 14646 9016 14648 9036
rect 14648 9016 14700 9036
rect 14700 9016 14702 9036
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 15474 9832 15530 9888
rect 15198 5208 15254 5264
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 15474 7792 15530 7848
rect 16302 13388 16358 13424
rect 16302 13368 16304 13388
rect 16304 13368 16356 13388
rect 16356 13368 16358 13388
rect 16302 11328 16358 11384
rect 16302 11228 16304 11248
rect 16304 11228 16356 11248
rect 16356 11228 16358 11248
rect 16302 11192 16358 11228
rect 16118 10920 16174 10976
rect 15474 5616 15530 5672
rect 15382 3440 15438 3496
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 16486 11056 16542 11112
rect 16578 10648 16634 10704
rect 16210 9696 16266 9752
rect 16210 9016 16266 9072
rect 16578 8356 16634 8392
rect 16578 8336 16580 8356
rect 16580 8336 16632 8356
rect 16632 8336 16634 8356
rect 17038 11872 17094 11928
rect 18694 20576 18750 20632
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 20258 22072 20314 22128
rect 19982 20168 20038 20224
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 17958 16904 18014 16960
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 17958 15036 17960 15056
rect 17960 15036 18012 15056
rect 18012 15036 18014 15056
rect 17958 15000 18014 15036
rect 19890 15952 19946 16008
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 17130 11736 17186 11792
rect 17038 10648 17094 10704
rect 16762 7248 16818 7304
rect 16854 4120 16910 4176
rect 17222 5788 17224 5808
rect 17224 5788 17276 5808
rect 17276 5788 17278 5808
rect 17222 5752 17278 5788
rect 18142 12280 18198 12336
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 17958 10376 18014 10432
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 17958 9460 17960 9480
rect 17960 9460 18012 9480
rect 18012 9460 18014 9480
rect 17958 9424 18014 9460
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18602 9968 18658 10024
rect 18418 8064 18474 8120
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 17774 6024 17830 6080
rect 17590 2896 17646 2952
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 17958 5752 18014 5808
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 17958 4664 18014 4720
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18418 3732 18474 3768
rect 18418 3712 18420 3732
rect 18420 3712 18472 3732
rect 18472 3712 18474 3732
rect 18234 3440 18290 3496
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 19246 14048 19302 14104
rect 19154 13676 19156 13696
rect 19156 13676 19208 13696
rect 19208 13676 19210 13696
rect 19154 13640 19210 13676
rect 18970 12144 19026 12200
rect 18970 9324 18972 9344
rect 18972 9324 19024 9344
rect 19024 9324 19026 9344
rect 18970 9288 19026 9324
rect 19430 12144 19486 12200
rect 19890 14612 19946 14648
rect 20166 19216 20222 19272
rect 20074 15544 20130 15600
rect 19890 14592 19892 14612
rect 19892 14592 19944 14612
rect 19944 14592 19946 14612
rect 19982 12144 20038 12200
rect 19614 9696 19670 9752
rect 18786 6060 18788 6080
rect 18788 6060 18840 6080
rect 18840 6060 18842 6080
rect 18786 6024 18842 6060
rect 19246 8880 19302 8936
rect 18970 7112 19026 7168
rect 19246 7792 19302 7848
rect 18602 4392 18658 4448
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 20626 21528 20682 21584
rect 20350 21120 20406 21176
rect 20534 18264 20590 18320
rect 20442 17312 20498 17368
rect 20718 19760 20774 19816
rect 20718 18808 20774 18864
rect 20810 18264 20866 18320
rect 20718 17856 20774 17912
rect 20258 13232 20314 13288
rect 20166 12688 20222 12744
rect 20442 12280 20498 12336
rect 20718 16496 20774 16552
rect 19890 7928 19946 7984
rect 19430 3712 19486 3768
rect 19246 2896 19302 2952
rect 5446 176 5502 232
rect 19430 992 19486 1048
rect 20626 10784 20682 10840
rect 20258 2916 20314 2952
rect 20258 2896 20260 2916
rect 20260 2896 20312 2916
rect 20312 2896 20314 2916
rect 20810 9832 20866 9888
rect 20166 1944 20222 2000
rect 20810 2488 20866 2544
rect 20902 1536 20958 1592
rect 19246 176 19302 232
<< metal3 >>
rect 0 22538 480 22568
rect 3141 22538 3207 22541
rect 0 22536 3207 22538
rect 0 22480 3146 22536
rect 3202 22480 3207 22536
rect 0 22478 3207 22480
rect 0 22448 480 22478
rect 3141 22475 3207 22478
rect 17217 22538 17283 22541
rect 22320 22538 22800 22568
rect 17217 22536 22800 22538
rect 17217 22480 17222 22536
rect 17278 22480 22800 22536
rect 17217 22478 22800 22480
rect 17217 22475 17283 22478
rect 22320 22448 22800 22478
rect 0 22130 480 22160
rect 3601 22130 3667 22133
rect 0 22128 3667 22130
rect 0 22072 3606 22128
rect 3662 22072 3667 22128
rect 0 22070 3667 22072
rect 0 22040 480 22070
rect 3601 22067 3667 22070
rect 20253 22130 20319 22133
rect 22320 22130 22800 22160
rect 20253 22128 22800 22130
rect 20253 22072 20258 22128
rect 20314 22072 22800 22128
rect 20253 22070 22800 22072
rect 20253 22067 20319 22070
rect 22320 22040 22800 22070
rect 0 21586 480 21616
rect 3049 21586 3115 21589
rect 0 21584 3115 21586
rect 0 21528 3054 21584
rect 3110 21528 3115 21584
rect 0 21526 3115 21528
rect 0 21496 480 21526
rect 3049 21523 3115 21526
rect 20621 21586 20687 21589
rect 22320 21586 22800 21616
rect 20621 21584 22800 21586
rect 20621 21528 20626 21584
rect 20682 21528 22800 21584
rect 20621 21526 22800 21528
rect 20621 21523 20687 21526
rect 22320 21496 22800 21526
rect 0 21178 480 21208
rect 2497 21178 2563 21181
rect 0 21176 2563 21178
rect 0 21120 2502 21176
rect 2558 21120 2563 21176
rect 0 21118 2563 21120
rect 0 21088 480 21118
rect 2497 21115 2563 21118
rect 20345 21178 20411 21181
rect 22320 21178 22800 21208
rect 20345 21176 22800 21178
rect 20345 21120 20350 21176
rect 20406 21120 22800 21176
rect 20345 21118 22800 21120
rect 20345 21115 20411 21118
rect 22320 21088 22800 21118
rect 0 20634 480 20664
rect 4061 20634 4127 20637
rect 0 20632 4127 20634
rect 0 20576 4066 20632
rect 4122 20576 4127 20632
rect 0 20574 4127 20576
rect 0 20544 480 20574
rect 4061 20571 4127 20574
rect 18689 20634 18755 20637
rect 22320 20634 22800 20664
rect 18689 20632 22800 20634
rect 18689 20576 18694 20632
rect 18750 20576 22800 20632
rect 18689 20574 22800 20576
rect 18689 20571 18755 20574
rect 22320 20544 22800 20574
rect 0 20226 480 20256
rect 2773 20226 2839 20229
rect 0 20224 2839 20226
rect 0 20168 2778 20224
rect 2834 20168 2839 20224
rect 0 20166 2839 20168
rect 0 20136 480 20166
rect 2773 20163 2839 20166
rect 19977 20226 20043 20229
rect 22320 20226 22800 20256
rect 19977 20224 22800 20226
rect 19977 20168 19982 20224
rect 20038 20168 22800 20224
rect 19977 20166 22800 20168
rect 19977 20163 20043 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 0 19818 480 19848
rect 1945 19818 2011 19821
rect 0 19816 2011 19818
rect 0 19760 1950 19816
rect 2006 19760 2011 19816
rect 0 19758 2011 19760
rect 0 19728 480 19758
rect 1945 19755 2011 19758
rect 20713 19818 20779 19821
rect 22320 19818 22800 19848
rect 20713 19816 22800 19818
rect 20713 19760 20718 19816
rect 20774 19760 22800 19816
rect 20713 19758 22800 19760
rect 20713 19755 20779 19758
rect 22320 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 1945 19274 2011 19277
rect 0 19272 2011 19274
rect 0 19216 1950 19272
rect 2006 19216 2011 19272
rect 0 19214 2011 19216
rect 0 19184 480 19214
rect 1945 19211 2011 19214
rect 20161 19274 20227 19277
rect 22320 19274 22800 19304
rect 20161 19272 22800 19274
rect 20161 19216 20166 19272
rect 20222 19216 22800 19272
rect 20161 19214 22800 19216
rect 20161 19211 20227 19214
rect 22320 19184 22800 19214
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 0 18866 480 18896
rect 1945 18866 2011 18869
rect 0 18864 2011 18866
rect 0 18808 1950 18864
rect 2006 18808 2011 18864
rect 0 18806 2011 18808
rect 0 18776 480 18806
rect 1945 18803 2011 18806
rect 20713 18866 20779 18869
rect 22320 18866 22800 18896
rect 20713 18864 22800 18866
rect 20713 18808 20718 18864
rect 20774 18808 22800 18864
rect 20713 18806 22800 18808
rect 20713 18803 20779 18806
rect 22320 18776 22800 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 480 18352
rect 1669 18322 1735 18325
rect 0 18320 1735 18322
rect 0 18264 1674 18320
rect 1730 18264 1735 18320
rect 0 18262 1735 18264
rect 0 18232 480 18262
rect 1669 18259 1735 18262
rect 19926 18260 19932 18324
rect 19996 18322 20002 18324
rect 20529 18322 20595 18325
rect 19996 18320 20595 18322
rect 19996 18264 20534 18320
rect 20590 18264 20595 18320
rect 19996 18262 20595 18264
rect 19996 18260 20002 18262
rect 20529 18259 20595 18262
rect 20805 18322 20871 18325
rect 22320 18322 22800 18352
rect 20805 18320 22800 18322
rect 20805 18264 20810 18320
rect 20866 18264 22800 18320
rect 20805 18262 22800 18264
rect 20805 18259 20871 18262
rect 22320 18232 22800 18262
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 1945 17914 2011 17917
rect 0 17912 2011 17914
rect 0 17856 1950 17912
rect 2006 17856 2011 17912
rect 0 17854 2011 17856
rect 0 17824 480 17854
rect 1945 17851 2011 17854
rect 20713 17914 20779 17917
rect 22320 17914 22800 17944
rect 20713 17912 22800 17914
rect 20713 17856 20718 17912
rect 20774 17856 22800 17912
rect 20713 17854 22800 17856
rect 20713 17851 20779 17854
rect 22320 17824 22800 17854
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1853 17370 1919 17373
rect 0 17368 1919 17370
rect 0 17312 1858 17368
rect 1914 17312 1919 17368
rect 0 17310 1919 17312
rect 0 17280 480 17310
rect 1853 17307 1919 17310
rect 20437 17370 20503 17373
rect 22320 17370 22800 17400
rect 20437 17368 22800 17370
rect 20437 17312 20442 17368
rect 20498 17312 22800 17368
rect 20437 17310 22800 17312
rect 20437 17307 20503 17310
rect 22320 17280 22800 17310
rect 0 16962 480 16992
rect 3693 16962 3759 16965
rect 0 16960 3759 16962
rect 0 16904 3698 16960
rect 3754 16904 3759 16960
rect 0 16902 3759 16904
rect 0 16872 480 16902
rect 3693 16899 3759 16902
rect 17953 16962 18019 16965
rect 22320 16962 22800 16992
rect 17953 16960 22800 16962
rect 17953 16904 17958 16960
rect 18014 16904 22800 16960
rect 17953 16902 22800 16904
rect 17953 16899 18019 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 22320 16872 22800 16902
rect 14672 16831 14992 16832
rect 0 16554 480 16584
rect 1945 16554 2011 16557
rect 0 16552 2011 16554
rect 0 16496 1950 16552
rect 2006 16496 2011 16552
rect 0 16494 2011 16496
rect 0 16464 480 16494
rect 1945 16491 2011 16494
rect 20713 16554 20779 16557
rect 22320 16554 22800 16584
rect 20713 16552 22800 16554
rect 20713 16496 20718 16552
rect 20774 16496 22800 16552
rect 20713 16494 22800 16496
rect 20713 16491 20779 16494
rect 22320 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 16010 480 16040
rect 1945 16010 2011 16013
rect 0 16008 2011 16010
rect 0 15952 1950 16008
rect 2006 15952 2011 16008
rect 0 15950 2011 15952
rect 0 15920 480 15950
rect 1945 15947 2011 15950
rect 19885 16010 19951 16013
rect 22320 16010 22800 16040
rect 19885 16008 22800 16010
rect 19885 15952 19890 16008
rect 19946 15952 22800 16008
rect 19885 15950 22800 15952
rect 19885 15947 19951 15950
rect 22320 15920 22800 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 480 15632
rect 2773 15602 2839 15605
rect 0 15600 2839 15602
rect 0 15544 2778 15600
rect 2834 15544 2839 15600
rect 0 15542 2839 15544
rect 0 15512 480 15542
rect 2773 15539 2839 15542
rect 20069 15602 20135 15605
rect 22320 15602 22800 15632
rect 20069 15600 22800 15602
rect 20069 15544 20074 15600
rect 20130 15544 22800 15600
rect 20069 15542 22800 15544
rect 20069 15539 20135 15542
rect 22320 15512 22800 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 480 15088
rect 1945 15058 2011 15061
rect 0 15056 2011 15058
rect 0 15000 1950 15056
rect 2006 15000 2011 15056
rect 0 14998 2011 15000
rect 0 14968 480 14998
rect 1945 14995 2011 14998
rect 17953 15058 18019 15061
rect 22320 15058 22800 15088
rect 17953 15056 22800 15058
rect 17953 15000 17958 15056
rect 18014 15000 22800 15056
rect 17953 14998 22800 15000
rect 17953 14995 18019 14998
rect 22320 14968 22800 14998
rect 7808 14720 8128 14721
rect 0 14650 480 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 2773 14650 2839 14653
rect 0 14648 2839 14650
rect 0 14592 2778 14648
rect 2834 14592 2839 14648
rect 0 14590 2839 14592
rect 0 14560 480 14590
rect 2773 14587 2839 14590
rect 19885 14650 19951 14653
rect 22320 14650 22800 14680
rect 19885 14648 22800 14650
rect 19885 14592 19890 14648
rect 19946 14592 22800 14648
rect 19885 14590 22800 14592
rect 19885 14587 19951 14590
rect 22320 14560 22800 14590
rect 4376 14176 4696 14177
rect 0 14106 480 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1577 14106 1643 14109
rect 0 14104 1643 14106
rect 0 14048 1582 14104
rect 1638 14048 1643 14104
rect 0 14046 1643 14048
rect 0 14016 480 14046
rect 1577 14043 1643 14046
rect 19241 14106 19307 14109
rect 22320 14106 22800 14136
rect 19241 14104 22800 14106
rect 19241 14048 19246 14104
rect 19302 14048 22800 14104
rect 19241 14046 22800 14048
rect 19241 14043 19307 14046
rect 22320 14016 22800 14046
rect 0 13698 480 13728
rect 1669 13698 1735 13701
rect 0 13696 1735 13698
rect 0 13640 1674 13696
rect 1730 13640 1735 13696
rect 0 13638 1735 13640
rect 0 13608 480 13638
rect 1669 13635 1735 13638
rect 19149 13698 19215 13701
rect 22320 13698 22800 13728
rect 19149 13696 22800 13698
rect 19149 13640 19154 13696
rect 19210 13640 22800 13696
rect 19149 13638 22800 13640
rect 19149 13635 19215 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22320 13608 22800 13638
rect 14672 13567 14992 13568
rect 3969 13426 4035 13429
rect 8293 13426 8359 13429
rect 3969 13424 8359 13426
rect 3969 13368 3974 13424
rect 4030 13368 8298 13424
rect 8354 13368 8359 13424
rect 3969 13366 8359 13368
rect 3969 13363 4035 13366
rect 8293 13363 8359 13366
rect 12801 13426 12867 13429
rect 16297 13426 16363 13429
rect 12801 13424 16363 13426
rect 12801 13368 12806 13424
rect 12862 13368 16302 13424
rect 16358 13368 16363 13424
rect 12801 13366 16363 13368
rect 12801 13363 12867 13366
rect 16297 13363 16363 13366
rect 0 13290 480 13320
rect 1577 13290 1643 13293
rect 0 13288 1643 13290
rect 0 13232 1582 13288
rect 1638 13232 1643 13288
rect 0 13230 1643 13232
rect 0 13200 480 13230
rect 1577 13227 1643 13230
rect 20253 13290 20319 13293
rect 22320 13290 22800 13320
rect 20253 13288 22800 13290
rect 20253 13232 20258 13288
rect 20314 13232 22800 13288
rect 20253 13230 22800 13232
rect 20253 13227 20319 13230
rect 22320 13200 22800 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 0 12746 480 12776
rect 4061 12746 4127 12749
rect 0 12744 4127 12746
rect 0 12688 4066 12744
rect 4122 12688 4127 12744
rect 0 12686 4127 12688
rect 0 12656 480 12686
rect 4061 12683 4127 12686
rect 20161 12746 20227 12749
rect 22320 12746 22800 12776
rect 20161 12744 22800 12746
rect 20161 12688 20166 12744
rect 20222 12688 22800 12744
rect 20161 12686 22800 12688
rect 20161 12683 20227 12686
rect 22320 12656 22800 12686
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 480 12368
rect 3969 12338 4035 12341
rect 0 12336 4035 12338
rect 0 12280 3974 12336
rect 4030 12280 4035 12336
rect 0 12278 4035 12280
rect 0 12248 480 12278
rect 3969 12275 4035 12278
rect 10593 12338 10659 12341
rect 14825 12338 14891 12341
rect 10593 12336 14891 12338
rect 10593 12280 10598 12336
rect 10654 12280 14830 12336
rect 14886 12280 14891 12336
rect 10593 12278 14891 12280
rect 10593 12275 10659 12278
rect 14825 12275 14891 12278
rect 15009 12338 15075 12341
rect 18137 12338 18203 12341
rect 15009 12336 18203 12338
rect 15009 12280 15014 12336
rect 15070 12280 18142 12336
rect 18198 12280 18203 12336
rect 15009 12278 18203 12280
rect 15009 12275 15075 12278
rect 18137 12275 18203 12278
rect 20437 12338 20503 12341
rect 22320 12338 22800 12368
rect 20437 12336 22800 12338
rect 20437 12280 20442 12336
rect 20498 12280 22800 12336
rect 20437 12278 22800 12280
rect 20437 12275 20503 12278
rect 22320 12248 22800 12278
rect 10041 12202 10107 12205
rect 12617 12202 12683 12205
rect 18965 12202 19031 12205
rect 10041 12200 19031 12202
rect 10041 12144 10046 12200
rect 10102 12144 12622 12200
rect 12678 12144 18970 12200
rect 19026 12144 19031 12200
rect 10041 12142 19031 12144
rect 10041 12139 10107 12142
rect 12617 12139 12683 12142
rect 18965 12139 19031 12142
rect 19425 12202 19491 12205
rect 19977 12202 20043 12205
rect 19425 12200 20043 12202
rect 19425 12144 19430 12200
rect 19486 12144 19982 12200
rect 20038 12144 20043 12200
rect 19425 12142 20043 12144
rect 19425 12139 19491 12142
rect 19977 12139 20043 12142
rect 5349 12066 5415 12069
rect 9213 12066 9279 12069
rect 5349 12064 9279 12066
rect 5349 12008 5354 12064
rect 5410 12008 9218 12064
rect 9274 12008 9279 12064
rect 5349 12006 9279 12008
rect 5349 12003 5415 12006
rect 9213 12003 9279 12006
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 9397 11930 9463 11933
rect 4846 11928 9463 11930
rect 4846 11872 9402 11928
rect 9458 11872 9463 11928
rect 4846 11870 9463 11872
rect 0 11794 480 11824
rect 4846 11794 4906 11870
rect 9397 11867 9463 11870
rect 12985 11930 13051 11933
rect 13353 11930 13419 11933
rect 17033 11930 17099 11933
rect 12985 11928 13419 11930
rect 12985 11872 12990 11928
rect 13046 11872 13358 11928
rect 13414 11872 13419 11928
rect 12985 11870 13419 11872
rect 12985 11867 13051 11870
rect 13353 11867 13419 11870
rect 13494 11928 17099 11930
rect 13494 11872 17038 11928
rect 17094 11872 17099 11928
rect 13494 11870 17099 11872
rect 0 11734 4906 11794
rect 6637 11794 6703 11797
rect 7097 11794 7163 11797
rect 8845 11794 8911 11797
rect 6637 11792 8911 11794
rect 6637 11736 6642 11792
rect 6698 11736 7102 11792
rect 7158 11736 8850 11792
rect 8906 11736 8911 11792
rect 6637 11734 8911 11736
rect 0 11704 480 11734
rect 6637 11731 6703 11734
rect 7097 11731 7163 11734
rect 8845 11731 8911 11734
rect 10501 11794 10567 11797
rect 11145 11794 11211 11797
rect 13494 11794 13554 11870
rect 17033 11867 17099 11870
rect 10501 11792 13554 11794
rect 10501 11736 10506 11792
rect 10562 11736 11150 11792
rect 11206 11736 13554 11792
rect 10501 11734 13554 11736
rect 17125 11794 17191 11797
rect 22320 11794 22800 11824
rect 17125 11792 22800 11794
rect 17125 11736 17130 11792
rect 17186 11736 22800 11792
rect 17125 11734 22800 11736
rect 10501 11731 10567 11734
rect 11145 11731 11211 11734
rect 17125 11731 17191 11734
rect 22320 11704 22800 11734
rect 4797 11658 4863 11661
rect 11605 11658 11671 11661
rect 4797 11656 11671 11658
rect 4797 11600 4802 11656
rect 4858 11600 11610 11656
rect 11666 11600 11671 11656
rect 4797 11598 11671 11600
rect 4797 11595 4863 11598
rect 11605 11595 11671 11598
rect 7808 11456 8128 11457
rect 0 11386 480 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 4061 11386 4127 11389
rect 0 11384 4127 11386
rect 0 11328 4066 11384
rect 4122 11328 4127 11384
rect 0 11326 4127 11328
rect 0 11296 480 11326
rect 4061 11323 4127 11326
rect 16297 11386 16363 11389
rect 22320 11386 22800 11416
rect 16297 11384 22800 11386
rect 16297 11328 16302 11384
rect 16358 11328 22800 11384
rect 16297 11326 22800 11328
rect 16297 11323 16363 11326
rect 22320 11296 22800 11326
rect 5809 11250 5875 11253
rect 9121 11250 9187 11253
rect 5809 11248 9187 11250
rect 5809 11192 5814 11248
rect 5870 11192 9126 11248
rect 9182 11192 9187 11248
rect 5809 11190 9187 11192
rect 5809 11187 5875 11190
rect 9121 11187 9187 11190
rect 12065 11250 12131 11253
rect 16297 11250 16363 11253
rect 12065 11248 16363 11250
rect 12065 11192 12070 11248
rect 12126 11192 16302 11248
rect 16358 11192 16363 11248
rect 12065 11190 16363 11192
rect 12065 11187 12131 11190
rect 16297 11187 16363 11190
rect 9489 11114 9555 11117
rect 16481 11114 16547 11117
rect 9489 11112 16547 11114
rect 9489 11056 9494 11112
rect 9550 11056 16486 11112
rect 16542 11056 16547 11112
rect 9489 11054 16547 11056
rect 9489 11051 9555 11054
rect 16070 10981 16130 11054
rect 16481 11051 16547 11054
rect 16070 10976 16179 10981
rect 16070 10920 16118 10976
rect 16174 10920 16179 10976
rect 16070 10918 16179 10920
rect 16113 10915 16179 10918
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 4061 10842 4127 10845
rect 0 10840 4127 10842
rect 0 10784 4066 10840
rect 4122 10784 4127 10840
rect 0 10782 4127 10784
rect 0 10752 480 10782
rect 4061 10779 4127 10782
rect 20621 10842 20687 10845
rect 22320 10842 22800 10872
rect 20621 10840 22800 10842
rect 20621 10784 20626 10840
rect 20682 10784 22800 10840
rect 20621 10782 22800 10784
rect 20621 10779 20687 10782
rect 22320 10752 22800 10782
rect 10593 10706 10659 10709
rect 16573 10706 16639 10709
rect 17033 10706 17099 10709
rect 10593 10704 17099 10706
rect 10593 10648 10598 10704
rect 10654 10648 16578 10704
rect 16634 10648 17038 10704
rect 17094 10648 17099 10704
rect 10593 10646 17099 10648
rect 10593 10643 10659 10646
rect 16573 10643 16639 10646
rect 17033 10643 17099 10646
rect 10225 10570 10291 10573
rect 14273 10570 14339 10573
rect 19926 10570 19932 10572
rect 10225 10568 19932 10570
rect 10225 10512 10230 10568
rect 10286 10512 14278 10568
rect 14334 10512 19932 10568
rect 10225 10510 19932 10512
rect 10225 10507 10291 10510
rect 14273 10507 14339 10510
rect 19926 10508 19932 10510
rect 19996 10508 20002 10572
rect 0 10434 480 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 480 10374
rect 4061 10371 4127 10374
rect 17953 10434 18019 10437
rect 22320 10434 22800 10464
rect 17953 10432 22800 10434
rect 17953 10376 17958 10432
rect 18014 10376 22800 10432
rect 17953 10374 22800 10376
rect 17953 10371 18019 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22320 10344 22800 10374
rect 14672 10303 14992 10304
rect 0 10026 480 10056
rect 3969 10026 4035 10029
rect 0 10024 4035 10026
rect 0 9968 3974 10024
rect 4030 9968 4035 10024
rect 0 9966 4035 9968
rect 0 9936 480 9966
rect 3969 9963 4035 9966
rect 18597 10026 18663 10029
rect 22320 10026 22800 10056
rect 18597 10024 22800 10026
rect 18597 9968 18602 10024
rect 18658 9968 22800 10024
rect 18597 9966 22800 9968
rect 18597 9963 18663 9966
rect 22320 9936 22800 9966
rect 12893 9890 12959 9893
rect 15469 9890 15535 9893
rect 20805 9890 20871 9893
rect 12893 9888 15535 9890
rect 12893 9832 12898 9888
rect 12954 9832 15474 9888
rect 15530 9832 15535 9888
rect 12893 9830 15535 9832
rect 12893 9827 12959 9830
rect 15469 9827 15535 9830
rect 19566 9888 20871 9890
rect 19566 9832 20810 9888
rect 20866 9832 20871 9888
rect 19566 9830 20871 9832
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 19566 9757 19626 9830
rect 20805 9827 20871 9830
rect 11973 9754 12039 9757
rect 16205 9754 16271 9757
rect 11973 9752 16271 9754
rect 11973 9696 11978 9752
rect 12034 9696 16210 9752
rect 16266 9696 16271 9752
rect 11973 9694 16271 9696
rect 19566 9752 19675 9757
rect 19566 9696 19614 9752
rect 19670 9696 19675 9752
rect 19566 9694 19675 9696
rect 11973 9691 12039 9694
rect 16205 9691 16271 9694
rect 19609 9691 19675 9694
rect 6085 9652 6151 9655
rect 5950 9650 6151 9652
rect 5950 9621 6090 9650
rect 5901 9616 6090 9621
rect 5901 9560 5906 9616
rect 5962 9594 6090 9616
rect 6146 9594 6151 9650
rect 5962 9592 6151 9594
rect 5962 9560 6010 9592
rect 6085 9589 6151 9592
rect 5901 9558 6010 9560
rect 5901 9555 5967 9558
rect 0 9482 480 9512
rect 3877 9482 3943 9485
rect 0 9480 3943 9482
rect 0 9424 3882 9480
rect 3938 9424 3943 9480
rect 0 9422 3943 9424
rect 0 9392 480 9422
rect 3877 9419 3943 9422
rect 4061 9484 4127 9485
rect 4061 9480 4108 9484
rect 4172 9482 4178 9484
rect 13445 9482 13511 9485
rect 17953 9482 18019 9485
rect 22320 9482 22800 9512
rect 4061 9424 4066 9480
rect 4061 9420 4108 9424
rect 4172 9422 4218 9482
rect 13445 9480 15210 9482
rect 13445 9424 13450 9480
rect 13506 9424 15210 9480
rect 13445 9422 15210 9424
rect 4172 9420 4178 9422
rect 4061 9419 4127 9420
rect 13445 9419 13511 9422
rect 15150 9346 15210 9422
rect 17953 9480 22800 9482
rect 17953 9424 17958 9480
rect 18014 9424 22800 9480
rect 17953 9422 22800 9424
rect 17953 9419 18019 9422
rect 22320 9392 22800 9422
rect 18965 9346 19031 9349
rect 15150 9344 19031 9346
rect 15150 9288 18970 9344
rect 19026 9288 19031 9344
rect 15150 9286 19031 9288
rect 18965 9283 19031 9286
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9074 480 9104
rect 4061 9074 4127 9077
rect 0 9072 4127 9074
rect 0 9016 4066 9072
rect 4122 9016 4127 9072
rect 0 9014 4127 9016
rect 0 8984 480 9014
rect 4061 9011 4127 9014
rect 12893 9074 12959 9077
rect 14641 9074 14707 9077
rect 12893 9072 14707 9074
rect 12893 9016 12898 9072
rect 12954 9016 14646 9072
rect 14702 9016 14707 9072
rect 12893 9014 14707 9016
rect 12893 9011 12959 9014
rect 14641 9011 14707 9014
rect 16205 9074 16271 9077
rect 22320 9074 22800 9104
rect 16205 9072 22800 9074
rect 16205 9016 16210 9072
rect 16266 9016 22800 9072
rect 16205 9014 22800 9016
rect 16205 9011 16271 9014
rect 22320 8984 22800 9014
rect 5257 8938 5323 8941
rect 8569 8938 8635 8941
rect 5257 8936 8635 8938
rect 5257 8880 5262 8936
rect 5318 8880 8574 8936
rect 8630 8880 8635 8936
rect 5257 8878 8635 8880
rect 5257 8875 5323 8878
rect 8569 8875 8635 8878
rect 12157 8938 12223 8941
rect 13905 8938 13971 8941
rect 19241 8938 19307 8941
rect 12157 8936 13971 8938
rect 12157 8880 12162 8936
rect 12218 8880 13910 8936
rect 13966 8880 13971 8936
rect 12157 8878 13971 8880
rect 12157 8875 12223 8878
rect 13905 8875 13971 8878
rect 17726 8936 19307 8938
rect 17726 8880 19246 8936
rect 19302 8880 19307 8936
rect 17726 8878 19307 8880
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 0 8530 480 8560
rect 3969 8530 4035 8533
rect 0 8528 4035 8530
rect 0 8472 3974 8528
rect 4030 8472 4035 8528
rect 0 8470 4035 8472
rect 0 8440 480 8470
rect 3969 8467 4035 8470
rect 10869 8530 10935 8533
rect 17726 8530 17786 8878
rect 19241 8875 19307 8878
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 22320 8530 22800 8560
rect 10869 8528 17786 8530
rect 10869 8472 10874 8528
rect 10930 8472 17786 8528
rect 10869 8470 17786 8472
rect 18094 8470 22800 8530
rect 10869 8467 10935 8470
rect 3969 8394 4035 8397
rect 4102 8394 4108 8396
rect 3969 8392 4108 8394
rect 3969 8336 3974 8392
rect 4030 8336 4108 8392
rect 3969 8334 4108 8336
rect 3969 8331 4035 8334
rect 4102 8332 4108 8334
rect 4172 8332 4178 8396
rect 4429 8394 4495 8397
rect 8477 8394 8543 8397
rect 4429 8392 8543 8394
rect 4429 8336 4434 8392
rect 4490 8336 8482 8392
rect 8538 8336 8543 8392
rect 4429 8334 8543 8336
rect 4429 8331 4495 8334
rect 8477 8331 8543 8334
rect 16573 8394 16639 8397
rect 18094 8394 18154 8470
rect 22320 8440 22800 8470
rect 16573 8392 18154 8394
rect 16573 8336 16578 8392
rect 16634 8336 18154 8392
rect 16573 8334 18154 8336
rect 16573 8331 16639 8334
rect 7808 8192 8128 8193
rect 0 8122 480 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 18413 8122 18479 8125
rect 22320 8122 22800 8152
rect 0 8062 4906 8122
rect 0 8032 480 8062
rect 4846 7986 4906 8062
rect 18413 8120 22800 8122
rect 18413 8064 18418 8120
rect 18474 8064 22800 8120
rect 18413 8062 22800 8064
rect 18413 8059 18479 8062
rect 22320 8032 22800 8062
rect 11973 7986 12039 7989
rect 4846 7984 12039 7986
rect 4846 7928 11978 7984
rect 12034 7928 12039 7984
rect 4846 7926 12039 7928
rect 11973 7923 12039 7926
rect 12617 7986 12683 7989
rect 19885 7986 19951 7989
rect 12617 7984 19951 7986
rect 12617 7928 12622 7984
rect 12678 7928 19890 7984
rect 19946 7928 19951 7984
rect 12617 7926 19951 7928
rect 12617 7923 12683 7926
rect 19885 7923 19951 7926
rect 10317 7850 10383 7853
rect 4110 7848 10383 7850
rect 4110 7792 10322 7848
rect 10378 7792 10383 7848
rect 4110 7790 10383 7792
rect 0 7578 480 7608
rect 4110 7578 4170 7790
rect 10317 7787 10383 7790
rect 12249 7850 12315 7853
rect 14365 7850 14431 7853
rect 15469 7850 15535 7853
rect 12249 7848 15535 7850
rect 12249 7792 12254 7848
rect 12310 7792 14370 7848
rect 14426 7792 15474 7848
rect 15530 7792 15535 7848
rect 12249 7790 15535 7792
rect 12249 7787 12315 7790
rect 14365 7787 14431 7790
rect 15469 7787 15535 7790
rect 19241 7850 19307 7853
rect 19241 7848 19442 7850
rect 19241 7792 19246 7848
rect 19302 7792 19442 7848
rect 19241 7790 19442 7792
rect 19241 7787 19307 7790
rect 4981 7714 5047 7717
rect 9121 7714 9187 7717
rect 4981 7712 9187 7714
rect 4981 7656 4986 7712
rect 5042 7656 9126 7712
rect 9182 7656 9187 7712
rect 4981 7654 9187 7656
rect 4981 7651 5047 7654
rect 9121 7651 9187 7654
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 0 7518 4170 7578
rect 5257 7578 5323 7581
rect 11053 7578 11119 7581
rect 5257 7576 11119 7578
rect 5257 7520 5262 7576
rect 5318 7520 11058 7576
rect 11114 7520 11119 7576
rect 5257 7518 11119 7520
rect 19382 7578 19442 7790
rect 22320 7578 22800 7608
rect 19382 7518 22800 7578
rect 0 7488 480 7518
rect 5257 7515 5323 7518
rect 11053 7515 11119 7518
rect 22320 7488 22800 7518
rect 5257 7442 5323 7445
rect 11513 7442 11579 7445
rect 5257 7440 11579 7442
rect 5257 7384 5262 7440
rect 5318 7384 11518 7440
rect 11574 7384 11579 7440
rect 5257 7382 11579 7384
rect 5257 7379 5323 7382
rect 11513 7379 11579 7382
rect 5993 7306 6059 7309
rect 16757 7306 16823 7309
rect 5993 7304 16823 7306
rect 5993 7248 5998 7304
rect 6054 7248 16762 7304
rect 16818 7248 16823 7304
rect 5993 7246 16823 7248
rect 5993 7243 6059 7246
rect 16757 7243 16823 7246
rect 0 7170 480 7200
rect 3969 7170 4035 7173
rect 0 7168 4035 7170
rect 0 7112 3974 7168
rect 4030 7112 4035 7168
rect 0 7110 4035 7112
rect 0 7080 480 7110
rect 3969 7107 4035 7110
rect 10777 7170 10843 7173
rect 12893 7170 12959 7173
rect 10777 7168 12959 7170
rect 10777 7112 10782 7168
rect 10838 7112 12898 7168
rect 12954 7112 12959 7168
rect 10777 7110 12959 7112
rect 10777 7107 10843 7110
rect 12893 7107 12959 7110
rect 18965 7170 19031 7173
rect 22320 7170 22800 7200
rect 18965 7168 22800 7170
rect 18965 7112 18970 7168
rect 19026 7112 22800 7168
rect 18965 7110 22800 7112
rect 18965 7107 19031 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 22320 7080 22800 7110
rect 14672 7039 14992 7040
rect 0 6762 480 6792
rect 7833 6762 7899 6765
rect 0 6760 7899 6762
rect 0 6704 7838 6760
rect 7894 6704 7899 6760
rect 0 6702 7899 6704
rect 0 6672 480 6702
rect 7833 6699 7899 6702
rect 11421 6762 11487 6765
rect 12525 6762 12591 6765
rect 11421 6760 12591 6762
rect 11421 6704 11426 6760
rect 11482 6704 12530 6760
rect 12586 6704 12591 6760
rect 11421 6702 12591 6704
rect 11421 6699 11487 6702
rect 12525 6699 12591 6702
rect 13077 6762 13143 6765
rect 22320 6762 22800 6792
rect 13077 6760 22800 6762
rect 13077 6704 13082 6760
rect 13138 6704 22800 6760
rect 13077 6702 22800 6704
rect 13077 6699 13143 6702
rect 22320 6672 22800 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 0 6218 480 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 480 6158
rect 4061 6155 4127 6158
rect 10501 6218 10567 6221
rect 22320 6218 22800 6248
rect 10501 6216 22800 6218
rect 10501 6160 10506 6216
rect 10562 6160 22800 6216
rect 10501 6158 22800 6160
rect 10501 6155 10567 6158
rect 22320 6128 22800 6158
rect 17769 6082 17835 6085
rect 18781 6084 18847 6085
rect 18781 6082 18828 6084
rect 17769 6080 18828 6082
rect 17769 6024 17774 6080
rect 17830 6024 18786 6080
rect 17769 6022 18828 6024
rect 17769 6019 17835 6022
rect 18781 6020 18828 6022
rect 18892 6020 18898 6084
rect 18781 6019 18847 6020
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 480 5750
rect 4061 5747 4127 5750
rect 10777 5810 10843 5813
rect 17217 5810 17283 5813
rect 10777 5808 17283 5810
rect 10777 5752 10782 5808
rect 10838 5752 17222 5808
rect 17278 5752 17283 5808
rect 10777 5750 17283 5752
rect 10777 5747 10843 5750
rect 17217 5747 17283 5750
rect 17953 5810 18019 5813
rect 22320 5810 22800 5840
rect 17953 5808 22800 5810
rect 17953 5752 17958 5808
rect 18014 5752 22800 5808
rect 17953 5750 22800 5752
rect 17953 5747 18019 5750
rect 22320 5720 22800 5750
rect 3693 5674 3759 5677
rect 15469 5674 15535 5677
rect 3693 5672 15535 5674
rect 3693 5616 3698 5672
rect 3754 5616 15474 5672
rect 15530 5616 15535 5672
rect 3693 5614 15535 5616
rect 3693 5611 3759 5614
rect 15469 5611 15535 5614
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 480 5296
rect 3877 5266 3943 5269
rect 15193 5266 15259 5269
rect 22320 5266 22800 5296
rect 0 5264 3943 5266
rect 0 5208 3882 5264
rect 3938 5208 3943 5264
rect 0 5206 3943 5208
rect 0 5176 480 5206
rect 3877 5203 3943 5206
rect 13862 5264 15259 5266
rect 13862 5208 15198 5264
rect 15254 5208 15259 5264
rect 13862 5206 15259 5208
rect 7189 5130 7255 5133
rect 10593 5130 10659 5133
rect 13862 5130 13922 5206
rect 15193 5203 15259 5206
rect 15334 5206 22800 5266
rect 15334 5130 15394 5206
rect 22320 5176 22800 5206
rect 7189 5128 13922 5130
rect 7189 5072 7194 5128
rect 7250 5072 10598 5128
rect 10654 5072 13922 5128
rect 7189 5070 13922 5072
rect 14414 5070 15394 5130
rect 7189 5067 7255 5070
rect 10593 5067 10659 5070
rect 11513 4994 11579 4997
rect 14414 4994 14474 5070
rect 11513 4992 14474 4994
rect 11513 4936 11518 4992
rect 11574 4936 14474 4992
rect 11513 4934 14474 4936
rect 11513 4931 11579 4934
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 3969 4858 4035 4861
rect 22320 4858 22800 4888
rect 0 4856 4035 4858
rect 0 4800 3974 4856
rect 4030 4800 4035 4856
rect 0 4798 4035 4800
rect 0 4768 480 4798
rect 3969 4795 4035 4798
rect 18094 4798 22800 4858
rect 3785 4722 3851 4725
rect 8845 4722 8911 4725
rect 3785 4720 8911 4722
rect 3785 4664 3790 4720
rect 3846 4664 8850 4720
rect 8906 4664 8911 4720
rect 3785 4662 8911 4664
rect 3785 4659 3851 4662
rect 8845 4659 8911 4662
rect 10593 4722 10659 4725
rect 17953 4722 18019 4725
rect 10593 4720 18019 4722
rect 10593 4664 10598 4720
rect 10654 4664 17958 4720
rect 18014 4664 18019 4720
rect 10593 4662 18019 4664
rect 10593 4659 10659 4662
rect 17953 4659 18019 4662
rect 13077 4586 13143 4589
rect 18094 4586 18154 4798
rect 22320 4768 22800 4798
rect 13077 4584 18154 4586
rect 13077 4528 13082 4584
rect 13138 4528 18154 4584
rect 13077 4526 18154 4528
rect 13077 4523 13143 4526
rect 18597 4448 18663 4453
rect 18597 4392 18602 4448
rect 18658 4392 18663 4448
rect 18597 4387 18663 4392
rect 4376 4384 4696 4385
rect 0 4314 480 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 4061 4314 4127 4317
rect 0 4312 4127 4314
rect 0 4256 4066 4312
rect 4122 4256 4127 4312
rect 0 4254 4127 4256
rect 18600 4314 18660 4387
rect 22320 4314 22800 4344
rect 18600 4254 22800 4314
rect 0 4224 480 4254
rect 4061 4251 4127 4254
rect 22320 4224 22800 4254
rect 12617 4178 12683 4181
rect 16849 4178 16915 4181
rect 12617 4176 16915 4178
rect 12617 4120 12622 4176
rect 12678 4120 16854 4176
rect 16910 4120 16915 4176
rect 12617 4118 16915 4120
rect 12617 4115 12683 4118
rect 16849 4115 16915 4118
rect 657 4042 723 4045
rect 10409 4042 10475 4045
rect 657 4040 10475 4042
rect 657 3984 662 4040
rect 718 3984 10414 4040
rect 10470 3984 10475 4040
rect 657 3982 10475 3984
rect 657 3979 723 3982
rect 10409 3979 10475 3982
rect 0 3906 480 3936
rect 3693 3906 3759 3909
rect 22320 3906 22800 3936
rect 0 3904 3759 3906
rect 0 3848 3698 3904
rect 3754 3848 3759 3904
rect 0 3846 3759 3848
rect 0 3816 480 3846
rect 3693 3843 3759 3846
rect 15150 3846 22800 3906
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 6177 3634 6243 3637
rect 11973 3634 12039 3637
rect 6177 3632 12039 3634
rect 6177 3576 6182 3632
rect 6238 3576 11978 3632
rect 12034 3576 12039 3632
rect 6177 3574 12039 3576
rect 6177 3571 6243 3574
rect 11973 3571 12039 3574
rect 12433 3634 12499 3637
rect 15150 3634 15210 3846
rect 22320 3816 22800 3846
rect 18413 3770 18479 3773
rect 19425 3770 19491 3773
rect 18413 3768 19491 3770
rect 18413 3712 18418 3768
rect 18474 3712 19430 3768
rect 19486 3712 19491 3768
rect 18413 3710 19491 3712
rect 18413 3707 18479 3710
rect 19425 3707 19491 3710
rect 12433 3632 15210 3634
rect 12433 3576 12438 3632
rect 12494 3576 15210 3632
rect 12433 3574 15210 3576
rect 12433 3571 12499 3574
rect 0 3498 480 3528
rect 2497 3498 2563 3501
rect 0 3496 2563 3498
rect 0 3440 2502 3496
rect 2558 3440 2563 3496
rect 0 3438 2563 3440
rect 0 3408 480 3438
rect 2497 3435 2563 3438
rect 6361 3498 6427 3501
rect 8293 3498 8359 3501
rect 15377 3498 15443 3501
rect 6361 3496 8359 3498
rect 6361 3440 6366 3496
rect 6422 3440 8298 3496
rect 8354 3440 8359 3496
rect 6361 3438 8359 3440
rect 6361 3435 6427 3438
rect 8293 3435 8359 3438
rect 11102 3496 15443 3498
rect 11102 3440 15382 3496
rect 15438 3440 15443 3496
rect 11102 3438 15443 3440
rect 5533 3362 5599 3365
rect 10685 3362 10751 3365
rect 11102 3362 11162 3438
rect 15377 3435 15443 3438
rect 18229 3498 18295 3501
rect 22320 3498 22800 3528
rect 18229 3496 22800 3498
rect 18229 3440 18234 3496
rect 18290 3440 22800 3496
rect 18229 3438 22800 3440
rect 18229 3435 18295 3438
rect 22320 3408 22800 3438
rect 5533 3360 11162 3362
rect 5533 3304 5538 3360
rect 5594 3304 10690 3360
rect 10746 3304 11162 3360
rect 5533 3302 11162 3304
rect 5533 3299 5599 3302
rect 10685 3299 10751 3302
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 11053 3090 11119 3093
rect 13077 3090 13143 3093
rect 11053 3088 13143 3090
rect 11053 3032 11058 3088
rect 11114 3032 13082 3088
rect 13138 3032 13143 3088
rect 11053 3030 13143 3032
rect 11053 3027 11119 3030
rect 13077 3027 13143 3030
rect 0 2954 480 2984
rect 4061 2954 4127 2957
rect 0 2952 4127 2954
rect 0 2896 4066 2952
rect 4122 2896 4127 2952
rect 0 2894 4127 2896
rect 0 2864 480 2894
rect 4061 2891 4127 2894
rect 17585 2954 17651 2957
rect 19241 2954 19307 2957
rect 17585 2952 19307 2954
rect 17585 2896 17590 2952
rect 17646 2896 19246 2952
rect 19302 2896 19307 2952
rect 17585 2894 19307 2896
rect 17585 2891 17651 2894
rect 19241 2891 19307 2894
rect 20253 2954 20319 2957
rect 22320 2954 22800 2984
rect 20253 2952 22800 2954
rect 20253 2896 20258 2952
rect 20314 2896 22800 2952
rect 20253 2894 22800 2896
rect 20253 2891 20319 2894
rect 22320 2864 22800 2894
rect 3049 2818 3115 2821
rect 7005 2818 7071 2821
rect 3049 2816 7071 2818
rect 3049 2760 3054 2816
rect 3110 2760 7010 2816
rect 7066 2760 7071 2816
rect 3049 2758 7071 2760
rect 3049 2755 3115 2758
rect 7005 2755 7071 2758
rect 12341 2818 12407 2821
rect 12801 2818 12867 2821
rect 12341 2816 12867 2818
rect 12341 2760 12346 2816
rect 12402 2760 12806 2816
rect 12862 2760 12867 2816
rect 12341 2758 12867 2760
rect 12341 2755 12407 2758
rect 12801 2755 12867 2758
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 480 2576
rect 2865 2546 2931 2549
rect 0 2544 2931 2546
rect 0 2488 2870 2544
rect 2926 2488 2931 2544
rect 0 2486 2931 2488
rect 0 2456 480 2486
rect 2865 2483 2931 2486
rect 20805 2546 20871 2549
rect 22320 2546 22800 2576
rect 20805 2544 22800 2546
rect 20805 2488 20810 2544
rect 20866 2488 22800 2544
rect 20805 2486 22800 2488
rect 20805 2483 20871 2486
rect 22320 2456 22800 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 480 2032
rect 3417 2002 3483 2005
rect 0 2000 3483 2002
rect 0 1944 3422 2000
rect 3478 1944 3483 2000
rect 0 1942 3483 1944
rect 0 1912 480 1942
rect 3417 1939 3483 1942
rect 20161 2002 20227 2005
rect 22320 2002 22800 2032
rect 20161 2000 22800 2002
rect 20161 1944 20166 2000
rect 20222 1944 22800 2000
rect 20161 1942 22800 1944
rect 20161 1939 20227 1942
rect 22320 1912 22800 1942
rect 0 1594 480 1624
rect 3325 1594 3391 1597
rect 0 1592 3391 1594
rect 0 1536 3330 1592
rect 3386 1536 3391 1592
rect 0 1534 3391 1536
rect 0 1504 480 1534
rect 3325 1531 3391 1534
rect 20897 1594 20963 1597
rect 22320 1594 22800 1624
rect 20897 1592 22800 1594
rect 20897 1536 20902 1592
rect 20958 1536 22800 1592
rect 20897 1534 22800 1536
rect 20897 1531 20963 1534
rect 22320 1504 22800 1534
rect 0 1050 480 1080
rect 3601 1050 3667 1053
rect 0 1048 3667 1050
rect 0 992 3606 1048
rect 3662 992 3667 1048
rect 0 990 3667 992
rect 0 960 480 990
rect 3601 987 3667 990
rect 19425 1050 19491 1053
rect 22320 1050 22800 1080
rect 19425 1048 22800 1050
rect 19425 992 19430 1048
rect 19486 992 22800 1048
rect 19425 990 22800 992
rect 19425 987 19491 990
rect 22320 960 22800 990
rect 0 642 480 672
rect 2957 642 3023 645
rect 0 640 3023 642
rect 0 584 2962 640
rect 3018 584 3023 640
rect 0 582 3023 584
rect 0 552 480 582
rect 2957 579 3023 582
rect 18822 580 18828 644
rect 18892 642 18898 644
rect 22320 642 22800 672
rect 18892 582 22800 642
rect 18892 580 18898 582
rect 22320 552 22800 582
rect 0 234 480 264
rect 5441 234 5507 237
rect 0 232 5507 234
rect 0 176 5446 232
rect 5502 176 5507 232
rect 0 174 5507 176
rect 0 144 480 174
rect 5441 171 5507 174
rect 19241 234 19307 237
rect 22320 234 22800 264
rect 19241 232 22800 234
rect 19241 176 19246 232
rect 19302 176 22800 232
rect 19241 174 22800 176
rect 19241 171 19307 174
rect 22320 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 19932 18260 19996 18324
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 19932 10508 19996 10572
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 4108 9480 4172 9484
rect 4108 9424 4122 9480
rect 4122 9424 4172 9480
rect 4108 9420 4172 9424
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 4108 8332 4172 8396
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 18828 6080 18892 6084
rect 18828 6024 18842 6080
rect 18842 6024 18892 6080
rect 18828 6020 18892 6024
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
rect 18828 580 18892 644
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4107 9484 4173 9485
rect 4107 9420 4108 9484
rect 4172 9420 4173 9484
rect 4107 9419 4173 9420
rect 4110 8397 4170 9419
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4107 8396 4173 8397
rect 4107 8332 4108 8396
rect 4172 8332 4173 8396
rect 4107 8331 4173 8332
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 19931 18324 19997 18325
rect 19931 18260 19932 18324
rect 19996 18260 19997 18324
rect 19931 18259 19997 18260
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 19934 10573 19994 18259
rect 19931 10572 19997 10573
rect 19931 10508 19932 10572
rect 19996 10508 19997 10572
rect 19931 10507 19997 10508
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18827 6084 18893 6085
rect 18827 6020 18828 6084
rect 18892 6020 18893 6084
rect 18827 6019 18893 6020
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
rect 18830 645 18890 6019
rect 18827 644 18893 645
rect 18827 580 18828 644
rect 18892 580 18893 644
rect 18827 579 18893 580
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2484 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2484 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _032_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3128 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1605641404
transform 1 0 4140 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23
timestamp 1605641404
transform 1 0 3220 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_21 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_31
timestamp 1605641404
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1605641404
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1605641404
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1605641404
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_42
timestamp 1605641404
transform 1 0 4968 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1605641404
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 8556 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 7728 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71
timestamp 1605641404
transform 1 0 7636 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1605641404
transform 1 0 8556 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_78
timestamp 1605641404
transform 1 0 8280 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10028 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 8832 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90
timestamp 1605641404
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1605641404
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_90
timestamp 1605641404
transform 1 0 9384 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_96
timestamp 1605641404
transform 1 0 9936 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1605641404
transform 1 0 11500 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_109
timestamp 1605641404
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11316 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _097_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10764 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1605641404
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1605641404
transform 1 0 11776 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1605641404
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13432 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13340 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14076 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1605641404
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_139
timestamp 1605641404
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1605641404
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_140
timestamp 1605641404
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1605641404
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_146
timestamp 1605641404
transform 1 0 14536 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1605641404
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1605641404
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14812 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1605641404
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1605641404
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_162
timestamp 1605641404
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 16100 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16192 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1605641404
transform 1 0 15548 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_170
timestamp 1605641404
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_172
timestamp 1605641404
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_176
timestamp 1605641404
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1605641404
transform 1 0 17112 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1605641404
transform 1 0 16928 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1605641404
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1605641404
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1605641404
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1605641404
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1605641404
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1605641404
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20148 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19044 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1605641404
transform 1 0 19688 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18676 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1605641404
transform 1 0 18676 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_204
timestamp 1605641404
transform 1 0 19872 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_188
timestamp 1605641404
transform 1 0 18400 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_200
timestamp 1605641404
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1605641404
transform 1 0 20700 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1605641404
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1605641404
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_211
timestamp 1605641404
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_217
timestamp 1605641404
transform 1 0 21068 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1605641404
transform 1 0 2576 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_15
timestamp 1605641404
transform 1 0 2484 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_25
timestamp 1605641404
transform 1 0 3404 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1605641404
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1605641404
transform 1 0 6348 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6808 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5060 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_52
timestamp 1605641404
transform 1 0 5888 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_56
timestamp 1605641404
transform 1 0 6256 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_60
timestamp 1605641404
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8464 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_78
timestamp 1605641404
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 10028 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1605641404
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11684 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_113
timestamp 1605641404
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_124
timestamp 1605641404
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1605641404
transform 1 0 13708 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1605641404
transform 1 0 12696 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14168 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_135
timestamp 1605641404
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_140
timestamp 1605641404
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1605641404
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 1605641404
transform 1 0 16100 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16468 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_2_183
timestamp 1605641404
transform 1 0 17940 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1605641404
transform 1 0 18584 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19596 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp 1605641404
transform 1 0 18492 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_199
timestamp 1605641404
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1605641404
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1605641404
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_218
timestamp 1605641404
transform 1 0 21160 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 2944 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1932 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_18
timestamp 1605641404
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4600 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_36
timestamp 1605641404
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 5612 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 1605641404
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1605641404
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7820 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1605641404
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10028 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_3_89
timestamp 1605641404
transform 1 0 9292 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1605641404
transform 1 0 11776 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1605641404
transform 1 0 11500 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1605641404
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13800 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_3_132
timestamp 1605641404
transform 1 0 13248 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15456 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_154
timestamp 1605641404
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1605641404
transform 1 0 16284 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1605641404
transform 1 0 16560 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_177
timestamp 1605641404
transform 1 0 17388 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1605641404
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1605641404
transform 1 0 18400 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1605641404
transform 1 0 18952 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 19964 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_192
timestamp 1605641404
transform 1 0 18768 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_203
timestamp 1605641404
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_214
timestamp 1605641404
transform 1 0 20792 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_19
timestamp 1605641404
transform 1 0 2852 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4508 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1605641404
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1605641404
transform 1 0 6532 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_53
timestamp 1605641404
transform 1 0 5980 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8096 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_68
timestamp 1605641404
transform 1 0 7360 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp 1605641404
transform 1 0 8924 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1605641404
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1605641404
transform 1 0 10488 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1605641404
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11408 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_110
timestamp 1605641404
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1605641404
transform 1 0 13064 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13524 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_128
timestamp 1605641404
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_133
timestamp 1605641404
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16100 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1605641404
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_158
timestamp 1605641404
transform 1 0 15640 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_162
timestamp 1605641404
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 17112 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_172
timestamp 1605641404
transform 1 0 16928 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 18768 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_190
timestamp 1605641404
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_208
timestamp 1605641404
transform 1 0 20240 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1605641404
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1605641404
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 1932 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 3680 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_5_25
timestamp 1605641404
transform 1 0 3404 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5336 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_44
timestamp 1605641404
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_55
timestamp 1605641404
transform 1 0 6164 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1605641404
transform 1 0 6992 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7544 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_5_67
timestamp 1605641404
transform 1 0 7268 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1605641404
transform 1 0 10120 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 9200 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_86
timestamp 1605641404
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_91
timestamp 1605641404
transform 1 0 9476 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_97
timestamp 1605641404
transform 1 0 10028 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1605641404
transform 1 0 11132 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_107
timestamp 1605641404
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1605641404
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13616 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1605641404
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_145
timestamp 1605641404
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1605641404
transform 1 0 16376 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14628 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_5_163
timestamp 1605641404
transform 1 0 16100 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1605641404
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1605641404
transform 1 0 16928 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_170
timestamp 1605641404
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1605641404
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 19596 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1605641404
transform 1 0 18584 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1605641404
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_199
timestamp 1605641404
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_217
timestamp 1605641404
transform 1 0 21068 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1748 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2300 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1605641404
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4784 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1605641404
transform 1 0 3404 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1605641404
transform 1 0 4508 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1605641404
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_32
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_40
timestamp 1605641404
transform 1 0 4784 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_23
timestamp 1605641404
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_34
timestamp 1605641404
transform 1 0 4232 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6624 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4968 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1605641404
transform 1 0 5796 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_59
timestamp 1605641404
transform 1 0 6532 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_56
timestamp 1605641404
transform 1 0 6256 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1605641404
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7820 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 8280 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_76
timestamp 1605641404
transform 1 0 8096 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1605641404
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_82
timestamp 1605641404
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8832 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1605641404
transform 1 0 9936 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1605641404
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1605641404
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_93
timestamp 1605641404
transform 1 0 9660 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_105
timestamp 1605641404
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_109
timestamp 1605641404
transform 1 0 11132 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10948 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_116
timestamp 1605641404
transform 1 0 11776 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_117
timestamp 1605641404
transform 1 0 11868 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1605641404
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12052 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12512 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1605641404
transform 1 0 13064 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13524 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1605641404
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_133
timestamp 1605641404
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1605641404
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 1605641404
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1605641404
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15180 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1605641404
transform 1 0 15456 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_162
timestamp 1605641404
transform 1 0 16008 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1605641404
transform 1 0 16376 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16008 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 17664 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1605641404
transform 1 0 16928 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 18216 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_178
timestamp 1605641404
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_170
timestamp 1605641404
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1605641404
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1605641404
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1605641404
transform 1 0 19320 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 20240 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1605641404
transform 1 0 19780 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19228 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_196
timestamp 1605641404
transform 1 0 19136 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_201
timestamp 1605641404
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_195
timestamp 1605641404
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_206
timestamp 1605641404
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1605641404
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1605641404
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1605641404
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_217
timestamp 1605641404
transform 1 0 21068 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1605641404
transform 1 0 2024 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1605641404
transform 1 0 1932 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_19
timestamp 1605641404
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1605641404
transform 1 0 3036 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_24
timestamp 1605641404
transform 1 0 3312 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1605641404
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1605641404
transform 1 0 4876 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1605641404
transform 1 0 6716 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5244 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 6440 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_54
timestamp 1605641404
transform 1 0 6072 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1605641404
transform 1 0 7728 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_70
timestamp 1605641404
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_81
timestamp 1605641404
transform 1 0 8556 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1605641404
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_102
timestamp 1605641404
transform 1 0 10488 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 11500 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_110
timestamp 1605641404
transform 1 0 11224 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1605641404
transform 1 0 13156 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13892 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1605641404
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_134
timestamp 1605641404
transform 1 0 13432 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_138
timestamp 1605641404
transform 1 0 13800 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1605641404
transform 1 0 16284 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1605641404
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1605641404
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1605641404
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 17756 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1605641404
transform 1 0 17296 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_174
timestamp 1605641404
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_179
timestamp 1605641404
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 19780 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1605641404
transform 1 0 18768 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_190
timestamp 1605641404
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1605641404
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1605641404
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1605641404
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1605641404
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2208 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_11
timestamp 1605641404
transform 1 0 2116 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 3220 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1605641404
transform 1 0 4416 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_21
timestamp 1605641404
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_32
timestamp 1605641404
transform 1 0 4048 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1605641404
transform 1 0 5520 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_45
timestamp 1605641404
transform 1 0 5244 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1605641404
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1605641404
transform 1 0 7820 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1605641404
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_82
timestamp 1605641404
transform 1 0 8648 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9016 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1605641404
transform 1 0 10672 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_102
timestamp 1605641404
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1605641404
transform 1 0 11500 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1605641404
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13432 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 14444 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1605641404
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_143
timestamp 1605641404
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14812 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15824 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_148
timestamp 1605641404
transform 1 0 14720 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_158
timestamp 1605641404
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1605641404
transform 1 0 16836 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1605641404
transform 1 0 18124 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1605641404
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_180
timestamp 1605641404
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_184
timestamp 1605641404
transform 1 0 18032 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1605641404
transform 1 0 20148 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 19136 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_194
timestamp 1605641404
transform 1 0 18952 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_205
timestamp 1605641404
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_216
timestamp 1605641404
transform 1 0 20976 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1605641404
transform 1 0 2024 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_9
timestamp 1605641404
transform 1 0 1932 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_19
timestamp 1605641404
transform 1 0 2852 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1605641404
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_25
timestamp 1605641404
transform 1 0 3404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1605641404
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1605641404
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1605641404
transform 1 0 6072 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1605641404
transform 1 0 5060 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1605641404
transform 1 0 6532 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1605641404
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_57
timestamp 1605641404
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7912 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_10_68
timestamp 1605641404
transform 1 0 7360 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1605641404
transform 1 0 10672 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1605641404
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1605641404
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12144 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_10_113
timestamp 1605641404
transform 1 0 11500 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_119
timestamp 1605641404
transform 1 0 12052 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13156 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_129
timestamp 1605641404
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_140
timestamp 1605641404
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1605641404
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16928 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_170
timestamp 1605641404
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1605641404
transform 1 0 20240 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 18584 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1605641404
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_206
timestamp 1605641404
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1605641404
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1605641404
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_218
timestamp 1605641404
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1748 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1605641404
transform 1 0 4600 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 3588 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_23
timestamp 1605641404
transform 1 0 3220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_36
timestamp 1605641404
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1605641404
transform 1 0 5612 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_47
timestamp 1605641404
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_58
timestamp 1605641404
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1605641404
transform 1 0 7820 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1605641404
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_82
timestamp 1605641404
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9108 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9936 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 8832 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1605641404
transform 1 0 10764 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1605641404
transform 1 0 11316 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_108
timestamp 1605641404
transform 1 0 11040 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1605641404
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14076 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_139
timestamp 1605641404
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1605641404
transform 1 0 15732 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1605641404
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_157
timestamp 1605641404
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_162
timestamp 1605641404
transform 1 0 16008 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1605641404
transform 1 0 17388 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1605641404
transform 1 0 18124 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1605641404
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1605641404
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_184
timestamp 1605641404
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1605641404
transform 1 0 19136 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 19688 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp 1605641404
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1605641404
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_218
timestamp 1605641404
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1605641404
transform 1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1605641404
transform 1 0 1932 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_18
timestamp 1605641404
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1605641404
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1605641404
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6440 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5060 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_12_52
timestamp 1605641404
transform 1 0 5888 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1605641404
transform 1 0 8096 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_74
timestamp 1605641404
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10580 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1605641404
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1605641404
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1605641404
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12420 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 14076 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_139
timestamp 1605641404
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_144
timestamp 1605641404
transform 1 0 14352 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16284 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1605641404
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1605641404
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 17388 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_12_174
timestamp 1605641404
transform 1 0 17112 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19044 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19780 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1605641404
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_201
timestamp 1605641404
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1605641404
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1605641404
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_218
timestamp 1605641404
transform 1 0 21160 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1656 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2852 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1840 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_6
timestamp 1605641404
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_17
timestamp 1605641404
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4324 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4416 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_28
timestamp 1605641404
transform 1 0 3680 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_22
timestamp 1605641404
transform 1 0 3128 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1605641404
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5980 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5428 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_45
timestamp 1605641404
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_56
timestamp 1605641404
transform 1 0 6256 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1605641404
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_62
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_51
timestamp 1605641404
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8740 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7912 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6900 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 7636 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_72
timestamp 1605641404
transform 1 0 7728 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_80
timestamp 1605641404
transform 1 0 8464 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_69
timestamp 1605641404
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10580 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10396 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1605641404
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1605641404
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_96
timestamp 1605641404
transform 1 0 9936 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_102
timestamp 1605641404
transform 1 0 10488 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12604 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11592 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11408 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1605641404
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1605641404
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_123
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_112
timestamp 1605641404
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_123
timestamp 1605641404
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13984 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14260 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12788 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_136
timestamp 1605641404
transform 1 0 13616 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1605641404
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 15456 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15640 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1605641404
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1605641404
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 17112 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16652 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1605641404
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_167
timestamp 1605641404
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1605641404
transform 1 0 17480 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1605641404
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_184
timestamp 1605641404
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_172
timestamp 1605641404
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 19136 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 19504 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18492 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_188
timestamp 1605641404
transform 1 0 18400 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_198
timestamp 1605641404
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1605641404
transform 1 0 18584 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1605641404
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_216
timestamp 1605641404
transform 1 0 20976 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1605641404
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1605641404
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1605641404
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1840 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1605641404
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1605641404
transform 1 0 3496 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4140 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1605641404
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_29
timestamp 1605641404
transform 1 0 3772 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1605641404
transform 1 0 5796 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_49
timestamp 1605641404
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_54
timestamp 1605641404
transform 1 0 6072 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1605641404
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_78
timestamp 1605641404
transform 1 0 8280 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10488 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8832 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_100
timestamp 1605641404
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1605641404
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 14076 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_139
timestamp 1605641404
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1605641404
transform 1 0 16100 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15088 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_150
timestamp 1605641404
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_161
timestamp 1605641404
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1605641404
transform 1 0 17112 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1605641404
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_172
timestamp 1605641404
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_177
timestamp 1605641404
transform 1 0 17388 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1605641404
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 18492 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1605641404
transform 1 0 20148 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_188
timestamp 1605641404
transform 1 0 18400 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_205
timestamp 1605641404
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_216
timestamp 1605641404
transform 1 0 20976 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2024 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1605641404
transform 1 0 1932 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1605641404
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 3036 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4784 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1605641404
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_32
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6440 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_49
timestamp 1605641404
transform 1 0 5612 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_57
timestamp 1605641404
transform 1 0 6348 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1605641404
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7452 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_67
timestamp 1605641404
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_78
timestamp 1605641404
transform 1 0 8280 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1605641404
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_102
timestamp 1605641404
transform 1 0 10488 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 11132 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_108
timestamp 1605641404
transform 1 0 11040 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1605641404
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12788 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13800 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_136
timestamp 1605641404
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1605641404
transform 1 0 15824 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 14812 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1605641404
transform 1 0 15548 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_147
timestamp 1605641404
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1605641404
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 17112 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_169
timestamp 1605641404
transform 1 0 16652 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_173
timestamp 1605641404
transform 1 0 17020 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1605641404
transform 1 0 20240 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1605641404
transform 1 0 19136 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1605641404
transform 1 0 18584 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_205
timestamp 1605641404
transform 1 0 19964 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1605641404
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1605641404
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1605641404
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_218
timestamp 1605641404
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1605641404
transform 1 0 1932 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1605641404
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_18
timestamp 1605641404
transform 1 0 2760 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 3312 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_40
timestamp 1605641404
transform 1 0 4784 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_53
timestamp 1605641404
transform 1 0 5980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7084 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1605641404
transform 1 0 8740 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1605641404
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1605641404
transform 1 0 10672 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_92
timestamp 1605641404
transform 1 0 9568 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1605641404
transform 1 0 11868 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1605641404
transform 1 0 11500 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1605641404
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 13432 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1605641404
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_143
timestamp 1605641404
transform 1 0 14260 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16284 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15272 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_151
timestamp 1605641404
transform 1 0 14996 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_163
timestamp 1605641404
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1605641404
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1605641404
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1605641404
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 19596 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_193
timestamp 1605641404
transform 1 0 18860 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_217
timestamp 1605641404
transform 1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1605641404
transform 1 0 1472 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1605641404
transform 1 0 2024 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_8
timestamp 1605641404
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_19
timestamp 1605641404
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 3036 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1605641404
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1605641404
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5060 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1605641404
transform 1 0 6716 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1605641404
transform 1 0 6532 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7912 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_70
timestamp 1605641404
transform 1 0 7544 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_83
timestamp 1605641404
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10672 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1605641404
transform 1 0 8924 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1605641404
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1605641404
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1605641404
transform 1 0 11684 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1605641404
transform 1 0 12512 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1605641404
transform 1 0 12236 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_113
timestamp 1605641404
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_118
timestamp 1605641404
transform 1 0 11960 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1605641404
transform 1 0 13524 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_133
timestamp 1605641404
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_138
timestamp 1605641404
transform 1 0 13800 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1605641404
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_163
timestamp 1605641404
transform 1 0 16100 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16836 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1605641404
transform 1 0 17848 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_180
timestamp 1605641404
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1605641404
transform 1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1605641404
transform 1 0 19596 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1605641404
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_191
timestamp 1605641404
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_196
timestamp 1605641404
transform 1 0 19136 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1605641404
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1605641404
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1605641404
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1605641404
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1605641404
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1748 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1605641404
transform 1 0 1932 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_18
timestamp 1605641404
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_16
timestamp 1605641404
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 2760 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4140 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4692 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_34
timestamp 1605641404
transform 1 0 4232 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_38
timestamp 1605641404
transform 1 0 4600 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1605641404
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_32
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6624 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5704 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_48
timestamp 1605641404
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1605641404
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_49
timestamp 1605641404
transform 1 0 5612 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_57
timestamp 1605641404
transform 1 0 6348 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8648 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7636 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_78
timestamp 1605641404
transform 1 0 8280 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_69
timestamp 1605641404
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1605641404
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10672 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 9752 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_98
timestamp 1605641404
transform 1 0 10120 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12512 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11408 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1605641404
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_123
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1605641404
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_121
timestamp 1605641404
transform 1 0 12236 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 13524 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12880 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 13892 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_127
timestamp 1605641404
transform 1 0 12788 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_137
timestamp 1605641404
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 1605641404
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15272 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15548 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_148
timestamp 1605641404
transform 1 0 14720 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1605641404
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_166
timestamp 1605641404
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 17848 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16560 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16928 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1605641404
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1605641404
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1605641404
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_177
timestamp 1605641404
transform 1 0 17388 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_181
timestamp 1605641404
transform 1 0 17756 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18860 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19780 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_19_190
timestamp 1605641404
transform 1 0 18584 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_198
timestamp 1605641404
transform 1 0 19320 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_202
timestamp 1605641404
transform 1 0 19688 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20516 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1605641404
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_209
timestamp 1605641404
transform 1 0 20332 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_217
timestamp 1605641404
transform 1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1605641404
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1605641404
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1605641404
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1605641404
transform 1 0 2392 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2944 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1656 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1605641404
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_18
timestamp 1605641404
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4600 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_36
timestamp 1605641404
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_47
timestamp 1605641404
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1605641404
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1605641404
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6992 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_73
timestamp 1605641404
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_78
timestamp 1605641404
transform 1 0 8280 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1605641404
transform 1 0 10304 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_90
timestamp 1605641404
transform 1 0 9384 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_98
timestamp 1605641404
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11316 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_109
timestamp 1605641404
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_117
timestamp 1605641404
transform 1 0 11868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1605641404
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1605641404
transform 1 0 14444 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12788 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_143
timestamp 1605641404
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15272 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_21_148
timestamp 1605641404
transform 1 0 14720 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16928 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1605641404
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_170
timestamp 1605641404
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1605641404
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1605641404
transform 1 0 18952 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20240 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19504 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_190
timestamp 1605641404
transform 1 0 18584 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_198
timestamp 1605641404
transform 1 0 19320 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1605641404
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_214
timestamp 1605641404
transform 1 0 20792 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1605641404
transform 1 0 2576 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1840 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1605641404
transform 1 0 1748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_14
timestamp 1605641404
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_25
timestamp 1605641404
transform 1 0 3404 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 6348 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1605641404
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_56
timestamp 1605641404
transform 1 0 6256 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7728 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_63
timestamp 1605641404
transform 1 0 6900 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_71
timestamp 1605641404
transform 1 0 7636 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1605641404
transform 1 0 10304 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1605641404
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1605641404
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_93
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_99
timestamp 1605641404
transform 1 0 10212 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11316 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_109
timestamp 1605641404
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12972 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_127
timestamp 1605641404
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1605641404
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16100 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_154
timestamp 1605641404
transform 1 0 15272 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_162
timestamp 1605641404
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 17756 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_179
timestamp 1605641404
transform 1 0 17572 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1605641404
transform 1 0 20240 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1605641404
transform 1 0 19688 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1605641404
transform 1 0 19228 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_201
timestamp 1605641404
transform 1 0 19596 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1605641404
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1605641404
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1605641404
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1605641404
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1605641404
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1605641404
transform 1 0 2852 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1605641404
transform 1 0 2300 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1605641404
transform 1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1605641404
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1605641404
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_17
timestamp 1605641404
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1605641404
transform 1 0 3404 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1605641404
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_29
timestamp 1605641404
transform 1 0 3772 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_41
timestamp 1605641404
transform 1 0 4876 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1605641404
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1605641404
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1605641404
transform 1 0 6348 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1605641404
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1605641404
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1605641404
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1605641404
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1605641404
transform 1 0 11592 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1605641404
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_110
timestamp 1605641404
transform 1 0 11224 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1605641404
transform 1 0 11960 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1605641404
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 13616 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_135
timestamp 1605641404
transform 1 0 13524 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_145
timestamp 1605641404
transform 1 0 14444 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_157
timestamp 1605641404
transform 1 0 15548 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1605641404
transform 1 0 16928 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1605641404
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_169
timestamp 1605641404
transform 1 0 16652 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_175
timestamp 1605641404
transform 1 0 17204 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1605641404
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1605641404
transform 1 0 19412 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1605641404
transform 1 0 19964 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_196
timestamp 1605641404
transform 1 0 19136 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_203
timestamp 1605641404
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1605641404
transform 1 0 20516 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1605641404
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1605641404
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1605641404
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1605641404
transform 1 0 2300 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1605641404
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1605641404
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1605641404
transform 1 0 2116 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_17
timestamp 1605641404
transform 1 0 2668 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1605641404
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1605641404
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_38
timestamp 1605641404
transform 1 0 4600 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_50
timestamp 1605641404
transform 1 0 5704 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_62
timestamp 1605641404
transform 1 0 6808 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_74
timestamp 1605641404
transform 1 0 7912 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1605641404
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_86
timestamp 1605641404
transform 1 0 9016 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1605641404
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1605641404
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1605641404
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13432 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_129
timestamp 1605641404
transform 1 0 12972 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_133
timestamp 1605641404
transform 1 0 13340 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_140
timestamp 1605641404
transform 1 0 13984 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1605641404
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1605641404
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1605641404
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1605641404
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1605641404
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1605641404
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1605641404
transform 1 0 19688 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1605641404
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1605641404
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1605641404
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1605641404
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1605641404
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1605641404
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1605641404
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1605641404
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1605641404
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_11
timestamp 1605641404
transform 1 0 2116 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1605641404
transform 1 0 3496 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_23
timestamp 1605641404
transform 1 0 3220 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_30
timestamp 1605641404
transform 1 0 3864 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1605641404
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_42
timestamp 1605641404
transform 1 0 4968 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_54
timestamp 1605641404
transform 1 0 6072 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1605641404
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1605641404
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1605641404
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1605641404
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1605641404
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1605641404
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1605641404
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1605641404
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1605641404
transform 1 0 14352 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1605641404
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_143
timestamp 1605641404
transform 1 0 14260 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_148
timestamp 1605641404
transform 1 0 14720 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_160
timestamp 1605641404
transform 1 0 15824 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1605641404
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_172
timestamp 1605641404
transform 1 0 16928 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1605641404
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1605641404
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1605641404
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_208
timestamp 1605641404
transform 1 0 20240 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1605641404
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1605641404
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1605641404
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1605641404
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1605641404
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1605641404
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1605641404
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1605641404
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1605641404
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_11
timestamp 1605641404
transform 1 0 2116 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1605641404
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1605641404
transform 1 0 2116 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1605641404
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1605641404
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1605641404
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1605641404
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1605641404
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1605641404
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1605641404
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1605641404
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_47
timestamp 1605641404
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1605641404
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1605641404
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1605641404
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1605641404
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1605641404
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1605641404
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1605641404
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1605641404
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1605641404
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1605641404
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1605641404
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1605641404
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1605641404
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1605641404
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1605641404
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1605641404
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1605641404
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1605641404
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1605641404
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1605641404
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1605641404
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1605641404
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1605641404
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1605641404
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1605641404
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1605641404
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1605641404
transform 1 0 19964 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1605641404
transform 1 0 20240 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1605641404
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_202
timestamp 1605641404
transform 1 0 19688 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_196
timestamp 1605641404
transform 1 0 19136 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_204
timestamp 1605641404
transform 1 0 19872 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1605641404
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1605641404
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1605641404
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1605641404
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1605641404
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1605641404
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1605641404
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1605641404
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1605641404
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1605641404
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1605641404
transform 1 0 1564 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2116 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1605641404
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1605641404
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_9
timestamp 1605641404
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_17
timestamp 1605641404
transform 1 0 2668 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1605641404
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1605641404
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1605641404
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1605641404
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1605641404
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1605641404
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1605641404
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1605641404
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1605641404
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1605641404
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1605641404
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1605641404
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1605641404
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1605641404
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1605641404
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1605641404
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1605641404
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19596 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_190
timestamp 1605641404
transform 1 0 18584 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_198
timestamp 1605641404
transform 1 0 19320 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_207
timestamp 1605641404
transform 1 0 20148 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1605641404
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1605641404
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1605641404
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1605641404
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1605641404
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1605641404
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1605641404
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1605641404
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_11
timestamp 1605641404
transform 1 0 2116 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_23
timestamp 1605641404
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_35
timestamp 1605641404
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1605641404
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_47
timestamp 1605641404
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1605641404
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1605641404
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1605641404
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1605641404
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1605641404
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1605641404
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1605641404
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1605641404
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1605641404
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1605641404
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1605641404
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1605641404
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1605641404
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1605641404
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1605641404
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_208
timestamp 1605641404
transform 1 0 20240 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1605641404
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1605641404
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1605641404
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1605641404
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1605641404
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1605641404
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1605641404
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_11
timestamp 1605641404
transform 1 0 2116 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1605641404
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_23
timestamp 1605641404
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1605641404
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1605641404
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1605641404
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1605641404
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1605641404
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1605641404
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1605641404
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1605641404
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1605641404
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1605641404
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1605641404
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1605641404
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1605641404
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1605641404
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17572 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_178
timestamp 1605641404
transform 1 0 17480 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_185
timestamp 1605641404
transform 1 0 18124 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1605641404
transform 1 0 19228 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1605641404
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1605641404
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_209
timestamp 1605641404
transform 1 0 20332 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1605641404
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1605641404
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1605641404
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1605641404
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1605641404
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1605641404
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1605641404
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1605641404
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_17
timestamp 1605641404
transform 1 0 2668 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_29
timestamp 1605641404
transform 1 0 3772 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_41
timestamp 1605641404
transform 1 0 4876 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1605641404
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_53
timestamp 1605641404
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1605641404
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1605641404
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1605641404
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1605641404
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1605641404
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1605641404
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1605641404
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1605641404
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1605641404
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1605641404
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1605641404
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1605641404
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 1605641404
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1605641404
transform 1 0 18492 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_188
timestamp 1605641404
transform 1 0 18400 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1605641404
transform 1 0 18860 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_205
timestamp 1605641404
transform 1 0 19964 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1605641404
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1605641404
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1605641404
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1605641404
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1605641404
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1605641404
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1605641404
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1605641404
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1605641404
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1605641404
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1605641404
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1605641404
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1605641404
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1605641404
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1605641404
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1605641404
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1605641404
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1605641404
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1605641404
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1605641404
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1605641404
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1605641404
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1605641404
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1605641404
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1605641404
transform 1 0 14812 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1605641404
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1605641404
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1605641404
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1605641404
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1605641404
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1605641404
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1605641404
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1605641404
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_211
timestamp 1605641404
transform 1 0 20516 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1605641404
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 0 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_43_
port 1 nsew default input
rlabel metal2 s 1122 0 1178 480 6 bottom_left_grid_pin_44_
port 2 nsew default input
rlabel metal2 s 1582 0 1638 480 6 bottom_left_grid_pin_45_
port 3 nsew default input
rlabel metal2 s 2042 0 2098 480 6 bottom_left_grid_pin_46_
port 4 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_47_
port 5 nsew default input
rlabel metal2 s 3054 0 3110 480 6 bottom_left_grid_pin_48_
port 6 nsew default input
rlabel metal2 s 3514 0 3570 480 6 bottom_left_grid_pin_49_
port 7 nsew default input
rlabel metal2 s 11334 22320 11390 22800 6 ccff_head
port 8 nsew default input
rlabel metal2 s 18970 22320 19026 22800 6 ccff_tail
port 9 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[10]
port 11 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[11]
port 12 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[12]
port 13 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[13]
port 14 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[14]
port 15 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[15]
port 16 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[16]
port 17 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[17]
port 18 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[18]
port 19 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[19]
port 20 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[1]
port 21 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[2]
port 22 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[3]
port 23 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[4]
port 24 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[5]
port 25 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[6]
port 26 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[7]
port 27 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[8]
port 28 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[9]
port 29 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_out[0]
port 30 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[10]
port 31 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[11]
port 32 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[12]
port 33 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[13]
port 34 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[14]
port 35 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[15]
port 36 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[16]
port 37 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[17]
port 38 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[18]
port 39 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[19]
port 40 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[1]
port 41 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[2]
port 42 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[3]
port 43 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[4]
port 44 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[5]
port 45 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[6]
port 46 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[7]
port 47 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[8]
port 48 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[9]
port 49 nsew default tristate
rlabel metal3 s 22320 3816 22800 3936 6 chanx_right_in[0]
port 50 nsew default input
rlabel metal3 s 22320 8440 22800 8560 6 chanx_right_in[10]
port 51 nsew default input
rlabel metal3 s 22320 8984 22800 9104 6 chanx_right_in[11]
port 52 nsew default input
rlabel metal3 s 22320 9392 22800 9512 6 chanx_right_in[12]
port 53 nsew default input
rlabel metal3 s 22320 9936 22800 10056 6 chanx_right_in[13]
port 54 nsew default input
rlabel metal3 s 22320 10344 22800 10464 6 chanx_right_in[14]
port 55 nsew default input
rlabel metal3 s 22320 10752 22800 10872 6 chanx_right_in[15]
port 56 nsew default input
rlabel metal3 s 22320 11296 22800 11416 6 chanx_right_in[16]
port 57 nsew default input
rlabel metal3 s 22320 11704 22800 11824 6 chanx_right_in[17]
port 58 nsew default input
rlabel metal3 s 22320 12248 22800 12368 6 chanx_right_in[18]
port 59 nsew default input
rlabel metal3 s 22320 12656 22800 12776 6 chanx_right_in[19]
port 60 nsew default input
rlabel metal3 s 22320 4224 22800 4344 6 chanx_right_in[1]
port 61 nsew default input
rlabel metal3 s 22320 4768 22800 4888 6 chanx_right_in[2]
port 62 nsew default input
rlabel metal3 s 22320 5176 22800 5296 6 chanx_right_in[3]
port 63 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 chanx_right_in[4]
port 64 nsew default input
rlabel metal3 s 22320 6128 22800 6248 6 chanx_right_in[5]
port 65 nsew default input
rlabel metal3 s 22320 6672 22800 6792 6 chanx_right_in[6]
port 66 nsew default input
rlabel metal3 s 22320 7080 22800 7200 6 chanx_right_in[7]
port 67 nsew default input
rlabel metal3 s 22320 7488 22800 7608 6 chanx_right_in[8]
port 68 nsew default input
rlabel metal3 s 22320 8032 22800 8152 6 chanx_right_in[9]
port 69 nsew default input
rlabel metal3 s 22320 13200 22800 13320 6 chanx_right_out[0]
port 70 nsew default tristate
rlabel metal3 s 22320 17824 22800 17944 6 chanx_right_out[10]
port 71 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[11]
port 72 nsew default tristate
rlabel metal3 s 22320 18776 22800 18896 6 chanx_right_out[12]
port 73 nsew default tristate
rlabel metal3 s 22320 19184 22800 19304 6 chanx_right_out[13]
port 74 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 chanx_right_out[14]
port 75 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[15]
port 76 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 chanx_right_out[16]
port 77 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[17]
port 78 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[18]
port 79 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 chanx_right_out[19]
port 80 nsew default tristate
rlabel metal3 s 22320 13608 22800 13728 6 chanx_right_out[1]
port 81 nsew default tristate
rlabel metal3 s 22320 14016 22800 14136 6 chanx_right_out[2]
port 82 nsew default tristate
rlabel metal3 s 22320 14560 22800 14680 6 chanx_right_out[3]
port 83 nsew default tristate
rlabel metal3 s 22320 14968 22800 15088 6 chanx_right_out[4]
port 84 nsew default tristate
rlabel metal3 s 22320 15512 22800 15632 6 chanx_right_out[5]
port 85 nsew default tristate
rlabel metal3 s 22320 15920 22800 16040 6 chanx_right_out[6]
port 86 nsew default tristate
rlabel metal3 s 22320 16464 22800 16584 6 chanx_right_out[7]
port 87 nsew default tristate
rlabel metal3 s 22320 16872 22800 16992 6 chanx_right_out[8]
port 88 nsew default tristate
rlabel metal3 s 22320 17280 22800 17400 6 chanx_right_out[9]
port 89 nsew default tristate
rlabel metal2 s 3974 0 4030 480 6 chany_bottom_in[0]
port 90 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chany_bottom_in[10]
port 91 nsew default input
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_in[11]
port 92 nsew default input
rlabel metal2 s 9678 0 9734 480 6 chany_bottom_in[12]
port 93 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[13]
port 94 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[14]
port 95 nsew default input
rlabel metal2 s 11058 0 11114 480 6 chany_bottom_in[15]
port 96 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_in[16]
port 97 nsew default input
rlabel metal2 s 12070 0 12126 480 6 chany_bottom_in[17]
port 98 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[18]
port 99 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[19]
port 100 nsew default input
rlabel metal2 s 4434 0 4490 480 6 chany_bottom_in[1]
port 101 nsew default input
rlabel metal2 s 4894 0 4950 480 6 chany_bottom_in[2]
port 102 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_in[3]
port 103 nsew default input
rlabel metal2 s 5906 0 5962 480 6 chany_bottom_in[4]
port 104 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[5]
port 105 nsew default input
rlabel metal2 s 6826 0 6882 480 6 chany_bottom_in[6]
port 106 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[7]
port 107 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[8]
port 108 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[9]
port 109 nsew default input
rlabel metal2 s 13450 0 13506 480 6 chany_bottom_out[0]
port 110 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[10]
port 111 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 chany_bottom_out[11]
port 112 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chany_bottom_out[12]
port 113 nsew default tristate
rlabel metal2 s 19614 0 19670 480 6 chany_bottom_out[13]
port 114 nsew default tristate
rlabel metal2 s 20166 0 20222 480 6 chany_bottom_out[14]
port 115 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 chany_bottom_out[15]
port 116 nsew default tristate
rlabel metal2 s 21086 0 21142 480 6 chany_bottom_out[16]
port 117 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[17]
port 118 nsew default tristate
rlabel metal2 s 22006 0 22062 480 6 chany_bottom_out[18]
port 119 nsew default tristate
rlabel metal2 s 22466 0 22522 480 6 chany_bottom_out[19]
port 120 nsew default tristate
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_out[1]
port 121 nsew default tristate
rlabel metal2 s 14462 0 14518 480 6 chany_bottom_out[2]
port 122 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_out[3]
port 123 nsew default tristate
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_out[4]
port 124 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[5]
port 125 nsew default tristate
rlabel metal2 s 16302 0 16358 480 6 chany_bottom_out[6]
port 126 nsew default tristate
rlabel metal2 s 16762 0 16818 480 6 chany_bottom_out[7]
port 127 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_out[8]
port 128 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_out[9]
port 129 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 130 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 131 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_36_
port 132 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 133 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_38_
port 134 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 135 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_40_
port 136 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 137 nsew default input
rlabel metal3 s 0 22448 480 22568 6 left_top_grid_pin_1_
port 138 nsew default input
rlabel metal2 s 3790 22320 3846 22800 6 prog_clk
port 139 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_34_
port 140 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_35_
port 141 nsew default input
rlabel metal3 s 22320 960 22800 1080 6 right_bottom_grid_pin_36_
port 142 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_37_
port 143 nsew default input
rlabel metal3 s 22320 1912 22800 2032 6 right_bottom_grid_pin_38_
port 144 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_39_
port 145 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_40_
port 146 nsew default input
rlabel metal3 s 22320 3408 22800 3528 6 right_bottom_grid_pin_41_
port 147 nsew default input
rlabel metal3 s 22320 22448 22800 22568 6 right_top_grid_pin_1_
port 148 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 149 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
