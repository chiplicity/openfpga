* NGSPICE file created from sb_3__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt sb_3__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ chanx_left_in[0] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4]
+ chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chany_top_in[0] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1] chany_top_out[2]
+ chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7]
+ chany_top_out[8] data_in enable left_bottom_grid_pin_11_ left_bottom_grid_pin_13_
+ left_bottom_grid_pin_15_ left_bottom_grid_pin_1_ left_bottom_grid_pin_3_ left_bottom_grid_pin_5_
+ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_ left_top_grid_pin_10_ top_left_grid_pin_13_
+ top_right_grid_pin_11_ top_right_grid_pin_13_ top_right_grid_pin_15_ top_right_grid_pin_1_
+ top_right_grid_pin_3_ top_right_grid_pin_5_ top_right_grid_pin_7_ top_right_grid_pin_9_
+ vpwr vgnd
XFILLER_36_19 vgnd vpwr scs8hd_decap_6
XFILLER_22_100 vpwr vgnd scs8hd_fill_2
XFILLER_22_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_7 vgnd vpwr scs8hd_decap_12
XFILLER_26_30 vgnd vpwr scs8hd_fill_1
XFILLER_26_85 vpwr vgnd scs8hd_fill_2
XFILLER_42_40 vgnd vpwr scs8hd_decap_4
XFILLER_9_159 vgnd vpwr scs8hd_decap_12
XFILLER_36_236 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_7_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XFILLER_12_10 vgnd vpwr scs8hd_decap_4
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_239 vgnd vpwr scs8hd_decap_4
XANTENNA__108__B enable vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _190_/A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_209 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_42 vpwr vgnd scs8hd_fill_2
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_23_75 vpwr vgnd scs8hd_fill_2
X_131_ _129_/X _133_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XANTENNA__110__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA__119__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
X_114_ _113_/Y _115_/B vgnd vpwr scs8hd_buf_1
XFILLER_22_7 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _217_/HI _172_/Y mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_32 vpwr vgnd scs8hd_fill_2
XFILLER_20_43 vgnd vpwr scs8hd_decap_8
Xmux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _214_/HI _194_/Y mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_30 vpwr vgnd scs8hd_fill_2
XFILLER_29_52 vpwr vgnd scs8hd_fill_2
XFILLER_29_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_194 vgnd vpwr scs8hd_decap_8
XANTENNA__116__B _117_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XANTENNA__132__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_25_120 vpwr vgnd scs8hd_fill_2
XFILLER_40_167 vgnd vpwr scs8hd_fill_1
XFILLER_40_145 vgnd vpwr scs8hd_decap_8
XFILLER_31_75 vpwr vgnd scs8hd_fill_2
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XFILLER_31_123 vgnd vpwr scs8hd_decap_4
XANTENNA__127__A _096_/X vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_223 vpwr vgnd scs8hd_fill_2
XFILLER_39_212 vpwr vgnd scs8hd_fill_2
XFILLER_39_201 vpwr vgnd scs8hd_fill_2
XFILLER_22_145 vpwr vgnd scs8hd_fill_2
Xmem_top_track_4.LATCH_0_.latch data_in _177_/A _117_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XFILLER_42_63 vgnd vpwr scs8hd_decap_8
XFILLER_36_248 vgnd vpwr scs8hd_decap_12
XFILLER_36_215 vgnd vpwr scs8hd_decap_4
XFILLER_27_204 vgnd vpwr scs8hd_decap_12
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XANTENNA__230__A _230_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.tap_buf4_0_.scs8hd_inv_1 mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _206_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XANTENNA__124__B _124_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XANTENNA__140__A _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_251 vpwr vgnd scs8hd_fill_2
Xmux_top_track_6.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_5_ mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
X_130_ _123_/A _115_/B _100_/A _169_/A _133_/B vgnd vpwr scs8hd_or4_4
XANTENNA__110__D _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XANTENNA__119__B _120_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
XANTENNA__135__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_5.tap_buf4_0_.scs8hd_inv_1 mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _232_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_10 vpwr vgnd scs8hd_fill_2
XFILLER_34_42 vgnd vpwr scs8hd_decap_4
XFILLER_11_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd vpwr
+ scs8hd_diode_2
X_113_ address[2] _113_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_7 vgnd vpwr scs8hd_decap_4
Xmux_top_track_6.tap_buf4_0_.scs8hd_inv_1 mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_22 vgnd vpwr scs8hd_decap_8
XFILLER_20_88 vpwr vgnd scs8hd_fill_2
XFILLER_28_162 vgnd vpwr scs8hd_decap_4
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _193_/A mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_187 vgnd vpwr scs8hd_decap_4
Xmem_left_track_5.LATCH_1_.latch data_in _194_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_11 vgnd vpwr scs8hd_fill_1
XFILLER_15_22 vgnd vpwr scs8hd_decap_4
XFILLER_15_33 vpwr vgnd scs8hd_fill_2
XFILLER_15_44 vgnd vpwr scs8hd_decap_4
XFILLER_15_55 vgnd vpwr scs8hd_decap_6
XFILLER_15_66 vgnd vpwr scs8hd_decap_4
XFILLER_25_187 vpwr vgnd scs8hd_fill_2
XFILLER_31_98 vpwr vgnd scs8hd_fill_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XANTENNA__233__A _233_/A vgnd vpwr scs8hd_diode_2
XANTENNA__127__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
XFILLER_31_168 vpwr vgnd scs8hd_fill_2
XFILLER_31_102 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_15_ mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vgnd vpwr scs8hd_decap_12
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_168 vgnd vpwr scs8hd_decap_4
Xmux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _175_/Y mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_26_32 vpwr vgnd scs8hd_fill_2
XFILLER_42_53 vgnd vpwr scs8hd_decap_8
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_43 vpwr vgnd scs8hd_fill_2
XANTENNA__138__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_12_190 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _197_/Y mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_27_216 vgnd vpwr scs8hd_decap_12
XFILLER_10_105 vgnd vpwr scs8hd_decap_12
XFILLER_12_56 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_75 vpwr vgnd scs8hd_fill_2
XFILLER_37_53 vpwr vgnd scs8hd_fill_2
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XFILLER_41_230 vgnd vpwr scs8hd_decap_12
XANTENNA__140__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XANTENNA__241__A _241_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__135__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_3
XANTENNA__151__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _175_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_211 vgnd vpwr scs8hd_decap_3
XFILLER_18_44 vgnd vpwr scs8hd_decap_3
XFILLER_34_21 vgnd vpwr scs8hd_decap_8
XFILLER_18_88 vpwr vgnd scs8hd_fill_2
XFILLER_34_65 vgnd vpwr scs8hd_decap_8
X_112_ _117_/A _111_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__236__A _236_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_3_ mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__146__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_37_174 vpwr vgnd scs8hd_fill_2
XFILLER_34_122 vpwr vgnd scs8hd_fill_2
XFILLER_19_130 vgnd vpwr scs8hd_decap_4
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XFILLER_40_158 vgnd vpwr scs8hd_decap_3
XFILLER_25_100 vpwr vgnd scs8hd_fill_2
XFILLER_25_144 vpwr vgnd scs8hd_fill_2
XFILLER_16_166 vgnd vpwr scs8hd_decap_12
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_180 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_22 vpwr vgnd scs8hd_fill_2
XFILLER_26_66 vpwr vgnd scs8hd_fill_2
XFILLER_13_147 vgnd vpwr scs8hd_decap_12
XANTENNA__138__B _137_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _164_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _177_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_13_ mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_228 vgnd vpwr scs8hd_decap_12
XFILLER_10_117 vgnd vpwr scs8hd_decap_12
XFILLER_5_7 vgnd vpwr scs8hd_decap_12
XFILLER_37_21 vpwr vgnd scs8hd_fill_2
XFILLER_41_242 vpwr vgnd scs8hd_fill_2
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _225_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XFILLER_38_7 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_0_.latch data_in _173_/A _107_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_15.LATCH_0_.latch data_in _205_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__140__C _157_/C vgnd vpwr scs8hd_diode_2
XANTENNA__149__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XFILLER_23_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_188_ _188_/A _188_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__151__B _149_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_23 vpwr vgnd scs8hd_fill_2
XFILLER_18_67 vgnd vpwr scs8hd_decap_4
X_111_ _096_/X _111_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
XANTENNA__146__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_120 vpwr vgnd scs8hd_fill_2
XFILLER_29_109 vpwr vgnd scs8hd_fill_2
XFILLER_20_68 vgnd vpwr scs8hd_decap_4
XFILLER_29_77 vgnd vpwr scs8hd_decap_4
XFILLER_13_6 vpwr vgnd scs8hd_fill_2
XFILLER_19_120 vpwr vgnd scs8hd_fill_2
XFILLER_34_112 vgnd vpwr scs8hd_fill_1
XANTENNA__157__A _123_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_1_ mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_123 vgnd vpwr scs8hd_decap_4
XFILLER_25_178 vgnd vpwr scs8hd_decap_4
XFILLER_31_56 vgnd vpwr scs8hd_decap_3
XFILLER_31_34 vpwr vgnd scs8hd_fill_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XFILLER_16_112 vgnd vpwr scs8hd_decap_12
XFILLER_16_178 vgnd vpwr scs8hd_decap_12
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__143__C _157_/C vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _192_/Y mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_104 vpwr vgnd scs8hd_fill_2
XFILLER_22_115 vgnd vpwr scs8hd_decap_4
XFILLER_22_126 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.LATCH_1_.latch data_in _190_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _207_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_104 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_89 vgnd vpwr scs8hd_decap_3
XFILLER_13_159 vgnd vpwr scs8hd_decap_12
XFILLER_8_141 vgnd vpwr scs8hd_decap_12
XANTENNA__154__B _153_/X vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_129 vgnd vpwr scs8hd_decap_12
XFILLER_12_69 vgnd vpwr scs8hd_decap_4
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
XANTENNA__140__D _160_/D vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_232 vgnd vpwr scs8hd_decap_12
XFILLER_23_46 vpwr vgnd scs8hd_fill_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_23_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_11_ mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_17 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A _187_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_35 vpwr vgnd scs8hd_fill_2
X_110_ _104_/A _123_/B _123_/C _171_/A _111_/B vgnd vpwr scs8hd_or4_4
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
X_239_ _239_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__146__C _157_/C vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_3
XANTENNA__162__B _162_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_143 vpwr vgnd scs8hd_fill_2
XFILLER_37_198 vpwr vgnd scs8hd_fill_2
XFILLER_37_187 vpwr vgnd scs8hd_fill_2
XFILLER_20_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_12 vpwr vgnd scs8hd_fill_2
XFILLER_29_34 vgnd vpwr scs8hd_decap_4
XFILLER_29_56 vgnd vpwr scs8hd_decap_3
XFILLER_28_132 vpwr vgnd scs8hd_fill_2
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XFILLER_42_190 vgnd vpwr scs8hd_decap_8
XFILLER_34_168 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _209_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__157__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_14 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_31_13 vpwr vgnd scs8hd_fill_2
XFILLER_31_79 vgnd vpwr scs8hd_decap_4
XFILLER_31_149 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_102 vgnd vpwr scs8hd_decap_8
XFILLER_16_124 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__D _157_/D vgnd vpwr scs8hd_diode_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_216 vgnd vpwr scs8hd_decap_4
XFILLER_39_205 vgnd vpwr scs8hd_decap_4
XFILLER_39_249 vpwr vgnd scs8hd_fill_2
XFILLER_39_227 vgnd vpwr scs8hd_decap_12
XANTENNA__168__A _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_149 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _191_/A mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_116 vgnd vpwr scs8hd_decap_6
XFILLER_26_79 vgnd vpwr scs8hd_decap_4
XFILLER_42_23 vgnd vpwr scs8hd_decap_8
XFILLER_21_182 vgnd vpwr scs8hd_fill_1
XFILLER_36_219 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__170__B _169_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_230 vpwr vgnd scs8hd_fill_2
XFILLER_37_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
Xmem_top_track_8.LATCH_1_.latch data_in _180_/A _124_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _173_/Y mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__149__C _157_/C vgnd vpwr scs8hd_diode_2
XANTENNA__165__B _164_/B vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_23_25 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _195_/Y mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_29 vpwr vgnd scs8hd_fill_2
XFILLER_13_80 vgnd vpwr scs8hd_decap_12
X_186_ _186_/A _186_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_11.LATCH_0_.latch data_in _201_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_58 vpwr vgnd scs8hd_fill_2
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
X_238_ _238_/A chany_top_out[5] vgnd vpwr scs8hd_buf_2
X_169_ _169_/A _169_/B _165_/A _169_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_11.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_9_ mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__146__D _160_/D vgnd vpwr scs8hd_diode_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_3
XFILLER_37_111 vpwr vgnd scs8hd_fill_2
XFILLER_1_50 vgnd vpwr scs8hd_decap_8
Xmux_left_track_7.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_177 vgnd vpwr scs8hd_decap_8
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__157__C _157_/C vgnd vpwr scs8hd_diode_2
XFILLER_25_114 vgnd vpwr scs8hd_decap_4
XFILLER_40_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_117 vpwr vgnd scs8hd_fill_2
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_136 vgnd vpwr scs8hd_decap_12
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_80 vpwr vgnd scs8hd_fill_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_239 vgnd vpwr scs8hd_decap_4
XANTENNA__168__B _169_/B vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_47 vpwr vgnd scs8hd_fill_2
XFILLER_21_161 vpwr vgnd scs8hd_fill_2
XFILLER_21_172 vpwr vgnd scs8hd_fill_2
Xmem_top_track_14.LATCH_0_.latch data_in _187_/A _136_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XANTENNA__170__C _164_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_242 vpwr vgnd scs8hd_fill_2
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.tap_buf4_0_.scs8hd_inv_1 mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _236_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_201 vgnd vpwr scs8hd_decap_12
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XANTENNA__149__D _157_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XFILLER_3_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XFILLER_13_92 vgnd vpwr scs8hd_decap_12
X_185_ _185_/A _185_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_36 vgnd vpwr scs8hd_decap_4
XFILLER_7_208 vgnd vpwr scs8hd_decap_12
X_237_ _237_/A chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_168_ _169_/A _169_/B _164_/A _168_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
X_099_ address[4] address[5] _100_/A vgnd vpwr scs8hd_or2_4
XFILLER_37_178 vgnd vpwr scs8hd_decap_4
XFILLER_37_156 vpwr vgnd scs8hd_fill_2
XFILLER_37_123 vgnd vpwr scs8hd_decap_3
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_112 vpwr vgnd scs8hd_fill_2
XFILLER_28_145 vgnd vpwr scs8hd_decap_6
XANTENNA__097__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_18 vgnd vpwr scs8hd_decap_12
XFILLER_10_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_126 vpwr vgnd scs8hd_fill_2
XFILLER_34_104 vpwr vgnd scs8hd_fill_2
XFILLER_19_112 vpwr vgnd scs8hd_fill_2
XFILLER_19_134 vgnd vpwr scs8hd_fill_1
XFILLER_19_156 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_90 vpwr vgnd scs8hd_fill_2
XANTENNA__157__D _157_/D vgnd vpwr scs8hd_diode_2
XFILLER_25_104 vgnd vpwr scs8hd_fill_1
XFILLER_25_159 vpwr vgnd scs8hd_fill_2
XFILLER_16_148 vgnd vpwr scs8hd_decap_4
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_170 vgnd vpwr scs8hd_decap_8
Xmux_left_track_5.INVTX1_0_.scs8hd_inv_1 chany_top_in[7] mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_6 vpwr vgnd scs8hd_fill_2
XANTENNA__168__C _164_/A vgnd vpwr scs8hd_diode_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
XFILLER_26_26 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_36 vpwr vgnd scs8hd_fill_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_19 vgnd vpwr scs8hd_decap_12
XFILLER_29_240 vgnd vpwr scs8hd_decap_4
XFILLER_32_91 vgnd vpwr scs8hd_fill_1
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XFILLER_16_81 vpwr vgnd scs8hd_fill_2
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_17 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _208_/HI _190_/Y mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_41_202 vpwr vgnd scs8hd_fill_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XFILLER_32_257 vgnd vpwr scs8hd_decap_12
XFILLER_32_213 vgnd vpwr scs8hd_fill_1
XFILLER_17_232 vgnd vpwr scs8hd_decap_12
XFILLER_27_91 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_202 vgnd vpwr scs8hd_decap_12
X_184_ _184_/A _184_/Y vgnd vpwr scs8hd_inv_8
Xmem_top_track_4.LATCH_1_.latch data_in _176_/A _116_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_227 vgnd vpwr scs8hd_decap_12
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_236_ _236_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
X_167_ _166_/X _169_/B vgnd vpwr scs8hd_buf_1
X_098_ address[2] _123_/B vgnd vpwr scs8hd_buf_1
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _206_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_157 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_149 vgnd vpwr scs8hd_decap_4
XFILLER_19_146 vgnd vpwr scs8hd_decap_8
XFILLER_19_168 vgnd vpwr scs8hd_decap_12
XFILLER_42_171 vgnd vpwr scs8hd_decap_12
XFILLER_42_160 vgnd vpwr scs8hd_decap_8
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_193 vpwr vgnd scs8hd_fill_2
XFILLER_18_190 vgnd vpwr scs8hd_decap_12
XFILLER_31_38 vgnd vpwr scs8hd_decap_3
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_160 vgnd vpwr scs8hd_fill_1
XFILLER_21_93 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_171 vgnd vpwr scs8hd_decap_12
XFILLER_30_163 vgnd vpwr scs8hd_decap_8
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_21_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
XFILLER_12_141 vgnd vpwr scs8hd_decap_12
XFILLER_35_222 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.INVTX1_0_.scs8hd_inv_1 chany_top_in[8] mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
Xmem_top_track_10.LATCH_0_.latch data_in _183_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_269 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _234_/A vgnd vpwr scs8hd_inv_1
XFILLER_4_30 vgnd vpwr scs8hd_fill_1
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.tap_buf4_0_.scs8hd_inv_1 mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _242_/A vgnd vpwr scs8hd_inv_1
XFILLER_9_19 vgnd vpwr scs8hd_decap_12
X_183_ _183_/A _183_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_20_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_39 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_6 vpwr vgnd scs8hd_fill_2
X_235_ _235_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_24_71 vpwr vgnd scs8hd_fill_2
XFILLER_40_70 vgnd vpwr scs8hd_decap_3
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_097_ address[3] _104_/A vgnd vpwr scs8hd_buf_1
Xmux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _193_/Y mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_166_ address[3] address[2] address[4] _137_/Y _166_/X vgnd vpwr scs8hd_or4_4
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_18 vpwr vgnd scs8hd_fill_2
XFILLER_29_16 vgnd vpwr scs8hd_decap_3
XFILLER_29_38 vgnd vpwr scs8hd_fill_1
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_139 vgnd vpwr scs8hd_decap_8
XFILLER_19_93 vpwr vgnd scs8hd_fill_2
XFILLER_42_183 vgnd vpwr scs8hd_decap_3
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
X_149_ address[3] _115_/B _157_/C _157_/D _149_/X vgnd vpwr scs8hd_or4_4
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_17 vpwr vgnd scs8hd_fill_2
XFILLER_15_18 vpwr vgnd scs8hd_fill_2
XFILLER_15_29 vpwr vgnd scs8hd_fill_2
XFILLER_0_249 vgnd vpwr scs8hd_decap_12
XFILLER_31_109 vgnd vpwr scs8hd_decap_6
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_150 vgnd vpwr scs8hd_decap_3
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_197 vgnd vpwr scs8hd_decap_12
XFILLER_30_186 vpwr vgnd scs8hd_fill_2
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XFILLER_21_142 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XFILLER_35_234 vgnd vpwr scs8hd_decap_8
XFILLER_37_38 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_29 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_182_ _182_/A _182_/Y vgnd vpwr scs8hd_inv_8
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_13_62 vgnd vpwr scs8hd_decap_3
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _100_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _177_/Y vgnd vpwr
+ scs8hd_diode_2
X_165_ _165_/A _164_/B _165_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_251 vgnd vpwr scs8hd_decap_12
X_234_ _234_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_24_83 vpwr vgnd scs8hd_fill_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_3
X_096_ _096_/A _096_/X vgnd vpwr scs8hd_buf_1
XFILLER_37_115 vgnd vpwr scs8hd_decap_3
XFILLER_1_10 vpwr vgnd scs8hd_fill_2
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_1_.latch data_in _172_/A _105_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_15.LATCH_1_.latch data_in _204_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_30 vgnd vpwr scs8hd_fill_1
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XFILLER_19_126 vpwr vgnd scs8hd_fill_2
XFILLER_35_71 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.INVTX1_1_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd vpwr
+ scs8hd_diode_2
X_148_ _133_/A _146_/X _148_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_3 vgnd vpwr scs8hd_decap_3
XFILLER_33_140 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_73 vgnd vpwr scs8hd_decap_4
XFILLER_30_121 vgnd vpwr scs8hd_fill_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XFILLER_7_86 vgnd vpwr scs8hd_decap_12
XFILLER_7_31 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_110 vpwr vgnd scs8hd_fill_2
XFILLER_26_18 vpwr vgnd scs8hd_fill_2
XFILLER_21_165 vpwr vgnd scs8hd_fill_2
XFILLER_21_176 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _183_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_154 vgnd vpwr scs8hd_decap_12
XFILLER_32_72 vgnd vpwr scs8hd_fill_1
XFILLER_32_50 vgnd vpwr scs8hd_fill_1
XANTENNA__103__A _160_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
XFILLER_35_202 vpwr vgnd scs8hd_fill_2
XFILLER_37_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _179_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
X_181_ _181_/A _181_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_3
XFILLER_9_220 vgnd vpwr scs8hd_decap_12
XFILLER_34_29 vpwr vgnd scs8hd_fill_2
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_40 vgnd vpwr scs8hd_fill_1
X_164_ _164_/A _164_/B _164_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_263 vgnd vpwr scs8hd_decap_12
X_233_ _233_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
X_095_ address[0] _096_/A vgnd vpwr scs8hd_inv_8
XFILLER_34_8 vgnd vpwr scs8hd_decap_4
XANTENNA__111__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_116 vgnd vpwr scs8hd_decap_3
XFILLER_34_108 vpwr vgnd scs8hd_fill_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_3
XFILLER_19_116 vpwr vgnd scs8hd_fill_2
XFILLER_27_193 vpwr vgnd scs8hd_fill_2
XANTENNA__106__A address[0] vgnd vpwr scs8hd_diode_2
X_147_ _129_/X _146_/X _147_/Y vgnd vpwr scs8hd_nor2_4
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_30 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _188_/A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_7_43 vgnd vpwr scs8hd_decap_12
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
XFILLER_7_98 vgnd vpwr scs8hd_decap_12
XFILLER_38_200 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.INVTX1_1_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _206_/A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_166 vgnd vpwr scs8hd_decap_12
XFILLER_16_85 vgnd vpwr scs8hd_decap_4
XFILLER_32_84 vgnd vpwr scs8hd_decap_4
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_41_206 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_17_269 vgnd vpwr scs8hd_decap_8
XFILLER_27_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA__114__A _113_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
X_180_ _180_/A _180_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_232 vgnd vpwr scs8hd_decap_12
XANTENNA__109__A _157_/D vgnd vpwr scs8hd_diode_2
X_232_ _232_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_24_52 vpwr vgnd scs8hd_fill_2
XFILLER_40_84 vgnd vpwr scs8hd_decap_8
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
X_163_ _122_/A _113_/Y _160_/C _157_/D _164_/B vgnd vpwr scs8hd_or4_4
XANTENNA__111__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_128 vpwr vgnd scs8hd_fill_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_19_74 vpwr vgnd scs8hd_fill_2
XFILLER_42_142 vgnd vpwr scs8hd_decap_12
XFILLER_42_131 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
X_146_ address[3] _115_/B _157_/C _160_/D _146_/X vgnd vpwr scs8hd_or4_4
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_197 vgnd vpwr scs8hd_decap_4
XFILLER_33_175 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _191_/Y mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_track_11.LATCH_1_.latch data_in _200_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_120 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_145 vgnd vpwr scs8hd_decap_8
XFILLER_7_55 vgnd vpwr scs8hd_decap_6
X_129_ _096_/A _129_/X vgnd vpwr scs8hd_buf_1
XFILLER_30_3 vpwr vgnd scs8hd_fill_2
XFILLER_38_212 vpwr vgnd scs8hd_fill_2
XFILLER_21_123 vpwr vgnd scs8hd_fill_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XFILLER_16_64 vpwr vgnd scs8hd_fill_2
XFILLER_32_41 vpwr vgnd scs8hd_fill_2
XFILLER_8_105 vgnd vpwr scs8hd_decap_12
XFILLER_12_178 vgnd vpwr scs8hd_decap_12
XFILLER_7_171 vgnd vpwr scs8hd_decap_12
XFILLER_41_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
Xmux_top_track_10.INVTX1_1_.scs8hd_inv_1 chanx_left_in[4] mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
Xmem_left_track_7.LATCH_0_.latch data_in _197_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XANTENNA__130__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_251 vgnd vpwr scs8hd_decap_12
XFILLER_13_10 vpwr vgnd scs8hd_fill_2
XFILLER_13_21 vpwr vgnd scs8hd_fill_2
XFILLER_13_43 vgnd vpwr scs8hd_decap_12
XFILLER_13_76 vpwr vgnd scs8hd_fill_2
XFILLER_38_84 vgnd vpwr scs8hd_decap_8
Xmem_top_track_14.LATCH_1_.latch data_in _186_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_170 vgnd vpwr scs8hd_fill_1
X_231_ _231_/A chanx_left_out[3] vgnd vpwr scs8hd_buf_2
X_162_ _165_/A _162_/B _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_75 vpwr vgnd scs8hd_fill_2
XFILLER_40_41 vgnd vpwr scs8hd_decap_3
XFILLER_40_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_37_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_42_154 vgnd vpwr scs8hd_fill_1
XFILLER_19_97 vgnd vpwr scs8hd_decap_4
XFILLER_27_151 vpwr vgnd scs8hd_fill_2
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
X_145_ _133_/A _143_/X _145_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_154 vpwr vgnd scs8hd_fill_2
XFILLER_33_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_132 vpwr vgnd scs8hd_fill_2
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_6
XFILLER_24_187 vgnd vpwr scs8hd_decap_12
XFILLER_30_135 vpwr vgnd scs8hd_fill_2
XFILLER_30_113 vpwr vgnd scs8hd_fill_2
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XANTENNA__117__B _117_/B vgnd vpwr scs8hd_diode_2
X_128_ _117_/A _127_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__133__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_10.tap_buf4_0_.scs8hd_inv_1 mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _238_/A vgnd vpwr scs8hd_inv_1
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_16_21 vgnd vpwr scs8hd_decap_4
XFILLER_16_32 vgnd vpwr scs8hd_decap_3
XFILLER_32_64 vpwr vgnd scs8hd_fill_2
XFILLER_8_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_42 vpwr vgnd scs8hd_fill_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_68 vgnd vpwr scs8hd_decap_12
XANTENNA__130__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_263 vgnd vpwr scs8hd_decap_12
XFILLER_13_55 vgnd vpwr scs8hd_decap_6
XFILLER_38_30 vgnd vpwr scs8hd_fill_1
XANTENNA__231__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XANTENNA__125__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_193 vpwr vgnd scs8hd_fill_2
XFILLER_39_160 vgnd vpwr scs8hd_decap_8
XFILLER_40_20 vpwr vgnd scs8hd_fill_2
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
X_230_ _230_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XFILLER_24_10 vpwr vgnd scs8hd_fill_2
XFILLER_24_32 vpwr vgnd scs8hd_fill_2
XFILLER_24_87 vgnd vpwr scs8hd_decap_3
X_161_ _164_/A _162_/B _161_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_14 vgnd vpwr scs8hd_decap_12
XFILLER_1_58 vgnd vpwr scs8hd_decap_3
XANTENNA__136__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_130 vpwr vgnd scs8hd_fill_2
XFILLER_28_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XFILLER_19_21 vpwr vgnd scs8hd_fill_2
XFILLER_42_122 vpwr vgnd scs8hd_fill_2
XFILLER_35_97 vgnd vpwr scs8hd_decap_3
XFILLER_35_86 vpwr vgnd scs8hd_fill_2
XFILLER_35_75 vpwr vgnd scs8hd_fill_2
XFILLER_35_53 vpwr vgnd scs8hd_fill_2
XFILLER_35_20 vgnd vpwr scs8hd_decap_6
XFILLER_27_130 vgnd vpwr scs8hd_decap_4
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
X_144_ _129_/X _143_/X _144_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XFILLER_18_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_111 vgnd vpwr scs8hd_decap_6
XFILLER_24_199 vgnd vpwr scs8hd_decap_12
XFILLER_21_77 vgnd vpwr scs8hd_fill_1
XPHY_8 vgnd vpwr scs8hd_decap_3
X_127_ _096_/X _127_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__133__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_16_11 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XFILLER_16_44 vgnd vpwr scs8hd_decap_3
XFILLER_8_129 vgnd vpwr scs8hd_decap_12
XANTENNA__234__A _234_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_206 vgnd vpwr scs8hd_decap_12
XANTENNA__144__A _129_/X vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
XFILLER_26_206 vgnd vpwr scs8hd_decap_8
Xmux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _186_/A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XANTENNA__130__C _100_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _160_/C vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _204_/A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_31_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_34 vpwr vgnd scs8hd_fill_2
XFILLER_38_64 vgnd vpwr scs8hd_decap_3
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
Xmem_left_track_3.LATCH_0_.latch data_in _193_/A _148_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__141__B _140_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_10 vgnd vpwr scs8hd_fill_1
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
X_160_ _122_/A _113_/Y _160_/C _160_/D _162_/B vgnd vpwr scs8hd_or4_4
XANTENNA__242__A _242_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_26 vgnd vpwr scs8hd_decap_12
XANTENNA__136__B _135_/B vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _096_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_10.LATCH_1_.latch data_in _182_/A _127_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_27_120 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_fill_1
XANTENNA__237__A _237_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_65 vgnd vpwr scs8hd_decap_4
XFILLER_35_32 vgnd vpwr scs8hd_decap_4
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
XFILLER_27_164 vpwr vgnd scs8hd_fill_2
XFILLER_27_175 vpwr vgnd scs8hd_fill_2
XFILLER_27_197 vgnd vpwr scs8hd_decap_4
X_143_ _104_/A _123_/B _157_/C _157_/D _143_/X vgnd vpwr scs8hd_or4_4
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XANTENNA__147__A _129_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_145 vgnd vpwr scs8hd_decap_3
XFILLER_21_34 vgnd vpwr scs8hd_decap_8
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
X_126_ _123_/A _123_/B _123_/C _171_/A _127_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_21_148 vpwr vgnd scs8hd_fill_2
XFILLER_29_204 vgnd vpwr scs8hd_decap_12
XFILLER_16_89 vgnd vpwr scs8hd_fill_1
XFILLER_32_88 vgnd vpwr scs8hd_fill_1
XFILLER_35_218 vpwr vgnd scs8hd_fill_2
XANTENNA__144__B _143_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
XANTENNA__160__A _122_/A vgnd vpwr scs8hd_diode_2
X_109_ _157_/D _171_/A vgnd vpwr scs8hd_buf_1
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_77 vgnd vpwr scs8hd_decap_3
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XANTENNA__130__D _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_6 vgnd vpwr scs8hd_decap_12
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_38_98 vgnd vpwr scs8hd_decap_3
XFILLER_13_232 vgnd vpwr scs8hd_decap_12
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_39_184 vgnd vpwr scs8hd_fill_1
XFILLER_24_23 vgnd vpwr scs8hd_decap_8
XFILLER_24_56 vpwr vgnd scs8hd_fill_2
XFILLER_10_202 vgnd vpwr scs8hd_decap_12
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _189_/A mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_1_38 vgnd vpwr scs8hd_decap_12
XFILLER_39_3 vpwr vgnd scs8hd_fill_2
XFILLER_36_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _207_/A mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_19_34 vpwr vgnd scs8hd_fill_2
XFILLER_19_78 vpwr vgnd scs8hd_fill_2
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
X_142_ _133_/A _140_/X _142_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_15.tap_buf4_0_.scs8hd_inv_1 mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _227_/A vgnd vpwr scs8hd_inv_1
XFILLER_33_179 vpwr vgnd scs8hd_fill_2
XANTENNA__147__B _146_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_143 vgnd vpwr scs8hd_decap_8
XFILLER_18_154 vgnd vpwr scs8hd_decap_12
XANTENNA__163__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_190 vpwr vgnd scs8hd_fill_2
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_13 vpwr vgnd scs8hd_fill_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_135 vgnd vpwr scs8hd_decap_12
X_125_ _117_/A _124_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_30_7 vpwr vgnd scs8hd_fill_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_14_190 vgnd vpwr scs8hd_decap_12
XFILLER_21_138 vpwr vgnd scs8hd_fill_2
XANTENNA__158__A _164_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_216 vgnd vpwr scs8hd_decap_12
XFILLER_16_68 vpwr vgnd scs8hd_fill_2
XFILLER_32_45 vgnd vpwr scs8hd_decap_3
XFILLER_32_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_12 vpwr vgnd scs8hd_fill_2
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.tap_buf4_0_.scs8hd_inv_1 mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _231_/A vgnd vpwr scs8hd_inv_1
XFILLER_11_171 vgnd vpwr scs8hd_decap_12
X_108_ address[1] enable _157_/D vgnd vpwr scs8hd_nand2_4
XFILLER_21_3 vgnd vpwr scs8hd_fill_1
XANTENNA__160__B _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
XFILLER_8_80 vgnd vpwr scs8hd_decap_12
XFILLER_17_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_12 vpwr vgnd scs8hd_fill_2
XFILLER_27_34 vpwr vgnd scs8hd_fill_2
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_255 vgnd vpwr scs8hd_decap_12
XFILLER_31_200 vgnd vpwr scs8hd_fill_1
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XANTENNA__171__A _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_211 vgnd vpwr scs8hd_decap_3
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_44 vgnd vpwr scs8hd_decap_4
XFILLER_38_22 vgnd vpwr scs8hd_decap_8
XANTENNA__166__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _183_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _179_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_111 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_13 vpwr vgnd scs8hd_fill_2
XFILLER_42_125 vgnd vpwr scs8hd_decap_3
XFILLER_42_114 vgnd vpwr scs8hd_decap_8
XFILLER_42_103 vgnd vpwr scs8hd_decap_8
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
X_141_ _129_/X _140_/X _141_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _180_/A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_158 vgnd vpwr scs8hd_decap_6
XFILLER_33_136 vpwr vgnd scs8hd_fill_2
XFILLER_33_114 vpwr vgnd scs8hd_fill_2
XFILLER_33_103 vgnd vpwr scs8hd_decap_6
XFILLER_18_166 vgnd vpwr scs8hd_decap_12
XFILLER_41_191 vpwr vgnd scs8hd_fill_2
XANTENNA__163__B _113_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_117 vgnd vpwr scs8hd_decap_4
XFILLER_30_106 vpwr vgnd scs8hd_fill_2
XFILLER_15_147 vgnd vpwr scs8hd_decap_12
X_124_ _096_/X _124_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_139 vgnd vpwr scs8hd_decap_4
XFILLER_23_180 vgnd vpwr scs8hd_decap_3
XFILLER_11_91 vgnd vpwr scs8hd_decap_12
XFILLER_23_7 vgnd vpwr scs8hd_decap_3
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _157_/X vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_228 vgnd vpwr scs8hd_decap_12
XFILLER_12_117 vgnd vpwr scs8hd_decap_12
XFILLER_16_25 vgnd vpwr scs8hd_fill_1
XFILLER_32_68 vgnd vpwr scs8hd_decap_4
X_107_ _117_/A _107_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_110 vgnd vpwr scs8hd_decap_12
XANTENNA__160__C _160_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _185_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__169__A _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XFILLER_25_231 vgnd vpwr scs8hd_decap_12
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_267 vgnd vpwr scs8hd_decap_8
XFILLER_31_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _181_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__171__B _169_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _184_/A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XANTENNA__166__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__182__A _182_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _202_/A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XFILLER_24_36 vpwr vgnd scs8hd_fill_2
XFILLER_40_46 vgnd vpwr scs8hd_decap_3
XFILLER_40_24 vgnd vpwr scs8hd_decap_6
XFILLER_14_91 vgnd vpwr scs8hd_fill_1
Xmux_left_track_13.INVTX1_0_.scs8hd_inv_1 chany_top_in[3] mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_8
XFILLER_36_167 vgnd vpwr scs8hd_decap_8
XFILLER_36_145 vpwr vgnd scs8hd_fill_2
XFILLER_36_134 vpwr vgnd scs8hd_fill_2
XFILLER_36_189 vgnd vpwr scs8hd_decap_8
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_35_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_112 vpwr vgnd scs8hd_fill_2
X_140_ _104_/A _123_/B _157_/C _160_/D _140_/X vgnd vpwr scs8hd_or4_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _221_/HI _188_/Y mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_123 vgnd vpwr scs8hd_decap_4
XFILLER_18_134 vgnd vpwr scs8hd_decap_3
XFILLER_41_170 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_178 vgnd vpwr scs8hd_decap_12
XANTENNA__163__C _160_/C vgnd vpwr scs8hd_diode_2
Xmem_top_track_6.LATCH_0_.latch data_in _179_/A _120_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _206_/Y mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_104 vpwr vgnd scs8hd_fill_2
XFILLER_15_159 vgnd vpwr scs8hd_decap_12
X_123_ _123_/A _123_/B _123_/C _169_/A _124_/B vgnd vpwr scs8hd_or4_4
XFILLER_11_70 vgnd vpwr scs8hd_decap_3
XFILLER_16_7 vgnd vpwr scs8hd_decap_4
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_129 vgnd vpwr scs8hd_decap_12
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
X_106_ address[0] _117_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
XFILLER_22_91 vgnd vpwr scs8hd_fill_1
XANTENNA__160__D _160_/D vgnd vpwr scs8hd_diode_2
XANTENNA__169__B _169_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XFILLER_25_243 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_4_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__171__C _165_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XANTENNA__166__C address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_143 vpwr vgnd scs8hd_fill_2
XFILLER_39_121 vgnd vpwr scs8hd_fill_1
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XFILLER_40_58 vgnd vpwr scs8hd_decap_12
XFILLER_6_6 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
Xmem_left_track_7.LATCH_1_.latch data_in _196_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_168 vpwr vgnd scs8hd_fill_2
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_90 vgnd vpwr scs8hd_decap_4
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__163__D _157_/D vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _187_/A mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_3
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_11.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__098__A address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_171 vgnd vpwr scs8hd_decap_6
X_122_ _122_/A _123_/A vgnd vpwr scs8hd_buf_1
Xmux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _205_/A mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_241 vgnd vpwr scs8hd_decap_3
XFILLER_16_49 vgnd vpwr scs8hd_decap_12
XFILLER_20_130 vgnd vpwr scs8hd_decap_4
XFILLER_20_163 vgnd vpwr scs8hd_decap_12
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
X_105_ _096_/X _107_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
XFILLER_22_70 vpwr vgnd scs8hd_fill_2
XFILLER_34_200 vgnd vpwr scs8hd_decap_12
XANTENNA__169__C _165_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_17 vpwr vgnd scs8hd_fill_2
XFILLER_13_28 vgnd vpwr scs8hd_decap_4
XFILLER_13_39 vpwr vgnd scs8hd_fill_2
XFILLER_38_69 vgnd vpwr scs8hd_decap_4
XFILLER_38_36 vgnd vpwr scs8hd_decap_6
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XANTENNA__166__D _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_10_18 vgnd vpwr scs8hd_decap_12
XFILLER_19_38 vpwr vgnd scs8hd_fill_2
XFILLER_27_147 vpwr vgnd scs8hd_fill_2
XFILLER_35_191 vpwr vgnd scs8hd_fill_2
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_92 vpwr vgnd scs8hd_fill_2
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
XFILLER_24_128 vpwr vgnd scs8hd_fill_2
XFILLER_32_194 vgnd vpwr scs8hd_decap_4
XFILLER_21_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_19 vgnd vpwr scs8hd_decap_12
X_121_ address[3] _122_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _208_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _178_/A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_28 vgnd vpwr scs8hd_decap_3
XFILLER_32_27 vpwr vgnd scs8hd_fill_2
XFILLER_32_16 vgnd vpwr scs8hd_decap_4
XFILLER_20_175 vgnd vpwr scs8hd_decap_12
Xmem_top_track_2.LATCH_0_.latch data_in _175_/A _112_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
Xmem_left_track_17.LATCH_0_.latch data_in _207_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_104_ _104_/A _123_/B _123_/C _169_/A _107_/B vgnd vpwr scs8hd_or4_4
XFILLER_34_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_6 vpwr vgnd scs8hd_fill_2
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_27_16 vpwr vgnd scs8hd_fill_2
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_245 vgnd vpwr scs8hd_decap_12
XFILLER_27_38 vpwr vgnd scs8hd_fill_2
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_204 vpwr vgnd scs8hd_fill_2
XFILLER_17_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_81 vgnd vpwr scs8hd_decap_3
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_38_59 vgnd vpwr scs8hd_decap_3
XFILLER_9_208 vgnd vpwr scs8hd_decap_12
XFILLER_28_81 vpwr vgnd scs8hd_fill_2
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_39_189 vpwr vgnd scs8hd_fill_2
XFILLER_39_156 vpwr vgnd scs8hd_fill_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_4
XFILLER_39_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_83 vgnd vpwr scs8hd_decap_8
Xmux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _182_/A mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_71 vpwr vgnd scs8hd_fill_2
XFILLER_39_80 vpwr vgnd scs8hd_fill_2
XFILLER_19_17 vpwr vgnd scs8hd_fill_2
XFILLER_35_38 vpwr vgnd scs8hd_fill_2
XFILLER_27_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _220_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _200_/A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_25_71 vpwr vgnd scs8hd_fill_2
XFILLER_26_181 vgnd vpwr scs8hd_decap_4
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_41_151 vgnd vpwr scs8hd_decap_6
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _184_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _235_/A vgnd vpwr scs8hd_inv_1
XFILLER_24_107 vpwr vgnd scs8hd_fill_2
XFILLER_32_173 vpwr vgnd scs8hd_fill_2
XFILLER_17_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_3.LATCH_1_.latch data_in _192_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_120_ _117_/A _120_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
XFILLER_11_62 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _220_/HI _186_/Y mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_221 vgnd vpwr scs8hd_decap_12
XFILLER_20_110 vgnd vpwr scs8hd_decap_6
XFILLER_20_187 vgnd vpwr scs8hd_decap_12
XFILLER_11_121 vgnd vpwr scs8hd_fill_1
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_7_147 vgnd vpwr scs8hd_decap_12
X_103_ _160_/D _169_/A vgnd vpwr scs8hd_buf_1
XFILLER_22_50 vgnd vpwr scs8hd_decap_4
XFILLER_22_83 vpwr vgnd scs8hd_fill_2
Xmux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _204_/Y mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_30 vgnd vpwr scs8hd_fill_1
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_72 vgnd vpwr scs8hd_fill_1
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _181_/A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_28_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_5_31 vgnd vpwr scs8hd_decap_12
XFILLER_39_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_36_149 vgnd vpwr scs8hd_decap_4
XFILLER_36_138 vgnd vpwr scs8hd_decap_4
XANTENNA__101__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_116 vpwr vgnd scs8hd_fill_2
XFILLER_4_6 vgnd vpwr scs8hd_decap_12
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_41_71 vpwr vgnd scs8hd_fill_2
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_15_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_15_108 vgnd vpwr scs8hd_decap_12
XFILLER_23_196 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vgnd vpwr scs8hd_decap_4
XFILLER_14_141 vgnd vpwr scs8hd_decap_12
X_179_ _179_/A _179_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_233 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_3 vpwr vgnd scs8hd_fill_2
XFILLER_20_199 vgnd vpwr scs8hd_decap_12
Xmux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _185_/A mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_159 vgnd vpwr scs8hd_decap_12
X_102_ address[1] _101_/Y _160_/D vgnd vpwr scs8hd_or2_4
Xmux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _203_/A mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_27_29 vgnd vpwr scs8hd_decap_3
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_17_62 vgnd vpwr scs8hd_decap_3
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_13.LATCH_0_.latch data_in _203_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _189_/Y mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_28_61 vgnd vpwr scs8hd_fill_1
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_114 vgnd vpwr scs8hd_decap_4
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_5_43 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_11.tap_buf4_0_.scs8hd_inv_1 mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _207_/Y mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_30_62 vpwr vgnd scs8hd_fill_2
XFILLER_30_84 vgnd vpwr scs8hd_decap_4
XFILLER_39_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_left_in[5] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_106 vpwr vgnd scs8hd_fill_2
XFILLER_18_139 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XFILLER_41_175 vgnd vpwr scs8hd_decap_8
XFILLER_41_164 vgnd vpwr scs8hd_decap_4
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_26_161 vgnd vpwr scs8hd_decap_6
XFILLER_26_194 vgnd vpwr scs8hd_decap_12
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__112__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XFILLER_32_131 vgnd vpwr scs8hd_decap_3
Xmux_left_track_3.tap_buf4_0_.scs8hd_inv_1 mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _233_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in _189_/A _142_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_142 vgnd vpwr scs8hd_fill_1
XFILLER_11_75 vpwr vgnd scs8hd_fill_2
XFILLER_36_61 vgnd vpwr scs8hd_fill_1
Xmux_top_track_4.tap_buf4_0_.scs8hd_inv_1 mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _241_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__107__A _117_/A vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_13_ mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_145 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
X_101_ enable _101_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_41 vgnd vpwr scs8hd_decap_3
XFILLER_22_96 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _176_/A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XFILLER_17_52 vpwr vgnd scs8hd_fill_2
XFILLER_17_85 vpwr vgnd scs8hd_fill_2
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_73 vpwr vgnd scs8hd_fill_2
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__104__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vpwr vgnd scs8hd_fill_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _198_/A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_38_18 vpwr vgnd scs8hd_fill_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_28_51 vpwr vgnd scs8hd_fill_2
XFILLER_12_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_55 vgnd vpwr scs8hd_decap_6
XANTENNA__115__A _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _185_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _225_/HI _180_/Y mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
XFILLER_30_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_162 vpwr vgnd scs8hd_fill_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _181_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_198 vpwr vgnd scs8hd_fill_2
XFILLER_41_187 vpwr vgnd scs8hd_fill_2
XFILLER_41_143 vpwr vgnd scs8hd_fill_2
XFILLER_41_132 vpwr vgnd scs8hd_fill_2
XFILLER_41_40 vpwr vgnd scs8hd_fill_2
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_25_41 vgnd vpwr scs8hd_decap_3
XFILLER_25_96 vpwr vgnd scs8hd_fill_2
XPHY_52 vgnd vpwr scs8hd_decap_3
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__112__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_154 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
XFILLER_23_110 vpwr vgnd scs8hd_fill_2
XFILLER_23_132 vgnd vpwr scs8hd_decap_4
XFILLER_23_154 vpwr vgnd scs8hd_fill_2
XFILLER_11_21 vpwr vgnd scs8hd_fill_2
XFILLER_11_10 vpwr vgnd scs8hd_fill_2
XFILLER_36_84 vpwr vgnd scs8hd_fill_2
XFILLER_36_51 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd vpwr
+ scs8hd_diode_2
X_177_ _177_/A _177_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__107__B _107_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_6 vgnd vpwr scs8hd_decap_8
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_6.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_37_202 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XFILLER_28_213 vgnd vpwr scs8hd_fill_1
XFILLER_11_135 vgnd vpwr scs8hd_decap_12
X_100_ _100_/A _123_/C vgnd vpwr scs8hd_buf_1
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _104_/A vgnd vpwr scs8hd_diode_2
X_229_ _229_/A chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_10_190 vgnd vpwr scs8hd_decap_12
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_40_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _219_/HI _184_/Y mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _187_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_12.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_75 vgnd vpwr scs8hd_fill_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_6.LATCH_1_.latch data_in _178_/A _119_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__104__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _202_/Y mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_28_85 vgnd vpwr scs8hd_decap_4
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XANTENNA__115__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_127 vgnd vpwr scs8hd_fill_1
XANTENNA__131__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_10 vgnd vpwr scs8hd_decap_4
XFILLER_39_62 vgnd vpwr scs8hd_decap_3
XFILLER_39_51 vpwr vgnd scs8hd_fill_2
XFILLER_29_193 vpwr vgnd scs8hd_fill_2
Xmux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _179_/A mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _221_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_18_119 vpwr vgnd scs8hd_fill_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XFILLER_25_75 vpwr vgnd scs8hd_fill_2
XFILLER_41_96 vgnd vpwr scs8hd_decap_6
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_177 vpwr vgnd scs8hd_fill_2
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _173_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_177 vgnd vpwr scs8hd_fill_1
XFILLER_2_6 vgnd vpwr scs8hd_decap_12
XFILLER_14_166 vgnd vpwr scs8hd_decap_12
X_176_ _176_/A _176_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_103 vgnd vpwr scs8hd_decap_12
XFILLER_11_147 vgnd vpwr scs8hd_decap_12
XFILLER_22_21 vpwr vgnd scs8hd_fill_2
XFILLER_22_54 vgnd vpwr scs8hd_fill_1
XFILLER_22_87 vpwr vgnd scs8hd_fill_2
Xmem_top_track_12.LATCH_0_.latch data_in _185_/A _133_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_269 vgnd vpwr scs8hd_decap_8
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _115_/B vgnd vpwr scs8hd_diode_2
X_228_ _228_/A chanx_left_out[6] vgnd vpwr scs8hd_buf_2
X_159_ _165_/A _157_/X _159_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.INVTX1_1_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _183_/A mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_33_86 vpwr vgnd scs8hd_fill_2
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XFILLER_33_20 vpwr vgnd scs8hd_fill_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
XANTENNA__104__D _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA__129__A _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
Xmux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _201_/A mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_28_64 vgnd vpwr scs8hd_decap_4
XFILLER_28_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_202 vgnd vpwr scs8hd_decap_12
XANTENNA__115__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA__131__B _133_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_10.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_9_ mux_top_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__232__A _232_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _187_/Y mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__126__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_175 vpwr vgnd scs8hd_fill_2
XANTENNA__227__A _227_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_26_131 vgnd vpwr scs8hd_decap_3
XFILLER_41_75 vgnd vpwr scs8hd_decap_4
XFILLER_41_53 vgnd vpwr scs8hd_decap_6
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _205_/Y mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_32_145 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_97 vgnd vpwr scs8hd_fill_1
XFILLER_14_178 vgnd vpwr scs8hd_decap_12
X_175_ _175_/A _175_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_126 vpwr vgnd scs8hd_fill_2
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XFILLER_11_115 vgnd vpwr scs8hd_decap_6
XFILLER_11_159 vgnd vpwr scs8hd_decap_12
XFILLER_22_66 vpwr vgnd scs8hd_fill_2
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
X_227_ _227_/A chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
XANTENNA__118__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
X_158_ _164_/A _157_/X _158_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA__150__A _129_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_3
XFILLER_25_207 vgnd vpwr scs8hd_decap_12
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__235__A _235_/A vgnd vpwr scs8hd_diode_2
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_32 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_12
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _205_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_28_32 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.INVTX1_1_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _174_/A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__115__D _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_118 vgnd vpwr scs8hd_fill_1
XFILLER_10_6 vgnd vpwr scs8hd_decap_12
Xmem_top_track_2.LATCH_1_.latch data_in _174_/A _111_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_17.LATCH_1_.latch data_in _206_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _196_/A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_67 vgnd vpwr scs8hd_decap_3
XFILLER_30_11 vpwr vgnd scs8hd_fill_2
XFILLER_30_22 vpwr vgnd scs8hd_fill_2
XFILLER_30_66 vgnd vpwr scs8hd_decap_3
XFILLER_30_88 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_97 vpwr vgnd scs8hd_fill_2
XFILLER_29_140 vgnd vpwr scs8hd_fill_1
XFILLER_29_173 vpwr vgnd scs8hd_fill_2
XANTENNA__142__B _140_/X vgnd vpwr scs8hd_diode_2
XANTENNA__126__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_198 vpwr vgnd scs8hd_fill_2
XFILLER_35_187 vpwr vgnd scs8hd_fill_2
XFILLER_35_143 vpwr vgnd scs8hd_fill_2
XFILLER_35_121 vgnd vpwr scs8hd_fill_1
XFILLER_26_110 vpwr vgnd scs8hd_fill_2
XFILLER_41_102 vgnd vpwr scs8hd_fill_1
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_25_33 vpwr vgnd scs8hd_fill_2
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_41_21 vgnd vpwr scs8hd_decap_4
XANTENNA__243__A _243_/A vgnd vpwr scs8hd_diode_2
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_32_102 vgnd vpwr scs8hd_decap_12
XFILLER_17_121 vgnd vpwr scs8hd_fill_1
XFILLER_32_124 vgnd vpwr scs8hd_decap_4
Xmux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _224_/HI _178_/Y mux_top_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__153__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_79 vgnd vpwr scs8hd_decap_12
XFILLER_36_65 vgnd vpwr scs8hd_decap_8
XFILLER_36_32 vgnd vpwr scs8hd_decap_8
XANTENNA__238__A _238_/A vgnd vpwr scs8hd_diode_2
X_243_ _243_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd vpwr
+ scs8hd_diode_2
X_174_ _174_/A _174_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__D _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_7 vpwr vgnd scs8hd_fill_2
XANTENNA__148__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_116 vgnd vpwr scs8hd_fill_1
XFILLER_36_260 vgnd vpwr scs8hd_decap_12
XFILLER_28_205 vgnd vpwr scs8hd_decap_8
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _222_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
X_226_ _226_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_7_ mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_157_ _123_/A address[2] _157_/C _157_/D _157_/X vgnd vpwr scs8hd_or4_4
XANTENNA__134__C _100_/A vgnd vpwr scs8hd_diode_2
XANTENNA__118__D _171_/A vgnd vpwr scs8hd_diode_2
XANTENNA__150__B _149_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_fill_1
XFILLER_25_219 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _184_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_23 vgnd vpwr scs8hd_fill_1
XFILLER_17_56 vgnd vpwr scs8hd_decap_4
XFILLER_17_89 vpwr vgnd scs8hd_fill_2
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_99 vpwr vgnd scs8hd_fill_2
XFILLER_33_77 vpwr vgnd scs8hd_fill_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__145__B _143_/X vgnd vpwr scs8hd_diode_2
XANTENNA__161__A _164_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XFILLER_28_55 vgnd vpwr scs8hd_decap_6
XFILLER_28_77 vpwr vgnd scs8hd_fill_2
Xmux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _218_/HI _182_/Y mux_top_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XANTENNA__156__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_163 vpwr vgnd scs8hd_fill_2
XFILLER_14_35 vgnd vpwr scs8hd_decap_12
XFILLER_14_79 vpwr vgnd scs8hd_fill_2
XFILLER_30_45 vgnd vpwr scs8hd_decap_4
XFILLER_39_43 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_12.tap_buf4_0_.scs8hd_inv_1 mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _237_/A vgnd vpwr scs8hd_inv_1
XFILLER_39_76 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _209_/HI _200_/Y mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_152 vpwr vgnd scs8hd_fill_2
XANTENNA__126__D _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vpwr vgnd scs8hd_fill_2
XFILLER_41_136 vgnd vpwr scs8hd_decap_4
XFILLER_41_114 vpwr vgnd scs8hd_fill_2
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XFILLER_26_177 vpwr vgnd scs8hd_fill_2
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_32_114 vgnd vpwr scs8hd_fill_1
XFILLER_17_133 vgnd vpwr scs8hd_decap_12
XFILLER_40_191 vgnd vpwr scs8hd_decap_6
XANTENNA__153__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _177_/A mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_23_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _186_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_25 vgnd vpwr scs8hd_decap_12
XFILLER_36_88 vgnd vpwr scs8hd_decap_4
XFILLER_36_55 vgnd vpwr scs8hd_decap_6
X_173_ _173_/A _173_/Y vgnd vpwr scs8hd_inv_8
X_242_ _242_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _199_/A mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__148__B _146_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vpwr vgnd scs8hd_fill_2
XANTENNA__164__A _164_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_272 vgnd vpwr scs8hd_decap_3
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_22_46 vpwr vgnd scs8hd_fill_2
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
X_225_ _225_/HI _225_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
X_156_ _165_/A _153_/X _156_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__D _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_7 vgnd vpwr scs8hd_fill_1
XANTENNA__159__A _165_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_13 vpwr vgnd scs8hd_fill_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_35 vpwr vgnd scs8hd_fill_2
XFILLER_17_68 vgnd vpwr scs8hd_decap_4
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _181_/Y mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
X_139_ _160_/C _157_/C vgnd vpwr scs8hd_buf_1
XANTENNA__161__B _162_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_3 vgnd vpwr scs8hd_fill_1
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_5_ mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_23 vpwr vgnd scs8hd_fill_2
XFILLER_28_89 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _153_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _172_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_131 vgnd vpwr scs8hd_decap_4
XFILLER_14_47 vgnd vpwr scs8hd_decap_12
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XFILLER_39_55 vpwr vgnd scs8hd_fill_2
XFILLER_39_22 vpwr vgnd scs8hd_fill_2
XFILLER_29_197 vgnd vpwr scs8hd_decap_4
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XFILLER_35_123 vgnd vpwr scs8hd_decap_3
XANTENNA__167__A _166_/X vgnd vpwr scs8hd_diode_2
Xmem_left_track_13.LATCH_1_.latch data_in _202_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_26_145 vpwr vgnd scs8hd_fill_2
XFILLER_26_167 vgnd vpwr scs8hd_fill_1
XFILLER_41_159 vpwr vgnd scs8hd_fill_2
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_25_79 vpwr vgnd scs8hd_fill_2
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vpwr vgnd scs8hd_fill_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_4
XFILLER_17_145 vgnd vpwr scs8hd_decap_12
XANTENNA__153__C _157_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _185_/Y mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_11_37 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_172_ _172_/A _172_/Y vgnd vpwr scs8hd_inv_8
X_241_ _241_/A chany_top_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__164__B _164_/B vgnd vpwr scs8hd_diode_2
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_196 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _203_/Y mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_22_25 vgnd vpwr scs8hd_decap_6
Xmem_left_track_9.LATCH_0_.latch data_in _199_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_240 vgnd vpwr scs8hd_decap_4
X_224_ _224_/HI _224_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
X_155_ address[0] _165_/A vgnd vpwr scs8hd_buf_1
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
XFILLER_33_243 vgnd vpwr scs8hd_fill_1
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _157_/X vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_24 vpwr vgnd scs8hd_fill_2
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_1_.latch data_in _188_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_207_ _207_/A _207_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_213 vgnd vpwr scs8hd_fill_1
X_138_ address[4] _137_/Y _160_/C vgnd vpwr scs8hd_nand2_4
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_21_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XFILLER_12_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_110 vpwr vgnd scs8hd_fill_2
XFILLER_14_59 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_3_ mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_102 vgnd vpwr scs8hd_decap_3
XFILLER_35_179 vgnd vpwr scs8hd_decap_4
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _172_/A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _243_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_26_102 vpwr vgnd scs8hd_fill_2
XFILLER_26_157 vpwr vgnd scs8hd_fill_2
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_2_18 vgnd vpwr scs8hd_decap_12
XFILLER_17_102 vpwr vgnd scs8hd_fill_2
XFILLER_17_113 vpwr vgnd scs8hd_fill_2
XFILLER_40_171 vgnd vpwr scs8hd_decap_12
XFILLER_32_149 vgnd vpwr scs8hd_decap_4
XFILLER_17_157 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _194_/A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__153__D _160_/D vgnd vpwr scs8hd_diode_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_138 vgnd vpwr scs8hd_decap_4
XFILLER_31_193 vgnd vpwr scs8hd_decap_4
XFILLER_16_190 vgnd vpwr scs8hd_decap_12
XFILLER_11_49 vgnd vpwr scs8hd_decap_12
X_240_ _240_/A chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
X_171_ _171_/A _169_/B _165_/A _171_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_13_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _223_/HI _176_/Y mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
X_223_ _223_/HI _223_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_141 vgnd vpwr scs8hd_decap_12
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
X_154_ _164_/A _153_/X _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _216_/HI _198_/Y mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_211 vgnd vpwr scs8hd_decap_3
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_36 vpwr vgnd scs8hd_fill_2
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
X_206_ _206_/A _206_/Y vgnd vpwr scs8hd_inv_8
X_137_ address[5] _137_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XFILLER_28_36 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_26 vgnd vpwr scs8hd_decap_4
XFILLER_29_177 vgnd vpwr scs8hd_decap_4
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_158 vpwr vgnd scs8hd_fill_2
XFILLER_35_114 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _187_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _230_/A vgnd vpwr scs8hd_inv_1
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vpwr vgnd scs8hd_fill_2
XFILLER_25_37 vpwr vgnd scs8hd_fill_2
XFILLER_26_114 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_41_36 vpwr vgnd scs8hd_fill_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_17_169 vgnd vpwr scs8hd_decap_12
XFILLER_40_183 vgnd vpwr scs8hd_decap_4
XFILLER_32_128 vgnd vpwr scs8hd_fill_1
XFILLER_15_70 vgnd vpwr scs8hd_fill_1
XFILLER_25_191 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_1_ mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_17 vpwr vgnd scs8hd_fill_2
XFILLER_39_261 vpwr vgnd scs8hd_fill_2
X_170_ _171_/A _169_/B _164_/A _170_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_14_117 vgnd vpwr scs8hd_decap_12
XFILLER_37_209 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_110 vgnd vpwr scs8hd_decap_12
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _223_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_42_201 vgnd vpwr scs8hd_decap_12
Xmux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _175_/A mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_222_ _222_/HI _222_/LO vgnd vpwr scs8hd_conb_1
XFILLER_8_18 vgnd vpwr scs8hd_decap_12
X_153_ _123_/A address[2] _157_/C _160_/D _153_/X vgnd vpwr scs8hd_or4_4
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
XFILLER_26_8 vgnd vpwr scs8hd_fill_1
XFILLER_37_90 vpwr vgnd scs8hd_fill_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _197_/A mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _173_/Y vgnd vpwr
+ scs8hd_diode_2
X_205_ _205_/A _205_/Y vgnd vpwr scs8hd_inv_8
Xmem_left_track_5.LATCH_0_.latch data_in _195_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd vpwr
+ scs8hd_diode_2
X_136_ _133_/A _135_/B _136_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_19 vgnd vpwr scs8hd_decap_12
Xmux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _179_/Y mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_119_ _096_/X _120_/B _119_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_12.LATCH_1_.latch data_in _184_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_145 vpwr vgnd scs8hd_fill_2
XFILLER_38_189 vgnd vpwr scs8hd_decap_8
XFILLER_38_178 vgnd vpwr scs8hd_decap_8
XFILLER_38_167 vgnd vpwr scs8hd_decap_8
XFILLER_14_17 vgnd vpwr scs8hd_decap_12
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_14 vpwr vgnd scs8hd_fill_2
XFILLER_29_156 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_118 vpwr vgnd scs8hd_fill_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
XFILLER_15_82 vpwr vgnd scs8hd_fill_2
XFILLER_15_93 vpwr vgnd scs8hd_fill_2
XFILLER_25_170 vpwr vgnd scs8hd_fill_2
XFILLER_31_140 vpwr vgnd scs8hd_fill_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_36_15 vpwr vgnd scs8hd_fill_2
XFILLER_14_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _175_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_74 vgnd vpwr scs8hd_decap_12
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_42_213 vgnd vpwr scs8hd_decap_4
Xmux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _183_/Y mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_154 vgnd vpwr scs8hd_decap_12
X_221_ _221_/HI _221_/LO vgnd vpwr scs8hd_conb_1
X_152_ _096_/A _164_/A vgnd vpwr scs8hd_buf_1
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_17 vgnd vpwr scs8hd_decap_6
XFILLER_17_39 vpwr vgnd scs8hd_fill_2
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _201_/Y mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_71 vpwr vgnd scs8hd_fill_2
X_135_ _129_/X _135_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_6 vpwr vgnd scs8hd_fill_2
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_227 vgnd vpwr scs8hd_decap_12
XFILLER_7_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
X_118_ _104_/A _115_/B _123_/C _171_/A _120_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_135 vgnd vpwr scs8hd_fill_1
XFILLER_22_3 vpwr vgnd scs8hd_fill_2
XFILLER_14_29 vpwr vgnd scs8hd_fill_2
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_39_26 vpwr vgnd scs8hd_fill_2
XFILLER_29_113 vgnd vpwr scs8hd_decap_3
XFILLER_20_72 vgnd vpwr scs8hd_fill_1
XFILLER_29_92 vpwr vgnd scs8hd_fill_2
XFILLER_6_30 vgnd vpwr scs8hd_fill_1
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_26_127 vpwr vgnd scs8hd_fill_2
XFILLER_26_149 vgnd vpwr scs8hd_decap_4
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_9_7 vgnd vpwr scs8hd_decap_12
XFILLER_25_182 vgnd vpwr scs8hd_fill_1
XFILLER_40_163 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _205_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_130 vpwr vgnd scs8hd_fill_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_42_81 vgnd vpwr scs8hd_decap_12
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_86 vgnd vpwr scs8hd_decap_12
XFILLER_3_31 vgnd vpwr scs8hd_decap_12
XFILLER_36_200 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _192_/A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
X_220_ _220_/HI _220_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_166 vgnd vpwr scs8hd_decap_12
X_151_ _133_/A _149_/X _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _222_/HI _174_/Y mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
X_134_ _123_/A _115_/B _100_/A _171_/A _135_/B vgnd vpwr scs8hd_or4_4
XFILLER_0_10 vgnd vpwr scs8hd_decap_4
XFILLER_0_21 vgnd vpwr scs8hd_decap_8
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _215_/HI _196_/Y mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_239 vgnd vpwr scs8hd_decap_12
X_117_ _117_/A _117_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _207_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_114 vgnd vpwr scs8hd_decap_4
Xmem_left_track_1.LATCH_0_.latch data_in _191_/A _145_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_136 vgnd vpwr scs8hd_decap_4
XFILLER_37_191 vpwr vgnd scs8hd_fill_2
XFILLER_29_169 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XFILLER_20_51 vpwr vgnd scs8hd_fill_2
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XFILLER_29_71 vgnd vpwr scs8hd_decap_4
XFILLER_35_139 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_19_180 vgnd vpwr scs8hd_decap_3
XFILLER_26_106 vpwr vgnd scs8hd_fill_2
XFILLER_41_17 vpwr vgnd scs8hd_fill_2
XFILLER_34_183 vpwr vgnd scs8hd_fill_2
XFILLER_17_106 vpwr vgnd scs8hd_fill_2
XFILLER_17_117 vpwr vgnd scs8hd_fill_2
XFILLER_15_40 vpwr vgnd scs8hd_fill_2
XFILLER_15_51 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_31_197 vgnd vpwr scs8hd_fill_1
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XFILLER_31_164 vpwr vgnd scs8hd_fill_2
XFILLER_39_253 vgnd vpwr scs8hd_decap_4
XFILLER_22_164 vpwr vgnd scs8hd_fill_2
XFILLER_22_175 vgnd vpwr scs8hd_decap_12
XFILLER_42_71 vgnd vpwr scs8hd_fill_1
XFILLER_9_135 vgnd vpwr scs8hd_decap_12
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_3_43 vgnd vpwr scs8hd_decap_12
XFILLER_36_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_190 vgnd vpwr scs8hd_decap_12
XFILLER_27_201 vgnd vpwr scs8hd_fill_1
XFILLER_27_245 vgnd vpwr scs8hd_decap_12
X_150_ _129_/X _149_/X _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_178 vgnd vpwr scs8hd_decap_12
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_37_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_215 vgnd vpwr scs8hd_decap_12
XFILLER_33_204 vgnd vpwr scs8hd_decap_8
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
X_133_ _133_/A _133_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _186_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__110__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _173_/A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_9_31 vgnd vpwr scs8hd_decap_12
XFILLER_9_86 vgnd vpwr scs8hd_decap_12
XFILLER_28_18 vgnd vpwr scs8hd_decap_3
XFILLER_20_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _195_/A mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_62 vgnd vpwr scs8hd_decap_3
XFILLER_34_61 vpwr vgnd scs8hd_fill_2
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
X_116_ _096_/X _117_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_39 vpwr vgnd scs8hd_fill_2
XFILLER_20_30 vgnd vpwr scs8hd_fill_1
XFILLER_35_118 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _177_/Y mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_25_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in _181_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_129 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_fill_1
XFILLER_40_132 vgnd vpwr scs8hd_decap_4
XFILLER_25_140 vpwr vgnd scs8hd_fill_2
XFILLER_25_195 vgnd vpwr scs8hd_decap_12
XANTENNA__102__B _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_261 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _199_/Y mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_121 vgnd vpwr scs8hd_fill_1
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_265 vgnd vpwr scs8hd_decap_12
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_22_121 vpwr vgnd scs8hd_fill_2
XFILLER_22_154 vgnd vpwr scs8hd_fill_1
XFILLER_22_187 vgnd vpwr scs8hd_decap_12
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _172_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_62 vpwr vgnd scs8hd_fill_2
XFILLER_42_61 vgnd vpwr scs8hd_fill_1
XFILLER_9_147 vgnd vpwr scs8hd_decap_12
XANTENNA__113__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_36_224 vgnd vpwr scs8hd_decap_8
XFILLER_3_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _224_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_3 vpwr vgnd scs8hd_fill_2
XFILLER_12_64 vgnd vpwr scs8hd_decap_3
XFILLER_18_202 vgnd vpwr scs8hd_decap_12
XFILLER_37_94 vpwr vgnd scs8hd_fill_2
XFILLER_33_227 vgnd vpwr scs8hd_decap_12
XANTENNA__108__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vpwr vgnd scs8hd_fill_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
X_132_ address[0] _133_/A vgnd vpwr scs8hd_buf_1
XFILLER_23_96 vgnd vpwr scs8hd_decap_3
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XANTENNA__110__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_43 vgnd vpwr scs8hd_decap_12
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
XFILLER_9_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_263 vgnd vpwr scs8hd_decap_12
XFILLER_34_84 vgnd vpwr scs8hd_decap_6
XANTENNA__105__B _107_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
X_115_ _104_/A _115_/B _123_/C _169_/A _117_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_127 vpwr vgnd scs8hd_fill_2
XANTENNA__121__A address[3] vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in _198_/A _158_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_149 vgnd vpwr scs8hd_decap_4
XFILLER_39_18 vpwr vgnd scs8hd_fill_2
XFILLER_37_160 vgnd vpwr scs8hd_decap_3
XFILLER_37_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_20_64 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_20_3 vpwr vgnd scs8hd_fill_2
XFILLER_34_163 vgnd vpwr scs8hd_decap_3
XFILLER_15_86 vgnd vpwr scs8hd_decap_4
XFILLER_15_97 vpwr vgnd scs8hd_fill_2
XFILLER_25_163 vgnd vpwr scs8hd_decap_4
XFILLER_25_174 vpwr vgnd scs8hd_fill_2
XFILLER_31_85 vpwr vgnd scs8hd_fill_2
XFILLER_31_52 vpwr vgnd scs8hd_fill_2
XFILLER_31_30 vpwr vgnd scs8hd_fill_2
XFILLER_0_273 vgnd vpwr scs8hd_decap_4
XFILLER_16_152 vgnd vpwr scs8hd_fill_1
XFILLER_31_144 vgnd vpwr scs8hd_decap_3
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

