magic
tech sky130A
magscale 1 2
timestamp 1606226223
<< locali >>
rect 17785 17051 17819 17221
rect 16773 15963 16807 16133
rect 15025 15351 15059 15657
rect 16221 15351 16255 15453
rect 16221 14807 16255 15113
rect 13553 13787 13587 14025
rect 13185 10047 13219 10149
rect 14473 9367 14507 9469
rect 14013 5151 14047 5321
rect 11437 3451 11471 3621
rect 6561 2839 6595 3077
rect 10517 3043 10551 3145
<< viali >>
rect 9045 20009 9079 20043
rect 11897 20009 11931 20043
rect 12817 20009 12851 20043
rect 13369 20009 13403 20043
rect 14565 20009 14599 20043
rect 15761 20009 15795 20043
rect 16865 20009 16899 20043
rect 17417 20009 17451 20043
rect 18521 20009 18555 20043
rect 19073 20009 19107 20043
rect 19625 20009 19659 20043
rect 11989 19941 12023 19975
rect 9137 19873 9171 19907
rect 10149 19873 10183 19907
rect 12633 19873 12667 19907
rect 13185 19873 13219 19907
rect 13829 19873 13863 19907
rect 14381 19873 14415 19907
rect 15577 19873 15611 19907
rect 16129 19873 16163 19907
rect 16681 19873 16715 19907
rect 17233 19873 17267 19907
rect 18337 19873 18371 19907
rect 18889 19873 18923 19907
rect 19441 19873 19475 19907
rect 19993 19873 20027 19907
rect 20545 19873 20579 19907
rect 9229 19805 9263 19839
rect 10241 19805 10275 19839
rect 10333 19805 10367 19839
rect 12173 19805 12207 19839
rect 16313 19737 16347 19771
rect 8677 19669 8711 19703
rect 9781 19669 9815 19703
rect 11529 19669 11563 19703
rect 14013 19669 14047 19703
rect 20177 19669 20211 19703
rect 20729 19669 20763 19703
rect 19073 19465 19107 19499
rect 8401 19261 8435 19295
rect 10057 19261 10091 19295
rect 11713 19261 11747 19295
rect 12449 19261 12483 19295
rect 14105 19261 14139 19295
rect 14657 19261 14691 19295
rect 15209 19261 15243 19295
rect 15761 19261 15795 19295
rect 16497 19261 16531 19295
rect 17141 19261 17175 19295
rect 17417 19261 17451 19295
rect 18061 19261 18095 19295
rect 18889 19261 18923 19295
rect 19441 19261 19475 19295
rect 19993 19261 20027 19295
rect 20545 19261 20579 19295
rect 8668 19193 8702 19227
rect 10302 19193 10336 19227
rect 12694 19193 12728 19227
rect 9781 19125 9815 19159
rect 11437 19125 11471 19159
rect 11897 19125 11931 19159
rect 13829 19125 13863 19159
rect 14289 19125 14323 19159
rect 14841 19125 14875 19159
rect 15393 19125 15427 19159
rect 15945 19125 15979 19159
rect 16681 19125 16715 19159
rect 18245 19125 18279 19159
rect 19625 19125 19659 19159
rect 20177 19125 20211 19159
rect 20729 19125 20763 19159
rect 9045 18921 9079 18955
rect 10149 18921 10183 18955
rect 11989 18921 12023 18955
rect 15669 18921 15703 18955
rect 10876 18853 10910 18887
rect 12900 18853 12934 18887
rect 19165 18853 19199 18887
rect 19901 18853 19935 18887
rect 7665 18785 7699 18819
rect 7932 18785 7966 18819
rect 12633 18785 12667 18819
rect 14657 18785 14691 18819
rect 15485 18785 15519 18819
rect 16293 18785 16327 18819
rect 18061 18785 18095 18819
rect 18889 18785 18923 18819
rect 19625 18785 19659 18819
rect 10609 18717 10643 18751
rect 16037 18717 16071 18751
rect 18153 18717 18187 18751
rect 18337 18717 18371 18751
rect 14013 18581 14047 18615
rect 14841 18581 14875 18615
rect 17417 18581 17451 18615
rect 17693 18581 17727 18615
rect 17601 18377 17635 18411
rect 18061 18377 18095 18411
rect 9873 18309 9907 18343
rect 9321 18241 9355 18275
rect 9505 18241 9539 18275
rect 10517 18241 10551 18275
rect 11529 18241 11563 18275
rect 13369 18241 13403 18275
rect 18613 18241 18647 18275
rect 10241 18173 10275 18207
rect 11253 18173 11287 18207
rect 13737 18173 13771 18207
rect 14004 18173 14038 18207
rect 15393 18173 15427 18207
rect 17417 18173 17451 18207
rect 19257 18173 19291 18207
rect 19809 18173 19843 18207
rect 20545 18173 20579 18207
rect 15638 18105 15672 18139
rect 20085 18105 20119 18139
rect 8861 18037 8895 18071
rect 9229 18037 9263 18071
rect 10333 18037 10367 18071
rect 12725 18037 12759 18071
rect 13093 18037 13127 18071
rect 13185 18037 13219 18071
rect 15117 18037 15151 18071
rect 16773 18037 16807 18071
rect 18429 18037 18463 18071
rect 18521 18037 18555 18071
rect 19441 18037 19475 18071
rect 20729 18037 20763 18071
rect 8769 17833 8803 17867
rect 10701 17833 10735 17867
rect 13001 17833 13035 17867
rect 18337 17833 18371 17867
rect 18613 17833 18647 17867
rect 13369 17765 13403 17799
rect 14749 17765 14783 17799
rect 16497 17765 16531 17799
rect 18981 17765 19015 17799
rect 19993 17765 20027 17799
rect 7389 17697 7423 17731
rect 7656 17697 7690 17731
rect 10609 17697 10643 17731
rect 11253 17697 11287 17731
rect 11529 17697 11563 17731
rect 11989 17697 12023 17731
rect 12265 17697 12299 17731
rect 14013 17697 14047 17731
rect 14289 17697 14323 17731
rect 15853 17697 15887 17731
rect 17224 17697 17258 17731
rect 19717 17697 19751 17731
rect 10885 17629 10919 17663
rect 13461 17629 13495 17663
rect 13553 17629 13587 17663
rect 15945 17629 15979 17663
rect 16129 17629 16163 17663
rect 16957 17629 16991 17663
rect 19073 17629 19107 17663
rect 19165 17629 19199 17663
rect 10241 17493 10275 17527
rect 15485 17493 15519 17527
rect 8401 17289 8435 17323
rect 12541 17289 12575 17323
rect 15393 17289 15427 17323
rect 10701 17221 10735 17255
rect 17049 17221 17083 17255
rect 17785 17221 17819 17255
rect 7021 17153 7055 17187
rect 9229 17153 9263 17187
rect 10241 17153 10275 17187
rect 11253 17153 11287 17187
rect 13001 17153 13035 17187
rect 13185 17153 13219 17187
rect 14105 17153 14139 17187
rect 15945 17153 15979 17187
rect 11161 17085 11195 17119
rect 15853 17085 15887 17119
rect 16865 17085 16899 17119
rect 17417 17085 17451 17119
rect 19993 17153 20027 17187
rect 20821 17153 20855 17187
rect 18061 17085 18095 17119
rect 19809 17085 19843 17119
rect 20545 17085 20579 17119
rect 7288 17017 7322 17051
rect 10057 17017 10091 17051
rect 11897 17017 11931 17051
rect 13921 17017 13955 17051
rect 15761 17017 15795 17051
rect 16405 17017 16439 17051
rect 17785 17017 17819 17051
rect 18328 17017 18362 17051
rect 8677 16949 8711 16983
rect 9045 16949 9079 16983
rect 9137 16949 9171 16983
rect 9689 16949 9723 16983
rect 10149 16949 10183 16983
rect 11069 16949 11103 16983
rect 12909 16949 12943 16983
rect 13553 16949 13587 16983
rect 14013 16949 14047 16983
rect 17601 16949 17635 16983
rect 19441 16949 19475 16983
rect 7021 16745 7055 16779
rect 8585 16745 8619 16779
rect 9137 16745 9171 16779
rect 12449 16745 12483 16779
rect 13093 16745 13127 16779
rect 13461 16745 13495 16779
rect 14197 16745 14231 16779
rect 14657 16745 14691 16779
rect 16589 16745 16623 16779
rect 18245 16745 18279 16779
rect 18613 16745 18647 16779
rect 19257 16745 19291 16779
rect 7389 16677 7423 16711
rect 12541 16677 12575 16711
rect 14565 16677 14599 16711
rect 15853 16677 15887 16711
rect 19625 16677 19659 16711
rect 20913 16677 20947 16711
rect 6837 16609 6871 16643
rect 7481 16609 7515 16643
rect 8493 16609 8527 16643
rect 10333 16609 10367 16643
rect 10692 16609 10726 16643
rect 15761 16609 15795 16643
rect 16405 16609 16439 16643
rect 16957 16609 16991 16643
rect 17509 16609 17543 16643
rect 17785 16609 17819 16643
rect 18705 16609 18739 16643
rect 20269 16609 20303 16643
rect 7665 16541 7699 16575
rect 8677 16541 8711 16575
rect 10425 16541 10459 16575
rect 12633 16541 12667 16575
rect 13553 16541 13587 16575
rect 13737 16541 13771 16575
rect 14841 16541 14875 16575
rect 15945 16541 15979 16575
rect 18889 16541 18923 16575
rect 19717 16541 19751 16575
rect 19809 16541 19843 16575
rect 8125 16473 8159 16507
rect 15393 16473 15427 16507
rect 10149 16405 10183 16439
rect 11805 16405 11839 16439
rect 12081 16405 12115 16439
rect 17141 16405 17175 16439
rect 20453 16405 20487 16439
rect 19441 16201 19475 16235
rect 16773 16133 16807 16167
rect 16865 16133 16899 16167
rect 19717 16133 19751 16167
rect 8953 16065 8987 16099
rect 11621 16065 11655 16099
rect 11713 16065 11747 16099
rect 12449 16065 12483 16099
rect 16497 16065 16531 16099
rect 6837 15997 6871 16031
rect 8677 15997 8711 16031
rect 9505 15997 9539 16031
rect 11529 15997 11563 16031
rect 14197 15997 14231 16031
rect 14464 15997 14498 16031
rect 16313 15997 16347 16031
rect 17509 16065 17543 16099
rect 20269 16065 20303 16099
rect 18061 15997 18095 16031
rect 18328 15997 18362 16031
rect 20729 15997 20763 16031
rect 7104 15929 7138 15963
rect 9772 15929 9806 15963
rect 12716 15929 12750 15963
rect 16773 15929 16807 15963
rect 17325 15929 17359 15963
rect 20177 15929 20211 15963
rect 8217 15861 8251 15895
rect 10885 15861 10919 15895
rect 11161 15861 11195 15895
rect 13829 15861 13863 15895
rect 15577 15861 15611 15895
rect 15853 15861 15887 15895
rect 16221 15861 16255 15895
rect 17233 15861 17267 15895
rect 20085 15861 20119 15895
rect 20913 15861 20947 15895
rect 7849 15657 7883 15691
rect 10701 15657 10735 15691
rect 15025 15657 15059 15691
rect 15669 15657 15703 15691
rect 17969 15657 18003 15691
rect 11161 15589 11195 15623
rect 13820 15589 13854 15623
rect 6469 15521 6503 15555
rect 6736 15521 6770 15555
rect 9689 15521 9723 15555
rect 9965 15521 9999 15555
rect 11069 15521 11103 15555
rect 12081 15521 12115 15555
rect 12817 15521 12851 15555
rect 13093 15521 13127 15555
rect 11345 15453 11379 15487
rect 12173 15453 12207 15487
rect 12357 15453 12391 15487
rect 13553 15453 13587 15487
rect 15761 15589 15795 15623
rect 18696 15589 18730 15623
rect 16497 15521 16531 15555
rect 16856 15521 16890 15555
rect 18429 15521 18463 15555
rect 20085 15521 20119 15555
rect 15853 15453 15887 15487
rect 16221 15453 16255 15487
rect 16589 15453 16623 15487
rect 20269 15453 20303 15487
rect 15301 15385 15335 15419
rect 11713 15317 11747 15351
rect 14933 15317 14967 15351
rect 15025 15317 15059 15351
rect 16221 15317 16255 15351
rect 16313 15317 16347 15351
rect 19809 15317 19843 15351
rect 9137 15113 9171 15147
rect 9413 15113 9447 15147
rect 12449 15113 12483 15147
rect 16221 15113 16255 15147
rect 16405 15113 16439 15147
rect 6193 14977 6227 15011
rect 6377 14977 6411 15011
rect 7757 14977 7791 15011
rect 9965 14977 9999 15011
rect 10885 14977 10919 15011
rect 11805 14977 11839 15011
rect 11989 14977 12023 15011
rect 13093 14977 13127 15011
rect 13645 14977 13679 15011
rect 15853 14977 15887 15011
rect 16037 14977 16071 15011
rect 6101 14909 6135 14943
rect 10609 14909 10643 14943
rect 13912 14909 13946 14943
rect 8024 14841 8058 14875
rect 9873 14841 9907 14875
rect 12909 14841 12943 14875
rect 15761 14841 15795 14875
rect 19441 15045 19475 15079
rect 16865 14977 16899 15011
rect 17049 14977 17083 15011
rect 18889 14977 18923 15011
rect 19073 14977 19107 15011
rect 19993 14977 20027 15011
rect 20729 14977 20763 15011
rect 16773 14909 16807 14943
rect 20453 14909 20487 14943
rect 17417 14841 17451 14875
rect 19901 14841 19935 14875
rect 5733 14773 5767 14807
rect 9781 14773 9815 14807
rect 11345 14773 11379 14807
rect 11713 14773 11747 14807
rect 12817 14773 12851 14807
rect 15025 14773 15059 14807
rect 15393 14773 15427 14807
rect 16221 14773 16255 14807
rect 18429 14773 18463 14807
rect 18797 14773 18831 14807
rect 19809 14773 19843 14807
rect 8585 14569 8619 14603
rect 9045 14569 9079 14603
rect 9689 14569 9723 14603
rect 12449 14569 12483 14603
rect 14105 14569 14139 14603
rect 15301 14569 15335 14603
rect 15669 14569 15703 14603
rect 15761 14569 15795 14603
rect 17693 14569 17727 14603
rect 7196 14501 7230 14535
rect 8953 14501 8987 14535
rect 11336 14501 11370 14535
rect 12970 14501 13004 14535
rect 14657 14501 14691 14535
rect 18880 14501 18914 14535
rect 10057 14433 10091 14467
rect 10977 14433 11011 14467
rect 12725 14433 12759 14467
rect 14381 14433 14415 14467
rect 16580 14433 16614 14467
rect 18613 14433 18647 14467
rect 20269 14433 20303 14467
rect 6929 14365 6963 14399
rect 9229 14365 9263 14399
rect 10149 14365 10183 14399
rect 10241 14365 10275 14399
rect 11069 14365 11103 14399
rect 15853 14365 15887 14399
rect 16313 14365 16347 14399
rect 17969 14365 18003 14399
rect 20913 14365 20947 14399
rect 8309 14297 8343 14331
rect 10793 14229 10827 14263
rect 19993 14229 20027 14263
rect 20453 14229 20487 14263
rect 11345 14025 11379 14059
rect 12725 14025 12759 14059
rect 13553 14025 13587 14059
rect 13737 14025 13771 14059
rect 15945 14025 15979 14059
rect 17601 14025 17635 14059
rect 19717 14025 19751 14059
rect 20913 14025 20947 14059
rect 9229 13889 9263 13923
rect 11805 13889 11839 13923
rect 11989 13889 12023 13923
rect 13185 13889 13219 13923
rect 13369 13889 13403 13923
rect 9496 13821 9530 13855
rect 14197 13889 14231 13923
rect 14381 13889 14415 13923
rect 15577 13889 15611 13923
rect 18613 13889 18647 13923
rect 20269 13889 20303 13923
rect 15393 13821 15427 13855
rect 16121 13821 16155 13855
rect 16221 13821 16255 13855
rect 16488 13821 16522 13855
rect 20177 13821 20211 13855
rect 20729 13821 20763 13855
rect 8769 13753 8803 13787
rect 13093 13753 13127 13787
rect 13553 13753 13587 13787
rect 18521 13753 18555 13787
rect 20085 13753 20119 13787
rect 10609 13685 10643 13719
rect 11713 13685 11747 13719
rect 14105 13685 14139 13719
rect 14933 13685 14967 13719
rect 15301 13685 15335 13719
rect 18061 13685 18095 13719
rect 18429 13685 18463 13719
rect 9781 13481 9815 13515
rect 11253 13481 11287 13515
rect 13185 13481 13219 13515
rect 14565 13481 14599 13515
rect 16773 13481 16807 13515
rect 17233 13481 17267 13515
rect 17785 13481 17819 13515
rect 18153 13481 18187 13515
rect 18245 13481 18279 13515
rect 18797 13481 18831 13515
rect 19809 13481 19843 13515
rect 11161 13413 11195 13447
rect 13553 13413 13587 13447
rect 15301 13413 15335 13447
rect 10149 13345 10183 13379
rect 12357 13345 12391 13379
rect 16129 13345 16163 13379
rect 16221 13345 16255 13379
rect 17141 13345 17175 13379
rect 19165 13345 19199 13379
rect 20177 13345 20211 13379
rect 10241 13277 10275 13311
rect 10333 13277 10367 13311
rect 11345 13277 11379 13311
rect 12449 13277 12483 13311
rect 12633 13277 12667 13311
rect 13645 13277 13679 13311
rect 13829 13277 13863 13311
rect 14657 13277 14691 13311
rect 14749 13277 14783 13311
rect 16313 13277 16347 13311
rect 17417 13277 17451 13311
rect 18337 13277 18371 13311
rect 19257 13277 19291 13311
rect 19349 13277 19383 13311
rect 20269 13277 20303 13311
rect 20361 13277 20395 13311
rect 10793 13141 10827 13175
rect 11989 13141 12023 13175
rect 14197 13141 14231 13175
rect 15761 13141 15795 13175
rect 9137 12937 9171 12971
rect 10793 12937 10827 12971
rect 11069 12937 11103 12971
rect 13369 12937 13403 12971
rect 16589 12937 16623 12971
rect 18337 12937 18371 12971
rect 20085 12937 20119 12971
rect 12081 12869 12115 12903
rect 9413 12801 9447 12835
rect 11529 12801 11563 12835
rect 11621 12801 11655 12835
rect 12725 12801 12759 12835
rect 13829 12801 13863 12835
rect 14013 12801 14047 12835
rect 17049 12801 17083 12835
rect 17233 12801 17267 12835
rect 18705 12801 18739 12835
rect 20913 12801 20947 12835
rect 9321 12733 9355 12767
rect 9680 12733 9714 12767
rect 12265 12733 12299 12767
rect 12449 12733 12483 12767
rect 14381 12733 14415 12767
rect 16405 12733 16439 12767
rect 16957 12733 16991 12767
rect 18153 12733 18187 12767
rect 18972 12733 19006 12767
rect 11437 12665 11471 12699
rect 14626 12665 14660 12699
rect 20821 12665 20855 12699
rect 13737 12597 13771 12631
rect 15761 12597 15795 12631
rect 16221 12597 16255 12631
rect 20361 12597 20395 12631
rect 20729 12597 20763 12631
rect 11069 12393 11103 12427
rect 12817 12393 12851 12427
rect 17877 12393 17911 12427
rect 19993 12393 20027 12427
rect 20453 12393 20487 12427
rect 7748 12325 7782 12359
rect 13728 12325 13762 12359
rect 16006 12325 16040 12359
rect 17785 12325 17819 12359
rect 9689 12257 9723 12291
rect 9956 12257 9990 12291
rect 11704 12257 11738 12291
rect 18880 12257 18914 12291
rect 20269 12257 20303 12291
rect 7481 12189 7515 12223
rect 9137 12189 9171 12223
rect 11437 12189 11471 12223
rect 13461 12189 13495 12223
rect 15301 12189 15335 12223
rect 15761 12189 15795 12223
rect 17969 12189 18003 12223
rect 18613 12189 18647 12223
rect 20913 12189 20947 12223
rect 8861 12053 8895 12087
rect 14841 12053 14875 12087
rect 17141 12053 17175 12087
rect 17417 12053 17451 12087
rect 10241 11849 10275 11883
rect 11345 11849 11379 11883
rect 13921 11849 13955 11883
rect 18705 11849 18739 11883
rect 8309 11781 8343 11815
rect 18337 11781 18371 11815
rect 8861 11713 8895 11747
rect 10885 11713 10919 11747
rect 11989 11713 12023 11747
rect 14565 11713 14599 11747
rect 15945 11713 15979 11747
rect 17509 11713 17543 11747
rect 19257 11713 19291 11747
rect 19717 11713 19751 11747
rect 9321 11645 9355 11679
rect 10609 11645 10643 11679
rect 12449 11645 12483 11679
rect 17233 11645 17267 11679
rect 18153 11645 18187 11679
rect 19073 11645 19107 11679
rect 9597 11577 9631 11611
rect 12694 11577 12728 11611
rect 14381 11577 14415 11611
rect 19984 11577 20018 11611
rect 8677 11509 8711 11543
rect 8769 11509 8803 11543
rect 10701 11509 10735 11543
rect 11713 11509 11747 11543
rect 11805 11509 11839 11543
rect 13829 11509 13863 11543
rect 14289 11509 14323 11543
rect 15393 11509 15427 11543
rect 15761 11509 15795 11543
rect 15853 11509 15887 11543
rect 16865 11509 16899 11543
rect 17325 11509 17359 11543
rect 19165 11509 19199 11543
rect 21097 11509 21131 11543
rect 9045 11305 9079 11339
rect 9781 11305 9815 11339
rect 12449 11305 12483 11339
rect 14381 11305 14415 11339
rect 15945 11305 15979 11339
rect 17969 11305 18003 11339
rect 19809 11305 19843 11339
rect 10149 11237 10183 11271
rect 10241 11237 10275 11271
rect 13093 11237 13127 11271
rect 16037 11237 16071 11271
rect 19165 11237 19199 11271
rect 7389 11169 7423 11203
rect 7656 11169 7690 11203
rect 10793 11169 10827 11203
rect 11060 11169 11094 11203
rect 16856 11169 16890 11203
rect 20177 11169 20211 11203
rect 10425 11101 10459 11135
rect 16221 11101 16255 11135
rect 16589 11101 16623 11135
rect 19257 11101 19291 11135
rect 19349 11101 19383 11135
rect 20269 11101 20303 11135
rect 20361 11101 20395 11135
rect 8769 11033 8803 11067
rect 12173 10965 12207 10999
rect 15577 10965 15611 10999
rect 18797 10965 18831 10999
rect 8493 10761 8527 10795
rect 12449 10761 12483 10795
rect 13277 10761 13311 10795
rect 15301 10761 15335 10795
rect 10609 10693 10643 10727
rect 9045 10625 9079 10659
rect 11161 10625 11195 10659
rect 11897 10625 11931 10659
rect 13093 10625 13127 10659
rect 13829 10625 13863 10659
rect 14933 10625 14967 10659
rect 15945 10625 15979 10659
rect 18061 10625 18095 10659
rect 19257 10625 19291 10659
rect 8953 10557 8987 10591
rect 9505 10557 9539 10591
rect 11621 10557 11655 10591
rect 13737 10557 13771 10591
rect 14749 10557 14783 10591
rect 15669 10557 15703 10591
rect 16313 10557 16347 10591
rect 16580 10557 16614 10591
rect 18981 10557 19015 10591
rect 19625 10557 19659 10591
rect 9781 10489 9815 10523
rect 14657 10489 14691 10523
rect 19073 10489 19107 10523
rect 19892 10489 19926 10523
rect 8861 10421 8895 10455
rect 10977 10421 11011 10455
rect 11069 10421 11103 10455
rect 12817 10421 12851 10455
rect 12909 10421 12943 10455
rect 13645 10421 13679 10455
rect 14289 10421 14323 10455
rect 15761 10421 15795 10455
rect 17693 10421 17727 10455
rect 18613 10421 18647 10455
rect 21005 10421 21039 10455
rect 11805 10217 11839 10251
rect 12357 10217 12391 10251
rect 13829 10217 13863 10251
rect 14381 10217 14415 10251
rect 14841 10217 14875 10251
rect 15761 10217 15795 10251
rect 17141 10217 17175 10251
rect 17601 10217 17635 10251
rect 18153 10217 18187 10251
rect 20545 10217 20579 10251
rect 7932 10149 7966 10183
rect 10692 10149 10726 10183
rect 13185 10149 13219 10183
rect 14749 10149 14783 10183
rect 16681 10149 16715 10183
rect 12725 10081 12759 10115
rect 13737 10081 13771 10115
rect 15669 10081 15703 10115
rect 16129 10081 16163 10115
rect 16405 10081 16439 10115
rect 17509 10081 17543 10115
rect 18521 10081 18555 10115
rect 19421 10081 19455 10115
rect 7665 10013 7699 10047
rect 9689 10013 9723 10047
rect 10425 10013 10459 10047
rect 12817 10013 12851 10047
rect 13001 10013 13035 10047
rect 13185 10013 13219 10047
rect 13921 10013 13955 10047
rect 14933 10013 14967 10047
rect 15853 10013 15887 10047
rect 17785 10013 17819 10047
rect 18613 10013 18647 10047
rect 18797 10013 18831 10047
rect 19165 10013 19199 10047
rect 15301 9945 15335 9979
rect 9045 9877 9079 9911
rect 13369 9877 13403 9911
rect 15945 9673 15979 9707
rect 11161 9605 11195 9639
rect 16221 9605 16255 9639
rect 18061 9605 18095 9639
rect 8033 9537 8067 9571
rect 16773 9537 16807 9571
rect 18613 9537 18647 9571
rect 19349 9537 19383 9571
rect 20453 9537 20487 9571
rect 20637 9537 20671 9571
rect 9781 9469 9815 9503
rect 12449 9469 12483 9503
rect 14289 9469 14323 9503
rect 14473 9469 14507 9503
rect 14565 9469 14599 9503
rect 19073 9469 19107 9503
rect 8300 9401 8334 9435
rect 10048 9401 10082 9435
rect 12716 9401 12750 9435
rect 14832 9401 14866 9435
rect 16681 9401 16715 9435
rect 18429 9401 18463 9435
rect 9413 9333 9447 9367
rect 11437 9333 11471 9367
rect 13829 9333 13863 9367
rect 14105 9333 14139 9367
rect 14473 9333 14507 9367
rect 16589 9333 16623 9367
rect 18521 9333 18555 9367
rect 19993 9333 20027 9367
rect 20361 9333 20395 9367
rect 8585 9129 8619 9163
rect 8953 9129 8987 9163
rect 10425 9129 10459 9163
rect 10701 9129 10735 9163
rect 11069 9129 11103 9163
rect 15301 9129 15335 9163
rect 15669 9129 15703 9163
rect 18429 9129 18463 9163
rect 20361 9129 20395 9163
rect 12173 9061 12207 9095
rect 13084 9061 13118 9095
rect 17316 9061 17350 9095
rect 18972 9061 19006 9095
rect 10609 8993 10643 9027
rect 11161 8993 11195 9027
rect 12081 8993 12115 9027
rect 12817 8993 12851 9027
rect 16957 8993 16991 9027
rect 9045 8925 9079 8959
rect 9229 8925 9263 8959
rect 11253 8925 11287 8959
rect 12265 8925 12299 8959
rect 15761 8925 15795 8959
rect 15853 8925 15887 8959
rect 17049 8925 17083 8959
rect 18705 8925 18739 8959
rect 16773 8857 16807 8891
rect 11713 8789 11747 8823
rect 14197 8789 14231 8823
rect 20085 8789 20119 8823
rect 8585 8585 8619 8619
rect 11345 8585 11379 8619
rect 16957 8585 16991 8619
rect 12633 8517 12667 8551
rect 14197 8517 14231 8551
rect 19533 8517 19567 8551
rect 9137 8449 9171 8483
rect 11897 8449 11931 8483
rect 13737 8449 13771 8483
rect 14749 8449 14783 8483
rect 15577 8449 15611 8483
rect 18613 8449 18647 8483
rect 20085 8449 20119 8483
rect 9045 8381 9079 8415
rect 9689 8381 9723 8415
rect 11713 8381 11747 8415
rect 12817 8381 12851 8415
rect 13553 8381 13587 8415
rect 14565 8381 14599 8415
rect 15393 8381 15427 8415
rect 18521 8381 18555 8415
rect 19901 8381 19935 8415
rect 8953 8313 8987 8347
rect 9956 8313 9990 8347
rect 13645 8313 13679 8347
rect 14657 8313 14691 8347
rect 15844 8313 15878 8347
rect 18429 8313 18463 8347
rect 11069 8245 11103 8279
rect 11805 8245 11839 8279
rect 13185 8245 13219 8279
rect 15209 8245 15243 8279
rect 17233 8245 17267 8279
rect 18061 8245 18095 8279
rect 19993 8245 20027 8279
rect 10149 8041 10183 8075
rect 14933 8041 14967 8075
rect 20269 8041 20303 8075
rect 20913 8041 20947 8075
rect 10517 7973 10551 8007
rect 11428 7973 11462 8007
rect 13820 7973 13854 8007
rect 16948 7973 16982 8007
rect 8861 7905 8895 7939
rect 10609 7905 10643 7939
rect 16037 7905 16071 7939
rect 18889 7905 18923 7939
rect 19156 7905 19190 7939
rect 9137 7837 9171 7871
rect 10793 7837 10827 7871
rect 11161 7837 11195 7871
rect 13553 7837 13587 7871
rect 16129 7837 16163 7871
rect 16313 7837 16347 7871
rect 16681 7837 16715 7871
rect 12541 7701 12575 7735
rect 15669 7701 15703 7735
rect 18061 7701 18095 7735
rect 10517 7497 10551 7531
rect 16681 7497 16715 7531
rect 16957 7497 16991 7531
rect 18061 7497 18095 7531
rect 20085 7497 20119 7531
rect 11989 7361 12023 7395
rect 13737 7361 13771 7395
rect 14749 7361 14783 7395
rect 15301 7361 15335 7395
rect 17509 7361 17543 7395
rect 18613 7361 18647 7395
rect 19625 7361 19659 7395
rect 20637 7361 20671 7395
rect 9137 7293 9171 7327
rect 11805 7293 11839 7327
rect 14657 7293 14691 7327
rect 15568 7293 15602 7327
rect 17325 7293 17359 7327
rect 17417 7293 17451 7327
rect 19441 7293 19475 7327
rect 20545 7293 20579 7327
rect 9404 7225 9438 7259
rect 11713 7225 11747 7259
rect 12725 7225 12759 7259
rect 13553 7225 13587 7259
rect 14565 7225 14599 7259
rect 18429 7225 18463 7259
rect 11345 7157 11379 7191
rect 13185 7157 13219 7191
rect 13645 7157 13679 7191
rect 14197 7157 14231 7191
rect 18521 7157 18555 7191
rect 19073 7157 19107 7191
rect 19533 7157 19567 7191
rect 20453 7157 20487 7191
rect 9689 6953 9723 6987
rect 14105 6953 14139 6987
rect 18521 6953 18555 6987
rect 20545 6953 20579 6987
rect 11796 6885 11830 6919
rect 15669 6885 15703 6919
rect 8208 6817 8242 6851
rect 10057 6817 10091 6851
rect 10977 6817 11011 6851
rect 14197 6817 14231 6851
rect 16957 6817 16991 6851
rect 17408 6817 17442 6851
rect 19432 6817 19466 6851
rect 7941 6749 7975 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 11529 6749 11563 6783
rect 14289 6749 14323 6783
rect 15761 6749 15795 6783
rect 15945 6749 15979 6783
rect 16313 6749 16347 6783
rect 17141 6749 17175 6783
rect 19165 6749 19199 6783
rect 9321 6681 9355 6715
rect 13737 6681 13771 6715
rect 16773 6681 16807 6715
rect 10793 6613 10827 6647
rect 12909 6613 12943 6647
rect 15301 6613 15335 6647
rect 9045 6409 9079 6443
rect 9321 6409 9355 6443
rect 10333 6409 10367 6443
rect 15301 6409 15335 6443
rect 18061 6409 18095 6443
rect 9873 6273 9907 6307
rect 10885 6273 10919 6307
rect 11897 6273 11931 6307
rect 13001 6273 13035 6307
rect 14105 6273 14139 6307
rect 15853 6273 15887 6307
rect 16865 6273 16899 6307
rect 18613 6273 18647 6307
rect 19717 6273 19751 6307
rect 19901 6273 19935 6307
rect 20821 6273 20855 6307
rect 7665 6205 7699 6239
rect 11713 6205 11747 6239
rect 16681 6205 16715 6239
rect 18429 6205 18463 6239
rect 20637 6205 20671 6239
rect 7910 6137 7944 6171
rect 9689 6137 9723 6171
rect 10701 6137 10735 6171
rect 11805 6137 11839 6171
rect 12817 6137 12851 6171
rect 13921 6137 13955 6171
rect 18521 6137 18555 6171
rect 20729 6137 20763 6171
rect 9781 6069 9815 6103
rect 10793 6069 10827 6103
rect 11345 6069 11379 6103
rect 12449 6069 12483 6103
rect 12909 6069 12943 6103
rect 13461 6069 13495 6103
rect 13829 6069 13863 6103
rect 15669 6069 15703 6103
rect 15761 6069 15795 6103
rect 16313 6069 16347 6103
rect 16773 6069 16807 6103
rect 19257 6069 19291 6103
rect 19625 6069 19659 6103
rect 20269 6069 20303 6103
rect 7849 5865 7883 5899
rect 9137 5865 9171 5899
rect 9689 5865 9723 5899
rect 13001 5865 13035 5899
rect 16681 5865 16715 5899
rect 18521 5865 18555 5899
rect 20913 5865 20947 5899
rect 6714 5797 6748 5831
rect 11152 5797 11186 5831
rect 15546 5797 15580 5831
rect 17386 5797 17420 5831
rect 19064 5797 19098 5831
rect 6469 5729 6503 5763
rect 10057 5729 10091 5763
rect 12909 5729 12943 5763
rect 13921 5729 13955 5763
rect 14013 5729 14047 5763
rect 15301 5729 15335 5763
rect 17141 5729 17175 5763
rect 18797 5729 18831 5763
rect 10149 5661 10183 5695
rect 10333 5661 10367 5695
rect 10885 5661 10919 5695
rect 13185 5661 13219 5695
rect 14105 5661 14139 5695
rect 12265 5593 12299 5627
rect 12541 5525 12575 5559
rect 13553 5525 13587 5559
rect 20177 5525 20211 5559
rect 10333 5321 10367 5355
rect 13829 5321 13863 5355
rect 14013 5321 14047 5355
rect 20637 5321 20671 5355
rect 10793 5185 10827 5219
rect 10977 5185 11011 5219
rect 12449 5185 12483 5219
rect 15945 5185 15979 5219
rect 18889 5185 18923 5219
rect 12716 5117 12750 5151
rect 14013 5117 14047 5151
rect 14105 5117 14139 5151
rect 14361 5117 14395 5151
rect 16212 5117 16246 5151
rect 18613 5117 18647 5151
rect 19257 5117 19291 5151
rect 10701 5049 10735 5083
rect 19524 5049 19558 5083
rect 11897 4981 11931 5015
rect 15485 4981 15519 5015
rect 17325 4981 17359 5015
rect 18245 4981 18279 5015
rect 18705 4981 18739 5015
rect 12449 4777 12483 4811
rect 12909 4777 12943 4811
rect 16037 4777 16071 4811
rect 18061 4777 18095 4811
rect 19625 4777 19659 4811
rect 19993 4777 20027 4811
rect 16129 4709 16163 4743
rect 12817 4641 12851 4675
rect 13829 4641 13863 4675
rect 13921 4641 13955 4675
rect 14473 4641 14507 4675
rect 18429 4641 18463 4675
rect 19073 4641 19107 4675
rect 13001 4573 13035 4607
rect 14105 4573 14139 4607
rect 16313 4573 16347 4607
rect 18521 4573 18555 4607
rect 18705 4573 18739 4607
rect 20085 4573 20119 4607
rect 20177 4573 20211 4607
rect 13461 4505 13495 4539
rect 14657 4437 14691 4471
rect 15669 4437 15703 4471
rect 19441 4233 19475 4267
rect 19717 4233 19751 4267
rect 14565 4097 14599 4131
rect 15853 4097 15887 4131
rect 20269 4097 20303 4131
rect 8953 4029 8987 4063
rect 9220 4029 9254 4063
rect 11793 4029 11827 4063
rect 12725 4029 12759 4063
rect 13001 4029 13035 4063
rect 15761 4029 15795 4063
rect 16313 4029 16347 4063
rect 17417 4029 17451 4063
rect 18061 4029 18095 4063
rect 20177 4029 20211 4063
rect 20729 4029 20763 4063
rect 13461 3961 13495 3995
rect 14289 3961 14323 3995
rect 15669 3961 15703 3995
rect 16589 3961 16623 3995
rect 18328 3961 18362 3995
rect 10333 3893 10367 3927
rect 10977 3893 11011 3927
rect 11989 3893 12023 3927
rect 13921 3893 13955 3927
rect 14381 3893 14415 3927
rect 15301 3893 15335 3927
rect 17601 3893 17635 3927
rect 20085 3893 20119 3927
rect 20913 3893 20947 3927
rect 13001 3689 13035 3723
rect 14657 3689 14691 3723
rect 16957 3689 16991 3723
rect 18613 3689 18647 3723
rect 10232 3621 10266 3655
rect 11437 3621 11471 3655
rect 11866 3621 11900 3655
rect 13522 3621 13556 3655
rect 15844 3621 15878 3655
rect 17478 3621 17512 3655
rect 9965 3485 9999 3519
rect 11621 3553 11655 3587
rect 13277 3553 13311 3587
rect 15577 3553 15611 3587
rect 17233 3553 17267 3587
rect 19073 3553 19107 3587
rect 19809 3553 19843 3587
rect 19349 3485 19383 3519
rect 20085 3485 20119 3519
rect 11345 3417 11379 3451
rect 11437 3417 11471 3451
rect 10333 3145 10367 3179
rect 10517 3145 10551 3179
rect 10701 3145 10735 3179
rect 13277 3145 13311 3179
rect 16497 3145 16531 3179
rect 18061 3145 18095 3179
rect 6561 3077 6595 3111
rect 15669 3077 15703 3111
rect 19533 3077 19567 3111
rect 10517 3009 10551 3043
rect 11345 3009 11379 3043
rect 13921 3009 13955 3043
rect 17141 3009 17175 3043
rect 18613 3009 18647 3043
rect 10149 2941 10183 2975
rect 11069 2941 11103 2975
rect 11805 2941 11839 2975
rect 12449 2941 12483 2975
rect 13645 2941 13679 2975
rect 14289 2941 14323 2975
rect 14556 2941 14590 2975
rect 15945 2941 15979 2975
rect 18521 2941 18555 2975
rect 19349 2941 19383 2975
rect 19993 2941 20027 2975
rect 20545 2941 20579 2975
rect 12725 2873 12759 2907
rect 16865 2873 16899 2907
rect 17509 2873 17543 2907
rect 18429 2873 18463 2907
rect 18889 2873 18923 2907
rect 6561 2805 6595 2839
rect 11161 2805 11195 2839
rect 11989 2805 12023 2839
rect 13737 2805 13771 2839
rect 16129 2805 16163 2839
rect 16957 2805 16991 2839
rect 20177 2805 20211 2839
rect 20729 2805 20763 2839
rect 10333 2601 10367 2635
rect 15853 2601 15887 2635
rect 15945 2601 15979 2635
rect 13645 2533 13679 2567
rect 10701 2465 10735 2499
rect 10793 2465 10827 2499
rect 11437 2465 11471 2499
rect 11989 2465 12023 2499
rect 12633 2465 12667 2499
rect 13369 2465 13403 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 16497 2465 16531 2499
rect 17325 2465 17359 2499
rect 18337 2465 18371 2499
rect 18981 2465 19015 2499
rect 19533 2465 19567 2499
rect 20361 2465 20395 2499
rect 10885 2397 10919 2431
rect 12817 2397 12851 2431
rect 16037 2397 16071 2431
rect 11621 2329 11655 2363
rect 14473 2329 14507 2363
rect 19717 2329 19751 2363
rect 12173 2261 12207 2295
rect 15025 2261 15059 2295
rect 15485 2261 15519 2295
rect 16681 2261 16715 2295
rect 17509 2261 17543 2295
rect 18521 2261 18555 2295
rect 19165 2261 19199 2295
rect 20545 2261 20579 2295
<< metal1 >>
rect 13262 20680 13268 20732
rect 13320 20720 13326 20732
rect 17954 20720 17960 20732
rect 13320 20692 17960 20720
rect 13320 20680 13326 20692
rect 17954 20680 17960 20692
rect 18012 20680 18018 20732
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 9033 20043 9091 20049
rect 9033 20009 9045 20043
rect 9079 20040 9091 20043
rect 9122 20040 9128 20052
rect 9079 20012 9128 20040
rect 9079 20009 9091 20012
rect 9033 20003 9091 20009
rect 9122 20000 9128 20012
rect 9180 20000 9186 20052
rect 11330 20000 11336 20052
rect 11388 20040 11394 20052
rect 11885 20043 11943 20049
rect 11885 20040 11897 20043
rect 11388 20012 11897 20040
rect 11388 20000 11394 20012
rect 11885 20009 11897 20012
rect 11931 20009 11943 20043
rect 11885 20003 11943 20009
rect 12526 20000 12532 20052
rect 12584 20040 12590 20052
rect 12805 20043 12863 20049
rect 12805 20040 12817 20043
rect 12584 20012 12817 20040
rect 12584 20000 12590 20012
rect 12805 20009 12817 20012
rect 12851 20009 12863 20043
rect 12805 20003 12863 20009
rect 13078 20000 13084 20052
rect 13136 20040 13142 20052
rect 13357 20043 13415 20049
rect 13357 20040 13369 20043
rect 13136 20012 13369 20040
rect 13136 20000 13142 20012
rect 13357 20009 13369 20012
rect 13403 20009 13415 20043
rect 13357 20003 13415 20009
rect 14553 20043 14611 20049
rect 14553 20009 14565 20043
rect 14599 20040 14611 20043
rect 15286 20040 15292 20052
rect 14599 20012 15292 20040
rect 14599 20009 14611 20012
rect 14553 20003 14611 20009
rect 15286 20000 15292 20012
rect 15344 20000 15350 20052
rect 15749 20043 15807 20049
rect 15749 20009 15761 20043
rect 15795 20009 15807 20043
rect 15749 20003 15807 20009
rect 16853 20043 16911 20049
rect 16853 20009 16865 20043
rect 16899 20040 16911 20043
rect 16942 20040 16948 20052
rect 16899 20012 16948 20040
rect 16899 20009 16911 20012
rect 16853 20003 16911 20009
rect 7466 19932 7472 19984
rect 7524 19972 7530 19984
rect 11606 19972 11612 19984
rect 7524 19944 11612 19972
rect 7524 19932 7530 19944
rect 11606 19932 11612 19944
rect 11664 19972 11670 19984
rect 11977 19975 12035 19981
rect 11977 19972 11989 19975
rect 11664 19944 11989 19972
rect 11664 19932 11670 19944
rect 11977 19941 11989 19944
rect 12023 19941 12035 19975
rect 15764 19972 15792 20003
rect 16942 20000 16948 20012
rect 17000 20000 17006 20052
rect 17405 20043 17463 20049
rect 17405 20009 17417 20043
rect 17451 20040 17463 20043
rect 17494 20040 17500 20052
rect 17451 20012 17500 20040
rect 17451 20009 17463 20012
rect 17405 20003 17463 20009
rect 17494 20000 17500 20012
rect 17552 20000 17558 20052
rect 18506 20040 18512 20052
rect 18467 20012 18512 20040
rect 18506 20000 18512 20012
rect 18564 20000 18570 20052
rect 19058 20040 19064 20052
rect 19019 20012 19064 20040
rect 19058 20000 19064 20012
rect 19116 20000 19122 20052
rect 19150 20000 19156 20052
rect 19208 20000 19214 20052
rect 19242 20000 19248 20052
rect 19300 20040 19306 20052
rect 19613 20043 19671 20049
rect 19613 20040 19625 20043
rect 19300 20012 19625 20040
rect 19300 20000 19306 20012
rect 19613 20009 19625 20012
rect 19659 20009 19671 20043
rect 19613 20003 19671 20009
rect 19168 19972 19196 20000
rect 15764 19944 19196 19972
rect 11977 19935 12035 19941
rect 6362 19864 6368 19916
rect 6420 19904 6426 19916
rect 9125 19907 9183 19913
rect 9125 19904 9137 19907
rect 6420 19876 9137 19904
rect 6420 19864 6426 19876
rect 9125 19873 9137 19876
rect 9171 19904 9183 19907
rect 9398 19904 9404 19916
rect 9171 19876 9404 19904
rect 9171 19873 9183 19876
rect 9125 19867 9183 19873
rect 9398 19864 9404 19876
rect 9456 19864 9462 19916
rect 10134 19904 10140 19916
rect 10095 19876 10140 19904
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 12250 19864 12256 19916
rect 12308 19904 12314 19916
rect 12621 19907 12679 19913
rect 12621 19904 12633 19907
rect 12308 19876 12633 19904
rect 12308 19864 12314 19876
rect 12621 19873 12633 19876
rect 12667 19873 12679 19907
rect 12621 19867 12679 19873
rect 12986 19864 12992 19916
rect 13044 19904 13050 19916
rect 13173 19907 13231 19913
rect 13173 19904 13185 19907
rect 13044 19876 13185 19904
rect 13044 19864 13050 19876
rect 13173 19873 13185 19876
rect 13219 19873 13231 19907
rect 13173 19867 13231 19873
rect 13817 19907 13875 19913
rect 13817 19873 13829 19907
rect 13863 19873 13875 19907
rect 13817 19867 13875 19873
rect 9214 19796 9220 19848
rect 9272 19836 9278 19848
rect 10226 19836 10232 19848
rect 9272 19808 9317 19836
rect 10187 19808 10232 19836
rect 9272 19796 9278 19808
rect 10226 19796 10232 19808
rect 10284 19796 10290 19848
rect 10318 19796 10324 19848
rect 10376 19836 10382 19848
rect 12161 19839 12219 19845
rect 10376 19808 10421 19836
rect 10376 19796 10382 19808
rect 12161 19805 12173 19839
rect 12207 19836 12219 19839
rect 12342 19836 12348 19848
rect 12207 19808 12348 19836
rect 12207 19805 12219 19808
rect 12161 19799 12219 19805
rect 12342 19796 12348 19808
rect 12400 19796 12406 19848
rect 13832 19836 13860 19867
rect 14274 19864 14280 19916
rect 14332 19904 14338 19916
rect 14369 19907 14427 19913
rect 14369 19904 14381 19907
rect 14332 19876 14381 19904
rect 14332 19864 14338 19876
rect 14369 19873 14381 19876
rect 14415 19873 14427 19907
rect 14369 19867 14427 19873
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15565 19907 15623 19913
rect 15565 19904 15577 19907
rect 15252 19876 15577 19904
rect 15252 19864 15258 19876
rect 15565 19873 15577 19876
rect 15611 19873 15623 19907
rect 15565 19867 15623 19873
rect 16022 19864 16028 19916
rect 16080 19904 16086 19916
rect 16117 19907 16175 19913
rect 16117 19904 16129 19907
rect 16080 19876 16129 19904
rect 16080 19864 16086 19876
rect 16117 19873 16129 19876
rect 16163 19873 16175 19907
rect 16666 19904 16672 19916
rect 16627 19876 16672 19904
rect 16117 19867 16175 19873
rect 16666 19864 16672 19876
rect 16724 19864 16730 19916
rect 16850 19864 16856 19916
rect 16908 19904 16914 19916
rect 17221 19907 17279 19913
rect 17221 19904 17233 19907
rect 16908 19876 17233 19904
rect 16908 19864 16914 19876
rect 17221 19873 17233 19876
rect 17267 19873 17279 19907
rect 17221 19867 17279 19873
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18782 19904 18788 19916
rect 18371 19876 18788 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 18782 19864 18788 19876
rect 18840 19864 18846 19916
rect 18877 19907 18935 19913
rect 18877 19873 18889 19907
rect 18923 19904 18935 19907
rect 19150 19904 19156 19916
rect 18923 19876 19156 19904
rect 18923 19873 18935 19876
rect 18877 19867 18935 19873
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 19426 19904 19432 19916
rect 19387 19876 19432 19904
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 19981 19907 20039 19913
rect 19981 19873 19993 19907
rect 20027 19873 20039 19907
rect 20530 19904 20536 19916
rect 20491 19876 20536 19904
rect 19981 19867 20039 19873
rect 16482 19836 16488 19848
rect 13832 19808 16488 19836
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 19996 19836 20024 19867
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 20898 19836 20904 19848
rect 19996 19808 20904 19836
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 16301 19771 16359 19777
rect 16301 19737 16313 19771
rect 16347 19768 16359 19771
rect 18598 19768 18604 19780
rect 16347 19740 18604 19768
rect 16347 19737 16359 19740
rect 16301 19731 16359 19737
rect 18598 19728 18604 19740
rect 18656 19728 18662 19780
rect 8662 19700 8668 19712
rect 8623 19672 8668 19700
rect 8662 19660 8668 19672
rect 8720 19660 8726 19712
rect 9766 19700 9772 19712
rect 9727 19672 9772 19700
rect 9766 19660 9772 19672
rect 9824 19660 9830 19712
rect 11517 19703 11575 19709
rect 11517 19669 11529 19703
rect 11563 19700 11575 19703
rect 11882 19700 11888 19712
rect 11563 19672 11888 19700
rect 11563 19669 11575 19672
rect 11517 19663 11575 19669
rect 11882 19660 11888 19672
rect 11940 19660 11946 19712
rect 14001 19703 14059 19709
rect 14001 19669 14013 19703
rect 14047 19700 14059 19703
rect 18506 19700 18512 19712
rect 14047 19672 18512 19700
rect 14047 19669 14059 19672
rect 14001 19663 14059 19669
rect 18506 19660 18512 19672
rect 18564 19660 18570 19712
rect 20165 19703 20223 19709
rect 20165 19669 20177 19703
rect 20211 19700 20223 19703
rect 20254 19700 20260 19712
rect 20211 19672 20260 19700
rect 20211 19669 20223 19672
rect 20165 19663 20223 19669
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 20622 19660 20628 19712
rect 20680 19700 20686 19712
rect 20717 19703 20775 19709
rect 20717 19700 20729 19703
rect 20680 19672 20729 19700
rect 20680 19660 20686 19672
rect 20717 19669 20729 19672
rect 20763 19669 20775 19703
rect 20717 19663 20775 19669
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 10226 19456 10232 19508
rect 10284 19496 10290 19508
rect 17770 19496 17776 19508
rect 10284 19468 17776 19496
rect 10284 19456 10290 19468
rect 17770 19456 17776 19468
rect 17828 19456 17834 19508
rect 18966 19456 18972 19508
rect 19024 19496 19030 19508
rect 19061 19499 19119 19505
rect 19061 19496 19073 19499
rect 19024 19468 19073 19496
rect 19024 19456 19030 19468
rect 19061 19465 19073 19468
rect 19107 19465 19119 19499
rect 19061 19459 19119 19465
rect 9968 19332 10180 19360
rect 8386 19292 8392 19304
rect 8347 19264 8392 19292
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 8478 19252 8484 19304
rect 8536 19292 8542 19304
rect 9968 19292 9996 19332
rect 8536 19264 9996 19292
rect 10045 19295 10103 19301
rect 8536 19252 8542 19264
rect 10045 19261 10057 19295
rect 10091 19261 10103 19295
rect 10152 19292 10180 19332
rect 12360 19332 12572 19360
rect 10152 19264 10456 19292
rect 10045 19255 10103 19261
rect 8656 19227 8714 19233
rect 8656 19193 8668 19227
rect 8702 19224 8714 19227
rect 9214 19224 9220 19236
rect 8702 19196 9220 19224
rect 8702 19193 8714 19196
rect 8656 19187 8714 19193
rect 9214 19184 9220 19196
rect 9272 19184 9278 19236
rect 9950 19184 9956 19236
rect 10008 19224 10014 19236
rect 10060 19224 10088 19255
rect 10008 19196 10088 19224
rect 10008 19184 10014 19196
rect 10226 19184 10232 19236
rect 10284 19233 10290 19236
rect 10284 19227 10348 19233
rect 10284 19193 10302 19227
rect 10336 19193 10348 19227
rect 10428 19224 10456 19264
rect 11698 19252 11704 19304
rect 11756 19292 11762 19304
rect 11756 19264 11801 19292
rect 11756 19252 11762 19264
rect 12360 19224 12388 19332
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19261 12495 19295
rect 12437 19255 12495 19261
rect 10428 19196 12388 19224
rect 10284 19187 10348 19193
rect 10284 19184 10290 19187
rect 12452 19168 12480 19255
rect 12544 19168 12572 19332
rect 14090 19292 14096 19304
rect 14051 19264 14096 19292
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 14182 19252 14188 19304
rect 14240 19292 14246 19304
rect 14240 19264 14504 19292
rect 14240 19252 14246 19264
rect 12618 19184 12624 19236
rect 12676 19233 12682 19236
rect 12676 19227 12740 19233
rect 12676 19193 12694 19227
rect 12728 19193 12740 19227
rect 12676 19187 12740 19193
rect 12676 19184 12682 19187
rect 13630 19184 13636 19236
rect 13688 19224 13694 19236
rect 13688 19196 14320 19224
rect 13688 19184 13694 19196
rect 2498 19116 2504 19168
rect 2556 19156 2562 19168
rect 9582 19156 9588 19168
rect 2556 19128 9588 19156
rect 2556 19116 2562 19128
rect 9582 19116 9588 19128
rect 9640 19116 9646 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 9769 19159 9827 19165
rect 9769 19156 9781 19159
rect 9732 19128 9781 19156
rect 9732 19116 9738 19128
rect 9769 19125 9781 19128
rect 9815 19125 9827 19159
rect 11422 19156 11428 19168
rect 11383 19128 11428 19156
rect 9769 19119 9827 19125
rect 11422 19116 11428 19128
rect 11480 19116 11486 19168
rect 11885 19159 11943 19165
rect 11885 19125 11897 19159
rect 11931 19156 11943 19159
rect 11974 19156 11980 19168
rect 11931 19128 11980 19156
rect 11931 19125 11943 19128
rect 11885 19119 11943 19125
rect 11974 19116 11980 19128
rect 12032 19116 12038 19168
rect 12434 19116 12440 19168
rect 12492 19116 12498 19168
rect 12526 19116 12532 19168
rect 12584 19116 12590 19168
rect 12894 19116 12900 19168
rect 12952 19156 12958 19168
rect 13538 19156 13544 19168
rect 12952 19128 13544 19156
rect 12952 19116 12958 19128
rect 13538 19116 13544 19128
rect 13596 19156 13602 19168
rect 14292 19165 14320 19196
rect 13817 19159 13875 19165
rect 13817 19156 13829 19159
rect 13596 19128 13829 19156
rect 13596 19116 13602 19128
rect 13817 19125 13829 19128
rect 13863 19125 13875 19159
rect 13817 19119 13875 19125
rect 14277 19159 14335 19165
rect 14277 19125 14289 19159
rect 14323 19125 14335 19159
rect 14476 19156 14504 19264
rect 14550 19252 14556 19304
rect 14608 19292 14614 19304
rect 14645 19295 14703 19301
rect 14645 19292 14657 19295
rect 14608 19264 14657 19292
rect 14608 19252 14614 19264
rect 14645 19261 14657 19264
rect 14691 19261 14703 19295
rect 14645 19255 14703 19261
rect 15197 19295 15255 19301
rect 15197 19261 15209 19295
rect 15243 19292 15255 19295
rect 15470 19292 15476 19304
rect 15243 19264 15476 19292
rect 15243 19261 15255 19264
rect 15197 19255 15255 19261
rect 15470 19252 15476 19264
rect 15528 19252 15534 19304
rect 15562 19252 15568 19304
rect 15620 19292 15626 19304
rect 15749 19295 15807 19301
rect 15749 19292 15761 19295
rect 15620 19264 15761 19292
rect 15620 19252 15626 19264
rect 15749 19261 15761 19264
rect 15795 19261 15807 19295
rect 15749 19255 15807 19261
rect 16485 19295 16543 19301
rect 16485 19261 16497 19295
rect 16531 19292 16543 19295
rect 16758 19292 16764 19304
rect 16531 19264 16764 19292
rect 16531 19261 16543 19264
rect 16485 19255 16543 19261
rect 16758 19252 16764 19264
rect 16816 19252 16822 19304
rect 17126 19292 17132 19304
rect 17087 19264 17132 19292
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 17405 19295 17463 19301
rect 17405 19261 17417 19295
rect 17451 19292 17463 19295
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17451 19264 18061 19292
rect 17451 19261 17463 19264
rect 17405 19255 17463 19261
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18877 19295 18935 19301
rect 18877 19292 18889 19295
rect 18049 19255 18107 19261
rect 18156 19264 18889 19292
rect 15286 19184 15292 19236
rect 15344 19224 15350 19236
rect 18156 19224 18184 19264
rect 18877 19261 18889 19264
rect 18923 19261 18935 19295
rect 18877 19255 18935 19261
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19429 19295 19487 19301
rect 19429 19292 19441 19295
rect 19392 19264 19441 19292
rect 19392 19252 19398 19264
rect 19429 19261 19441 19264
rect 19475 19261 19487 19295
rect 19978 19292 19984 19304
rect 19939 19264 19984 19292
rect 19429 19255 19487 19261
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 20346 19252 20352 19304
rect 20404 19292 20410 19304
rect 20533 19295 20591 19301
rect 20533 19292 20545 19295
rect 20404 19264 20545 19292
rect 20404 19252 20410 19264
rect 20533 19261 20545 19264
rect 20579 19261 20591 19295
rect 20533 19255 20591 19261
rect 15344 19196 18184 19224
rect 15344 19184 15350 19196
rect 18506 19184 18512 19236
rect 18564 19224 18570 19236
rect 21358 19224 21364 19236
rect 18564 19196 21364 19224
rect 18564 19184 18570 19196
rect 21358 19184 21364 19196
rect 21416 19184 21422 19236
rect 14829 19159 14887 19165
rect 14829 19156 14841 19159
rect 14476 19128 14841 19156
rect 14277 19119 14335 19125
rect 14829 19125 14841 19128
rect 14875 19125 14887 19159
rect 14829 19119 14887 19125
rect 15010 19116 15016 19168
rect 15068 19156 15074 19168
rect 15381 19159 15439 19165
rect 15381 19156 15393 19159
rect 15068 19128 15393 19156
rect 15068 19116 15074 19128
rect 15381 19125 15393 19128
rect 15427 19125 15439 19159
rect 15381 19119 15439 19125
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 15896 19128 15945 19156
rect 15896 19116 15902 19128
rect 15933 19125 15945 19128
rect 15979 19125 15991 19159
rect 15933 19119 15991 19125
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 16669 19159 16727 19165
rect 16669 19156 16681 19159
rect 16448 19128 16681 19156
rect 16448 19116 16454 19128
rect 16669 19125 16681 19128
rect 16715 19125 16727 19159
rect 16669 19119 16727 19125
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18690 19156 18696 19168
rect 18279 19128 18696 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 19242 19116 19248 19168
rect 19300 19156 19306 19168
rect 19613 19159 19671 19165
rect 19613 19156 19625 19159
rect 19300 19128 19625 19156
rect 19300 19116 19306 19128
rect 19613 19125 19625 19128
rect 19659 19125 19671 19159
rect 20162 19156 20168 19168
rect 20123 19128 20168 19156
rect 19613 19119 19671 19125
rect 20162 19116 20168 19128
rect 20220 19116 20226 19168
rect 20717 19159 20775 19165
rect 20717 19125 20729 19159
rect 20763 19156 20775 19159
rect 20806 19156 20812 19168
rect 20763 19128 20812 19156
rect 20763 19125 20775 19128
rect 20717 19119 20775 19125
rect 20806 19116 20812 19128
rect 20864 19116 20870 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 290 18912 296 18964
rect 348 18952 354 18964
rect 9033 18955 9091 18961
rect 348 18924 8984 18952
rect 348 18912 354 18924
rect 8386 18884 8392 18896
rect 7668 18856 8392 18884
rect 7374 18776 7380 18828
rect 7432 18816 7438 18828
rect 7668 18825 7696 18856
rect 8386 18844 8392 18856
rect 8444 18884 8450 18896
rect 8444 18856 8892 18884
rect 8444 18844 8450 18856
rect 7653 18819 7711 18825
rect 7653 18816 7665 18819
rect 7432 18788 7665 18816
rect 7432 18776 7438 18788
rect 7653 18785 7665 18788
rect 7699 18785 7711 18819
rect 7653 18779 7711 18785
rect 7920 18819 7978 18825
rect 7920 18785 7932 18819
rect 7966 18816 7978 18819
rect 8754 18816 8760 18828
rect 7966 18788 8760 18816
rect 7966 18785 7978 18788
rect 7920 18779 7978 18785
rect 8754 18776 8760 18788
rect 8812 18776 8818 18828
rect 1394 18708 1400 18760
rect 1452 18748 1458 18760
rect 1452 18720 6408 18748
rect 1452 18708 1458 18720
rect 4706 18572 4712 18624
rect 4764 18612 4770 18624
rect 6178 18612 6184 18624
rect 4764 18584 6184 18612
rect 4764 18572 4770 18584
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 6380 18612 6408 18720
rect 8864 18680 8892 18856
rect 8956 18748 8984 18924
rect 9033 18921 9045 18955
rect 9079 18952 9091 18955
rect 9214 18952 9220 18964
rect 9079 18924 9220 18952
rect 9079 18921 9091 18924
rect 9033 18915 9091 18921
rect 9214 18912 9220 18924
rect 9272 18912 9278 18964
rect 10134 18952 10140 18964
rect 10095 18924 10140 18952
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 11977 18955 12035 18961
rect 11977 18921 11989 18955
rect 12023 18952 12035 18955
rect 12342 18952 12348 18964
rect 12023 18924 12348 18952
rect 12023 18921 12035 18924
rect 11977 18915 12035 18921
rect 12342 18912 12348 18924
rect 12400 18912 12406 18964
rect 13630 18912 13636 18964
rect 13688 18952 13694 18964
rect 15562 18952 15568 18964
rect 13688 18924 15568 18952
rect 13688 18912 13694 18924
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 15657 18955 15715 18961
rect 15657 18921 15669 18955
rect 15703 18952 15715 18955
rect 20070 18952 20076 18964
rect 15703 18924 20076 18952
rect 15703 18921 15715 18924
rect 15657 18915 15715 18921
rect 20070 18912 20076 18924
rect 20128 18912 20134 18964
rect 9674 18844 9680 18896
rect 9732 18884 9738 18896
rect 10226 18884 10232 18896
rect 9732 18856 10232 18884
rect 9732 18844 9738 18856
rect 10226 18844 10232 18856
rect 10284 18844 10290 18896
rect 10502 18844 10508 18896
rect 10560 18884 10566 18896
rect 10864 18887 10922 18893
rect 10864 18884 10876 18887
rect 10560 18856 10876 18884
rect 10560 18844 10566 18856
rect 10864 18853 10876 18856
rect 10910 18884 10922 18887
rect 11422 18884 11428 18896
rect 10910 18856 11428 18884
rect 10910 18853 10922 18856
rect 10864 18847 10922 18853
rect 11422 18844 11428 18856
rect 11480 18844 11486 18896
rect 12894 18893 12900 18896
rect 12888 18884 12900 18893
rect 12855 18856 12900 18884
rect 12888 18847 12900 18856
rect 12894 18844 12900 18847
rect 12952 18844 12958 18896
rect 19150 18884 19156 18896
rect 19111 18856 19156 18884
rect 19150 18844 19156 18856
rect 19208 18844 19214 18896
rect 19426 18844 19432 18896
rect 19484 18884 19490 18896
rect 19889 18887 19947 18893
rect 19889 18884 19901 18887
rect 19484 18856 19901 18884
rect 19484 18844 19490 18856
rect 19889 18853 19901 18856
rect 19935 18853 19947 18887
rect 19889 18847 19947 18853
rect 9766 18776 9772 18828
rect 9824 18816 9830 18828
rect 10134 18816 10140 18828
rect 9824 18788 10140 18816
rect 9824 18776 9830 18788
rect 10134 18776 10140 18788
rect 10192 18776 10198 18828
rect 12434 18816 12440 18828
rect 10612 18788 12440 18816
rect 10226 18748 10232 18760
rect 8956 18720 10232 18748
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 10612 18757 10640 18788
rect 12434 18776 12440 18788
rect 12492 18816 12498 18828
rect 12621 18819 12679 18825
rect 12621 18816 12633 18819
rect 12492 18788 12633 18816
rect 12492 18776 12498 18788
rect 12621 18785 12633 18788
rect 12667 18785 12679 18819
rect 12621 18779 12679 18785
rect 14458 18776 14464 18828
rect 14516 18816 14522 18828
rect 14645 18819 14703 18825
rect 14645 18816 14657 18819
rect 14516 18788 14657 18816
rect 14516 18776 14522 18788
rect 14645 18785 14657 18788
rect 14691 18785 14703 18819
rect 14645 18779 14703 18785
rect 15473 18819 15531 18825
rect 15473 18785 15485 18819
rect 15519 18816 15531 18819
rect 15746 18816 15752 18828
rect 15519 18788 15752 18816
rect 15519 18785 15531 18788
rect 15473 18779 15531 18785
rect 15746 18776 15752 18788
rect 15804 18776 15810 18828
rect 16114 18776 16120 18828
rect 16172 18816 16178 18828
rect 16281 18819 16339 18825
rect 16281 18816 16293 18819
rect 16172 18788 16293 18816
rect 16172 18776 16178 18788
rect 16281 18785 16293 18788
rect 16327 18785 16339 18819
rect 16281 18779 16339 18785
rect 18049 18819 18107 18825
rect 18049 18785 18061 18819
rect 18095 18816 18107 18819
rect 18598 18816 18604 18828
rect 18095 18788 18604 18816
rect 18095 18785 18107 18788
rect 18049 18779 18107 18785
rect 18598 18776 18604 18788
rect 18656 18776 18662 18828
rect 18874 18816 18880 18828
rect 18835 18788 18880 18816
rect 18874 18776 18880 18788
rect 18932 18776 18938 18828
rect 19518 18776 19524 18828
rect 19576 18816 19582 18828
rect 19613 18819 19671 18825
rect 19613 18816 19625 18819
rect 19576 18788 19625 18816
rect 19576 18776 19582 18788
rect 19613 18785 19625 18788
rect 19659 18785 19671 18819
rect 19613 18779 19671 18785
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18717 10655 18751
rect 10597 18711 10655 18717
rect 9950 18680 9956 18692
rect 8864 18652 9956 18680
rect 9950 18640 9956 18652
rect 10008 18680 10014 18692
rect 10612 18680 10640 18711
rect 15378 18708 15384 18760
rect 15436 18748 15442 18760
rect 16025 18751 16083 18757
rect 16025 18748 16037 18751
rect 15436 18720 16037 18748
rect 15436 18708 15442 18720
rect 16025 18717 16037 18720
rect 16071 18717 16083 18751
rect 16025 18711 16083 18717
rect 17954 18708 17960 18760
rect 18012 18748 18018 18760
rect 18141 18751 18199 18757
rect 18141 18748 18153 18751
rect 18012 18720 18153 18748
rect 18012 18708 18018 18720
rect 18141 18717 18153 18720
rect 18187 18717 18199 18751
rect 18141 18711 18199 18717
rect 18325 18751 18383 18757
rect 18325 18717 18337 18751
rect 18371 18748 18383 18751
rect 18506 18748 18512 18760
rect 18371 18720 18512 18748
rect 18371 18717 18383 18720
rect 18325 18711 18383 18717
rect 18506 18708 18512 18720
rect 18564 18708 18570 18760
rect 19702 18680 19708 18692
rect 10008 18652 10640 18680
rect 17144 18652 19708 18680
rect 10008 18640 10014 18652
rect 11790 18612 11796 18624
rect 6380 18584 11796 18612
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 13998 18612 14004 18624
rect 13959 18584 14004 18612
rect 13998 18572 14004 18584
rect 14056 18572 14062 18624
rect 14829 18615 14887 18621
rect 14829 18581 14841 18615
rect 14875 18612 14887 18615
rect 17144 18612 17172 18652
rect 19702 18640 19708 18652
rect 19760 18640 19766 18692
rect 14875 18584 17172 18612
rect 14875 18581 14887 18584
rect 14829 18575 14887 18581
rect 17218 18572 17224 18624
rect 17276 18612 17282 18624
rect 17405 18615 17463 18621
rect 17405 18612 17417 18615
rect 17276 18584 17417 18612
rect 17276 18572 17282 18584
rect 17405 18581 17417 18584
rect 17451 18581 17463 18615
rect 17405 18575 17463 18581
rect 17681 18615 17739 18621
rect 17681 18581 17693 18615
rect 17727 18612 17739 18615
rect 19242 18612 19248 18624
rect 17727 18584 19248 18612
rect 17727 18581 17739 18584
rect 17681 18575 17739 18581
rect 19242 18572 19248 18584
rect 19300 18572 19306 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 8202 18368 8208 18420
rect 8260 18408 8266 18420
rect 12894 18408 12900 18420
rect 8260 18380 12900 18408
rect 8260 18368 8266 18380
rect 12894 18368 12900 18380
rect 12952 18368 12958 18420
rect 15286 18408 15292 18420
rect 13188 18380 15292 18408
rect 3050 18300 3056 18352
rect 3108 18340 3114 18352
rect 9861 18343 9919 18349
rect 3108 18312 9812 18340
rect 3108 18300 3114 18312
rect 8662 18232 8668 18284
rect 8720 18272 8726 18284
rect 9309 18275 9367 18281
rect 9309 18272 9321 18275
rect 8720 18244 9321 18272
rect 8720 18232 8726 18244
rect 9309 18241 9321 18244
rect 9355 18241 9367 18275
rect 9309 18235 9367 18241
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18272 9551 18275
rect 9674 18272 9680 18284
rect 9539 18244 9680 18272
rect 9539 18241 9551 18244
rect 9493 18235 9551 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 9784 18272 9812 18312
rect 9861 18309 9873 18343
rect 9907 18340 9919 18343
rect 11974 18340 11980 18352
rect 9907 18312 11980 18340
rect 9907 18309 9919 18312
rect 9861 18303 9919 18309
rect 11974 18300 11980 18312
rect 12032 18300 12038 18352
rect 10318 18272 10324 18284
rect 9784 18244 10324 18272
rect 10318 18232 10324 18244
rect 10376 18232 10382 18284
rect 10502 18272 10508 18284
rect 10463 18244 10508 18272
rect 10502 18232 10508 18244
rect 10560 18232 10566 18284
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 13188 18272 13216 18380
rect 15286 18368 15292 18380
rect 15344 18368 15350 18420
rect 15746 18368 15752 18420
rect 15804 18408 15810 18420
rect 17589 18411 17647 18417
rect 15804 18380 16528 18408
rect 15804 18368 15810 18380
rect 16500 18340 16528 18380
rect 17589 18377 17601 18411
rect 17635 18408 17647 18411
rect 17862 18408 17868 18420
rect 17635 18380 17868 18408
rect 17635 18377 17647 18380
rect 17589 18371 17647 18377
rect 17862 18368 17868 18380
rect 17920 18368 17926 18420
rect 17954 18368 17960 18420
rect 18012 18408 18018 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 18012 18380 18061 18408
rect 18012 18368 18018 18380
rect 18049 18377 18061 18380
rect 18095 18377 18107 18411
rect 18049 18371 18107 18377
rect 18138 18340 18144 18352
rect 16500 18312 18144 18340
rect 18138 18300 18144 18312
rect 18196 18300 18202 18352
rect 11563 18244 13216 18272
rect 13357 18275 13415 18281
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 13357 18241 13369 18275
rect 13403 18272 13415 18275
rect 13403 18244 13860 18272
rect 13403 18241 13415 18244
rect 13357 18235 13415 18241
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 4212 18176 9904 18204
rect 4212 18164 4218 18176
rect 3602 18096 3608 18148
rect 3660 18136 3666 18148
rect 8570 18136 8576 18148
rect 3660 18108 8576 18136
rect 3660 18096 3666 18108
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 8864 18108 9812 18136
rect 8864 18077 8892 18108
rect 9784 18080 9812 18108
rect 8849 18071 8907 18077
rect 8849 18037 8861 18071
rect 8895 18037 8907 18071
rect 8849 18031 8907 18037
rect 9217 18071 9275 18077
rect 9217 18037 9229 18071
rect 9263 18068 9275 18071
rect 9582 18068 9588 18080
rect 9263 18040 9588 18068
rect 9263 18037 9275 18040
rect 9217 18031 9275 18037
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 9766 18028 9772 18080
rect 9824 18028 9830 18080
rect 9876 18068 9904 18176
rect 10134 18164 10140 18216
rect 10192 18204 10198 18216
rect 10229 18207 10287 18213
rect 10229 18204 10241 18207
rect 10192 18176 10241 18204
rect 10192 18164 10198 18176
rect 10229 18173 10241 18176
rect 10275 18173 10287 18207
rect 10229 18167 10287 18173
rect 10686 18164 10692 18216
rect 10744 18204 10750 18216
rect 11241 18207 11299 18213
rect 11241 18204 11253 18207
rect 10744 18176 11253 18204
rect 10744 18164 10750 18176
rect 11241 18173 11253 18176
rect 11287 18173 11299 18207
rect 13722 18204 13728 18216
rect 13683 18176 13728 18204
rect 11241 18167 11299 18173
rect 13722 18164 13728 18176
rect 13780 18164 13786 18216
rect 13832 18204 13860 18244
rect 17218 18232 17224 18284
rect 17276 18272 17282 18284
rect 18601 18275 18659 18281
rect 18601 18272 18613 18275
rect 17276 18244 18613 18272
rect 17276 18232 17282 18244
rect 18601 18241 18613 18244
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 18966 18232 18972 18284
rect 19024 18272 19030 18284
rect 19150 18272 19156 18284
rect 19024 18244 19156 18272
rect 19024 18232 19030 18244
rect 19150 18232 19156 18244
rect 19208 18232 19214 18284
rect 13998 18213 14004 18216
rect 13992 18204 14004 18213
rect 13832 18176 14004 18204
rect 13992 18167 14004 18176
rect 13998 18164 14004 18167
rect 14056 18164 14062 18216
rect 15378 18204 15384 18216
rect 15028 18176 15384 18204
rect 13906 18136 13912 18148
rect 12728 18108 13912 18136
rect 9950 18068 9956 18080
rect 9876 18040 9956 18068
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 10042 18028 10048 18080
rect 10100 18068 10106 18080
rect 10321 18071 10379 18077
rect 10321 18068 10333 18071
rect 10100 18040 10333 18068
rect 10100 18028 10106 18040
rect 10321 18037 10333 18040
rect 10367 18037 10379 18071
rect 10321 18031 10379 18037
rect 10778 18028 10784 18080
rect 10836 18068 10842 18080
rect 12066 18068 12072 18080
rect 10836 18040 12072 18068
rect 10836 18028 10842 18040
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 12728 18077 12756 18108
rect 13906 18096 13912 18108
rect 13964 18096 13970 18148
rect 12713 18071 12771 18077
rect 12713 18037 12725 18071
rect 12759 18037 12771 18071
rect 13078 18068 13084 18080
rect 13039 18040 13084 18068
rect 12713 18031 12771 18037
rect 13078 18028 13084 18040
rect 13136 18028 13142 18080
rect 13170 18028 13176 18080
rect 13228 18068 13234 18080
rect 13228 18040 13273 18068
rect 13228 18028 13234 18040
rect 13722 18028 13728 18080
rect 13780 18068 13786 18080
rect 15028 18068 15056 18176
rect 15378 18164 15384 18176
rect 15436 18164 15442 18216
rect 17402 18204 17408 18216
rect 17363 18176 17408 18204
rect 17402 18164 17408 18176
rect 17460 18204 17466 18216
rect 17770 18204 17776 18216
rect 17460 18176 17776 18204
rect 17460 18164 17466 18176
rect 17770 18164 17776 18176
rect 17828 18164 17834 18216
rect 18046 18164 18052 18216
rect 18104 18204 18110 18216
rect 19245 18207 19303 18213
rect 19245 18204 19257 18207
rect 18104 18176 19257 18204
rect 18104 18164 18110 18176
rect 19245 18173 19257 18176
rect 19291 18173 19303 18207
rect 19794 18204 19800 18216
rect 19755 18176 19800 18204
rect 19245 18167 19303 18173
rect 19794 18164 19800 18176
rect 19852 18164 19858 18216
rect 19886 18164 19892 18216
rect 19944 18204 19950 18216
rect 20533 18207 20591 18213
rect 20533 18204 20545 18207
rect 19944 18176 20545 18204
rect 19944 18164 19950 18176
rect 20533 18173 20545 18176
rect 20579 18173 20591 18207
rect 20533 18167 20591 18173
rect 15626 18139 15684 18145
rect 15626 18136 15638 18139
rect 15120 18108 15638 18136
rect 15120 18077 15148 18108
rect 15626 18105 15638 18108
rect 15672 18136 15684 18139
rect 15930 18136 15936 18148
rect 15672 18108 15936 18136
rect 15672 18105 15684 18108
rect 15626 18099 15684 18105
rect 15930 18096 15936 18108
rect 15988 18096 15994 18148
rect 16298 18096 16304 18148
rect 16356 18136 16362 18148
rect 16356 18108 16896 18136
rect 16356 18096 16362 18108
rect 13780 18040 15056 18068
rect 15105 18071 15163 18077
rect 13780 18028 13786 18040
rect 15105 18037 15117 18071
rect 15151 18037 15163 18071
rect 15105 18031 15163 18037
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 16761 18071 16819 18077
rect 16761 18068 16773 18071
rect 16172 18040 16773 18068
rect 16172 18028 16178 18040
rect 16761 18037 16773 18040
rect 16807 18037 16819 18071
rect 16868 18068 16896 18108
rect 17954 18096 17960 18148
rect 18012 18136 18018 18148
rect 20073 18139 20131 18145
rect 20073 18136 20085 18139
rect 18012 18108 20085 18136
rect 18012 18096 18018 18108
rect 20073 18105 20085 18108
rect 20119 18105 20131 18139
rect 20073 18099 20131 18105
rect 18417 18071 18475 18077
rect 18417 18068 18429 18071
rect 16868 18040 18429 18068
rect 16761 18031 16819 18037
rect 18417 18037 18429 18040
rect 18463 18037 18475 18071
rect 18417 18031 18475 18037
rect 18509 18071 18567 18077
rect 18509 18037 18521 18071
rect 18555 18068 18567 18071
rect 18690 18068 18696 18080
rect 18555 18040 18696 18068
rect 18555 18037 18567 18040
rect 18509 18031 18567 18037
rect 18690 18028 18696 18040
rect 18748 18028 18754 18080
rect 19058 18028 19064 18080
rect 19116 18068 19122 18080
rect 19429 18071 19487 18077
rect 19429 18068 19441 18071
rect 19116 18040 19441 18068
rect 19116 18028 19122 18040
rect 19429 18037 19441 18040
rect 19475 18037 19487 18071
rect 20714 18068 20720 18080
rect 20675 18040 20720 18068
rect 19429 18031 19487 18037
rect 20714 18028 20720 18040
rect 20772 18028 20778 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 8754 17864 8760 17876
rect 8715 17836 8760 17864
rect 8754 17824 8760 17836
rect 8812 17824 8818 17876
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 10689 17867 10747 17873
rect 10689 17864 10701 17867
rect 9732 17836 10701 17864
rect 9732 17824 9738 17836
rect 10689 17833 10701 17836
rect 10735 17833 10747 17867
rect 10689 17827 10747 17833
rect 12989 17867 13047 17873
rect 12989 17833 13001 17867
rect 13035 17864 13047 17867
rect 13078 17864 13084 17876
rect 13035 17836 13084 17864
rect 13035 17833 13047 17836
rect 12989 17827 13047 17833
rect 13078 17824 13084 17836
rect 13136 17824 13142 17876
rect 18046 17864 18052 17876
rect 14844 17836 18052 17864
rect 842 17756 848 17808
rect 900 17796 906 17808
rect 13357 17799 13415 17805
rect 900 17768 11376 17796
rect 900 17756 906 17768
rect 7374 17728 7380 17740
rect 7335 17700 7380 17728
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 7644 17731 7702 17737
rect 7644 17697 7656 17731
rect 7690 17728 7702 17731
rect 8386 17728 8392 17740
rect 7690 17700 8392 17728
rect 7690 17697 7702 17700
rect 7644 17691 7702 17697
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 9950 17688 9956 17740
rect 10008 17728 10014 17740
rect 10597 17731 10655 17737
rect 10597 17728 10609 17731
rect 10008 17700 10609 17728
rect 10008 17688 10014 17700
rect 10597 17697 10609 17700
rect 10643 17697 10655 17731
rect 10597 17691 10655 17697
rect 11054 17688 11060 17740
rect 11112 17728 11118 17740
rect 11241 17731 11299 17737
rect 11241 17728 11253 17731
rect 11112 17700 11253 17728
rect 11112 17688 11118 17700
rect 11241 17697 11253 17700
rect 11287 17697 11299 17731
rect 11241 17691 11299 17697
rect 10870 17660 10876 17672
rect 10831 17632 10876 17660
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 10229 17527 10287 17533
rect 10229 17493 10241 17527
rect 10275 17524 10287 17527
rect 11146 17524 11152 17536
rect 10275 17496 11152 17524
rect 10275 17493 10287 17496
rect 10229 17487 10287 17493
rect 11146 17484 11152 17496
rect 11204 17484 11210 17536
rect 11348 17524 11376 17768
rect 13357 17765 13369 17799
rect 13403 17796 13415 17799
rect 14737 17799 14795 17805
rect 14737 17796 14749 17799
rect 13403 17768 14749 17796
rect 13403 17765 13415 17768
rect 13357 17759 13415 17765
rect 14737 17765 14749 17768
rect 14783 17765 14795 17799
rect 14737 17759 14795 17765
rect 11514 17728 11520 17740
rect 11475 17700 11520 17728
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 11974 17728 11980 17740
rect 11935 17700 11980 17728
rect 11974 17688 11980 17700
rect 12032 17688 12038 17740
rect 12253 17731 12311 17737
rect 12253 17697 12265 17731
rect 12299 17728 12311 17731
rect 12299 17700 13759 17728
rect 12299 17697 12311 17700
rect 12253 17691 12311 17697
rect 13354 17620 13360 17672
rect 13412 17660 13418 17672
rect 13449 17663 13507 17669
rect 13449 17660 13461 17663
rect 13412 17632 13461 17660
rect 13412 17620 13418 17632
rect 13449 17629 13461 17632
rect 13495 17629 13507 17663
rect 13449 17623 13507 17629
rect 13538 17620 13544 17672
rect 13596 17660 13602 17672
rect 13731 17660 13759 17700
rect 13906 17688 13912 17740
rect 13964 17728 13970 17740
rect 14001 17731 14059 17737
rect 14001 17728 14013 17731
rect 13964 17700 14013 17728
rect 13964 17688 13970 17700
rect 14001 17697 14013 17700
rect 14047 17697 14059 17731
rect 14001 17691 14059 17697
rect 14277 17731 14335 17737
rect 14277 17697 14289 17731
rect 14323 17728 14335 17731
rect 14844 17728 14872 17836
rect 18046 17824 18052 17836
rect 18104 17824 18110 17876
rect 18325 17867 18383 17873
rect 18325 17833 18337 17867
rect 18371 17864 18383 17867
rect 18414 17864 18420 17876
rect 18371 17836 18420 17864
rect 18371 17833 18383 17836
rect 18325 17827 18383 17833
rect 18414 17824 18420 17836
rect 18472 17824 18478 17876
rect 18598 17864 18604 17876
rect 18559 17836 18604 17864
rect 18598 17824 18604 17836
rect 18656 17824 18662 17876
rect 16485 17799 16543 17805
rect 16485 17765 16497 17799
rect 16531 17796 16543 17799
rect 18969 17799 19027 17805
rect 18969 17796 18981 17799
rect 16531 17768 18981 17796
rect 16531 17765 16543 17768
rect 16485 17759 16543 17765
rect 18969 17765 18981 17768
rect 19015 17765 19027 17799
rect 18969 17759 19027 17765
rect 19981 17799 20039 17805
rect 19981 17765 19993 17799
rect 20027 17796 20039 17799
rect 20530 17796 20536 17808
rect 20027 17768 20536 17796
rect 20027 17765 20039 17768
rect 19981 17759 20039 17765
rect 20530 17756 20536 17768
rect 20588 17756 20594 17808
rect 14323 17700 14872 17728
rect 14323 17697 14335 17700
rect 14277 17691 14335 17697
rect 15378 17688 15384 17740
rect 15436 17728 15442 17740
rect 17218 17737 17224 17740
rect 15841 17731 15899 17737
rect 15841 17728 15853 17731
rect 15436 17700 15853 17728
rect 15436 17688 15442 17700
rect 15841 17697 15853 17700
rect 15887 17697 15899 17731
rect 17212 17728 17224 17737
rect 17179 17700 17224 17728
rect 15841 17691 15899 17697
rect 17212 17691 17224 17700
rect 17276 17728 17282 17740
rect 17276 17700 19196 17728
rect 17218 17688 17224 17691
rect 17276 17688 17282 17700
rect 15562 17660 15568 17672
rect 13596 17632 13641 17660
rect 13731 17632 15568 17660
rect 13596 17620 13602 17632
rect 15562 17620 15568 17632
rect 15620 17620 15626 17672
rect 15654 17620 15660 17672
rect 15712 17660 15718 17672
rect 15933 17663 15991 17669
rect 15933 17660 15945 17663
rect 15712 17632 15945 17660
rect 15712 17620 15718 17632
rect 15933 17629 15945 17632
rect 15979 17629 15991 17663
rect 16114 17660 16120 17672
rect 16075 17632 16120 17660
rect 15933 17623 15991 17629
rect 16114 17620 16120 17632
rect 16172 17620 16178 17672
rect 16942 17660 16948 17672
rect 16903 17632 16948 17660
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 18138 17620 18144 17672
rect 18196 17660 18202 17672
rect 19168 17669 19196 17700
rect 19242 17688 19248 17740
rect 19300 17728 19306 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 19300 17700 19717 17728
rect 19300 17688 19306 17700
rect 19705 17697 19717 17700
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 19061 17663 19119 17669
rect 19061 17660 19073 17663
rect 18196 17632 19073 17660
rect 18196 17620 18202 17632
rect 19061 17629 19073 17632
rect 19107 17629 19119 17663
rect 19061 17623 19119 17629
rect 19153 17663 19211 17669
rect 19153 17629 19165 17663
rect 19199 17629 19211 17663
rect 19153 17623 19211 17629
rect 11606 17552 11612 17604
rect 11664 17592 11670 17604
rect 12250 17592 12256 17604
rect 11664 17564 12256 17592
rect 11664 17552 11670 17564
rect 12250 17552 12256 17564
rect 12308 17552 12314 17604
rect 12434 17552 12440 17604
rect 12492 17592 12498 17604
rect 16850 17592 16856 17604
rect 12492 17564 16856 17592
rect 12492 17552 12498 17564
rect 16850 17552 16856 17564
rect 16908 17552 16914 17604
rect 18598 17552 18604 17604
rect 18656 17592 18662 17604
rect 22462 17592 22468 17604
rect 18656 17564 22468 17592
rect 18656 17552 18662 17564
rect 22462 17552 22468 17564
rect 22520 17552 22526 17604
rect 14366 17524 14372 17536
rect 11348 17496 14372 17524
rect 14366 17484 14372 17496
rect 14424 17484 14430 17536
rect 15473 17527 15531 17533
rect 15473 17493 15485 17527
rect 15519 17524 15531 17527
rect 19794 17524 19800 17536
rect 15519 17496 19800 17524
rect 15519 17493 15531 17496
rect 15473 17487 15531 17493
rect 19794 17484 19800 17496
rect 19852 17484 19858 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 7374 17320 7380 17332
rect 7024 17292 7380 17320
rect 7024 17193 7052 17292
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 8386 17320 8392 17332
rect 8347 17292 8392 17320
rect 8386 17280 8392 17292
rect 8444 17280 8450 17332
rect 9306 17280 9312 17332
rect 9364 17320 9370 17332
rect 12434 17320 12440 17332
rect 9364 17292 12440 17320
rect 9364 17280 9370 17292
rect 12434 17280 12440 17292
rect 12492 17280 12498 17332
rect 12529 17323 12587 17329
rect 12529 17289 12541 17323
rect 12575 17320 12587 17323
rect 13170 17320 13176 17332
rect 12575 17292 13176 17320
rect 12575 17289 12587 17292
rect 12529 17283 12587 17289
rect 13170 17280 13176 17292
rect 13228 17280 13234 17332
rect 13354 17280 13360 17332
rect 13412 17320 13418 17332
rect 15194 17320 15200 17332
rect 13412 17292 15200 17320
rect 13412 17280 13418 17292
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 15378 17320 15384 17332
rect 15339 17292 15384 17320
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 15562 17280 15568 17332
rect 15620 17320 15626 17332
rect 20346 17320 20352 17332
rect 15620 17292 20352 17320
rect 15620 17280 15626 17292
rect 20346 17280 20352 17292
rect 20404 17280 20410 17332
rect 7009 17187 7067 17193
rect 7009 17153 7021 17187
rect 7055 17153 7067 17187
rect 8404 17184 8432 17280
rect 8754 17212 8760 17264
rect 8812 17252 8818 17264
rect 10689 17255 10747 17261
rect 8812 17224 10272 17252
rect 8812 17212 8818 17224
rect 8662 17184 8668 17196
rect 8404 17156 8668 17184
rect 7009 17147 7067 17153
rect 8662 17144 8668 17156
rect 8720 17184 8726 17196
rect 10244 17193 10272 17224
rect 10689 17221 10701 17255
rect 10735 17252 10747 17255
rect 11606 17252 11612 17264
rect 10735 17224 11612 17252
rect 10735 17221 10747 17224
rect 10689 17215 10747 17221
rect 11606 17212 11612 17224
rect 11664 17212 11670 17264
rect 12894 17212 12900 17264
rect 12952 17252 12958 17264
rect 16114 17252 16120 17264
rect 12952 17224 16120 17252
rect 12952 17212 12958 17224
rect 16114 17212 16120 17224
rect 16172 17212 16178 17264
rect 17037 17255 17095 17261
rect 17037 17221 17049 17255
rect 17083 17252 17095 17255
rect 17773 17255 17831 17261
rect 17773 17252 17785 17255
rect 17083 17224 17785 17252
rect 17083 17221 17095 17224
rect 17037 17215 17095 17221
rect 17773 17221 17785 17224
rect 17819 17221 17831 17255
rect 17773 17215 17831 17221
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 8720 17156 9229 17184
rect 8720 17144 8726 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 10229 17187 10287 17193
rect 10229 17153 10241 17187
rect 10275 17153 10287 17187
rect 11238 17184 11244 17196
rect 11199 17156 11244 17184
rect 10229 17147 10287 17153
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 11882 17144 11888 17196
rect 11940 17184 11946 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 11940 17156 13001 17184
rect 11940 17144 11946 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 13173 17187 13231 17193
rect 13173 17153 13185 17187
rect 13219 17184 13231 17187
rect 13538 17184 13544 17196
rect 13219 17156 13544 17184
rect 13219 17153 13231 17156
rect 13173 17147 13231 17153
rect 13538 17144 13544 17156
rect 13596 17144 13602 17196
rect 13906 17144 13912 17196
rect 13964 17184 13970 17196
rect 14093 17187 14151 17193
rect 14093 17184 14105 17187
rect 13964 17156 14105 17184
rect 13964 17144 13970 17156
rect 14093 17153 14105 17156
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 15746 17184 15752 17196
rect 15436 17156 15752 17184
rect 15436 17144 15442 17156
rect 15746 17144 15752 17156
rect 15804 17144 15810 17196
rect 15930 17184 15936 17196
rect 15891 17156 15936 17184
rect 15930 17144 15936 17156
rect 15988 17144 15994 17196
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 19978 17184 19984 17196
rect 17000 17156 18092 17184
rect 19939 17156 19984 17184
rect 17000 17144 17006 17156
rect 18064 17128 18092 17156
rect 19978 17144 19984 17156
rect 20036 17144 20042 17196
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17184 20867 17187
rect 20898 17184 20904 17196
rect 20855 17156 20904 17184
rect 20855 17153 20867 17156
rect 20809 17147 20867 17153
rect 20898 17144 20904 17156
rect 20956 17144 20962 17196
rect 11146 17116 11152 17128
rect 11107 17088 11152 17116
rect 11146 17076 11152 17088
rect 11204 17076 11210 17128
rect 13998 17076 14004 17128
rect 14056 17116 14062 17128
rect 14458 17116 14464 17128
rect 14056 17088 14464 17116
rect 14056 17076 14062 17088
rect 14458 17076 14464 17088
rect 14516 17116 14522 17128
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 14516 17088 15853 17116
rect 14516 17076 14522 17088
rect 15841 17085 15853 17088
rect 15887 17085 15899 17119
rect 15841 17079 15899 17085
rect 16853 17119 16911 17125
rect 16853 17085 16865 17119
rect 16899 17116 16911 17119
rect 17310 17116 17316 17128
rect 16899 17088 17316 17116
rect 16899 17085 16911 17088
rect 16853 17079 16911 17085
rect 17310 17076 17316 17088
rect 17368 17076 17374 17128
rect 17405 17119 17463 17125
rect 17405 17085 17417 17119
rect 17451 17116 17463 17119
rect 17954 17116 17960 17128
rect 17451 17088 17960 17116
rect 17451 17085 17463 17088
rect 17405 17079 17463 17085
rect 17954 17076 17960 17088
rect 18012 17076 18018 17128
rect 18046 17076 18052 17128
rect 18104 17116 18110 17128
rect 18598 17116 18604 17128
rect 18104 17088 18149 17116
rect 18248 17088 18604 17116
rect 18104 17076 18110 17088
rect 7276 17051 7334 17057
rect 7276 17017 7288 17051
rect 7322 17048 7334 17051
rect 7650 17048 7656 17060
rect 7322 17020 7656 17048
rect 7322 17017 7334 17020
rect 7276 17011 7334 17017
rect 7650 17008 7656 17020
rect 7708 17008 7714 17060
rect 10045 17051 10103 17057
rect 10045 17048 10057 17051
rect 8680 17020 10057 17048
rect 8680 16989 8708 17020
rect 10045 17017 10057 17020
rect 10091 17017 10103 17051
rect 10045 17011 10103 17017
rect 11885 17051 11943 17057
rect 11885 17017 11897 17051
rect 11931 17048 11943 17051
rect 13446 17048 13452 17060
rect 11931 17020 13452 17048
rect 11931 17017 11943 17020
rect 11885 17011 11943 17017
rect 13446 17008 13452 17020
rect 13504 17008 13510 17060
rect 13909 17051 13967 17057
rect 13909 17017 13921 17051
rect 13955 17048 13967 17051
rect 15286 17048 15292 17060
rect 13955 17020 15292 17048
rect 13955 17017 13967 17020
rect 13909 17011 13967 17017
rect 15286 17008 15292 17020
rect 15344 17008 15350 17060
rect 15749 17051 15807 17057
rect 15749 17017 15761 17051
rect 15795 17048 15807 17051
rect 16393 17051 16451 17057
rect 16393 17048 16405 17051
rect 15795 17020 16405 17048
rect 15795 17017 15807 17020
rect 15749 17011 15807 17017
rect 16393 17017 16405 17020
rect 16439 17017 16451 17051
rect 16393 17011 16451 17017
rect 17773 17051 17831 17057
rect 17773 17017 17785 17051
rect 17819 17048 17831 17051
rect 18248 17048 18276 17088
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 18690 17076 18696 17128
rect 18748 17116 18754 17128
rect 19797 17119 19855 17125
rect 19797 17116 19809 17119
rect 18748 17088 19809 17116
rect 18748 17076 18754 17088
rect 19797 17085 19809 17088
rect 19843 17085 19855 17119
rect 20530 17116 20536 17128
rect 20491 17088 20536 17116
rect 19797 17079 19855 17085
rect 20530 17076 20536 17088
rect 20588 17076 20594 17128
rect 17819 17020 18276 17048
rect 18316 17051 18374 17057
rect 17819 17017 17831 17020
rect 17773 17011 17831 17017
rect 18316 17017 18328 17051
rect 18362 17048 18374 17051
rect 18506 17048 18512 17060
rect 18362 17020 18512 17048
rect 18362 17017 18374 17020
rect 18316 17011 18374 17017
rect 18506 17008 18512 17020
rect 18564 17008 18570 17060
rect 20990 17048 20996 17060
rect 18616 17020 20996 17048
rect 8665 16983 8723 16989
rect 8665 16949 8677 16983
rect 8711 16949 8723 16983
rect 9030 16980 9036 16992
rect 8991 16952 9036 16980
rect 8665 16943 8723 16949
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 9125 16983 9183 16989
rect 9125 16949 9137 16983
rect 9171 16980 9183 16983
rect 9306 16980 9312 16992
rect 9171 16952 9312 16980
rect 9171 16949 9183 16952
rect 9125 16943 9183 16949
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 9674 16980 9680 16992
rect 9635 16952 9680 16980
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 10134 16980 10140 16992
rect 10095 16952 10140 16980
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 11054 16980 11060 16992
rect 11015 16952 11060 16980
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 12894 16980 12900 16992
rect 12855 16952 12900 16980
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 13538 16980 13544 16992
rect 13499 16952 13544 16980
rect 13538 16940 13544 16952
rect 13596 16940 13602 16992
rect 14001 16983 14059 16989
rect 14001 16949 14013 16983
rect 14047 16980 14059 16983
rect 16298 16980 16304 16992
rect 14047 16952 16304 16980
rect 14047 16949 14059 16952
rect 14001 16943 14059 16949
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 17218 16980 17224 16992
rect 16632 16952 17224 16980
rect 16632 16940 16638 16952
rect 17218 16940 17224 16952
rect 17276 16940 17282 16992
rect 17589 16983 17647 16989
rect 17589 16949 17601 16983
rect 17635 16980 17647 16983
rect 17954 16980 17960 16992
rect 17635 16952 17960 16980
rect 17635 16949 17647 16952
rect 17589 16943 17647 16949
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 18138 16940 18144 16992
rect 18196 16980 18202 16992
rect 18616 16980 18644 17020
rect 20990 17008 20996 17020
rect 21048 17008 21054 17060
rect 18196 16952 18644 16980
rect 19429 16983 19487 16989
rect 18196 16940 18202 16952
rect 19429 16949 19441 16983
rect 19475 16980 19487 16983
rect 19794 16980 19800 16992
rect 19475 16952 19800 16980
rect 19475 16949 19487 16952
rect 19429 16943 19487 16949
rect 19794 16940 19800 16952
rect 19852 16940 19858 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 7009 16779 7067 16785
rect 7009 16745 7021 16779
rect 7055 16776 7067 16779
rect 8573 16779 8631 16785
rect 8573 16776 8585 16779
rect 7055 16748 8585 16776
rect 7055 16745 7067 16748
rect 7009 16739 7067 16745
rect 8573 16745 8585 16748
rect 8619 16745 8631 16779
rect 8573 16739 8631 16745
rect 9030 16736 9036 16788
rect 9088 16776 9094 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 9088 16748 9137 16776
rect 9088 16736 9094 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9125 16739 9183 16745
rect 12437 16779 12495 16785
rect 12437 16745 12449 16779
rect 12483 16776 12495 16779
rect 13081 16779 13139 16785
rect 13081 16776 13093 16779
rect 12483 16748 13093 16776
rect 12483 16745 12495 16748
rect 12437 16739 12495 16745
rect 13081 16745 13093 16748
rect 13127 16745 13139 16779
rect 13446 16776 13452 16788
rect 13407 16748 13452 16776
rect 13081 16739 13139 16745
rect 13446 16736 13452 16748
rect 13504 16736 13510 16788
rect 14182 16776 14188 16788
rect 14143 16748 14188 16776
rect 14182 16736 14188 16748
rect 14240 16736 14246 16788
rect 14645 16779 14703 16785
rect 14645 16776 14657 16779
rect 14476 16748 14657 16776
rect 6914 16668 6920 16720
rect 6972 16708 6978 16720
rect 7377 16711 7435 16717
rect 7377 16708 7389 16711
rect 6972 16680 7389 16708
rect 6972 16668 6978 16680
rect 7377 16677 7389 16680
rect 7423 16677 7435 16711
rect 10134 16708 10140 16720
rect 7377 16671 7435 16677
rect 8128 16680 10140 16708
rect 5810 16600 5816 16652
rect 5868 16640 5874 16652
rect 6825 16643 6883 16649
rect 6825 16640 6837 16643
rect 5868 16612 6837 16640
rect 5868 16600 5874 16612
rect 6825 16609 6837 16612
rect 6871 16640 6883 16643
rect 7469 16643 7527 16649
rect 7469 16640 7481 16643
rect 6871 16612 7481 16640
rect 6871 16609 6883 16612
rect 6825 16603 6883 16609
rect 7469 16609 7481 16612
rect 7515 16640 7527 16643
rect 7558 16640 7564 16652
rect 7515 16612 7564 16640
rect 7515 16609 7527 16612
rect 7469 16603 7527 16609
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 7650 16572 7656 16584
rect 7611 16544 7656 16572
rect 7650 16532 7656 16544
rect 7708 16532 7714 16584
rect 8128 16513 8156 16680
rect 10134 16668 10140 16680
rect 10192 16668 10198 16720
rect 10870 16668 10876 16720
rect 10928 16668 10934 16720
rect 12529 16711 12587 16717
rect 12529 16677 12541 16711
rect 12575 16708 12587 16711
rect 13538 16708 13544 16720
rect 12575 16680 13544 16708
rect 12575 16677 12587 16680
rect 12529 16671 12587 16677
rect 13538 16668 13544 16680
rect 13596 16668 13602 16720
rect 14366 16668 14372 16720
rect 14424 16708 14430 16720
rect 14476 16708 14504 16748
rect 14645 16745 14657 16748
rect 14691 16745 14703 16779
rect 14645 16739 14703 16745
rect 16577 16779 16635 16785
rect 16577 16745 16589 16779
rect 16623 16776 16635 16779
rect 18138 16776 18144 16788
rect 16623 16748 18144 16776
rect 16623 16745 16635 16748
rect 16577 16739 16635 16745
rect 18138 16736 18144 16748
rect 18196 16736 18202 16788
rect 18233 16779 18291 16785
rect 18233 16745 18245 16779
rect 18279 16776 18291 16779
rect 18506 16776 18512 16788
rect 18279 16748 18512 16776
rect 18279 16745 18291 16748
rect 18233 16739 18291 16745
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 18601 16779 18659 16785
rect 18601 16745 18613 16779
rect 18647 16776 18659 16779
rect 19245 16779 19303 16785
rect 19245 16776 19257 16779
rect 18647 16748 19257 16776
rect 18647 16745 18659 16748
rect 18601 16739 18659 16745
rect 19245 16745 19257 16748
rect 19291 16745 19303 16779
rect 20990 16776 20996 16788
rect 19245 16739 19303 16745
rect 19536 16748 20996 16776
rect 14424 16680 14504 16708
rect 14553 16711 14611 16717
rect 14424 16668 14430 16680
rect 14553 16677 14565 16711
rect 14599 16708 14611 16711
rect 14734 16708 14740 16720
rect 14599 16680 14740 16708
rect 14599 16677 14611 16680
rect 14553 16671 14611 16677
rect 14734 16668 14740 16680
rect 14792 16668 14798 16720
rect 15841 16711 15899 16717
rect 15841 16677 15853 16711
rect 15887 16708 15899 16711
rect 16114 16708 16120 16720
rect 15887 16680 16120 16708
rect 15887 16677 15899 16680
rect 15841 16671 15899 16677
rect 16114 16668 16120 16680
rect 16172 16668 16178 16720
rect 19536 16708 19564 16748
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 16408 16680 19564 16708
rect 19613 16711 19671 16717
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16640 8539 16643
rect 9122 16640 9128 16652
rect 8527 16612 9128 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 10321 16643 10379 16649
rect 10321 16609 10333 16643
rect 10367 16640 10379 16643
rect 10502 16640 10508 16652
rect 10367 16612 10508 16640
rect 10367 16609 10379 16612
rect 10321 16603 10379 16609
rect 10502 16600 10508 16612
rect 10560 16600 10566 16652
rect 10680 16643 10738 16649
rect 10680 16609 10692 16643
rect 10726 16640 10738 16643
rect 10888 16640 10916 16668
rect 11790 16640 11796 16652
rect 10726 16612 11796 16640
rect 10726 16609 10738 16612
rect 10680 16603 10738 16609
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 16408 16649 16436 16680
rect 19613 16677 19625 16711
rect 19659 16708 19671 16711
rect 20901 16711 20959 16717
rect 20901 16708 20913 16711
rect 19659 16680 20913 16708
rect 19659 16677 19671 16680
rect 19613 16671 19671 16677
rect 20901 16677 20913 16680
rect 20947 16677 20959 16711
rect 20901 16671 20959 16677
rect 15749 16643 15807 16649
rect 15749 16609 15761 16643
rect 15795 16640 15807 16643
rect 16393 16643 16451 16649
rect 15795 16612 16344 16640
rect 15795 16609 15807 16612
rect 15749 16603 15807 16609
rect 8662 16572 8668 16584
rect 8623 16544 8668 16572
rect 8662 16532 8668 16544
rect 8720 16532 8726 16584
rect 10410 16572 10416 16584
rect 10371 16544 10416 16572
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 12621 16575 12679 16581
rect 12621 16572 12633 16575
rect 11808 16544 12633 16572
rect 8113 16507 8171 16513
rect 8113 16473 8125 16507
rect 8159 16473 8171 16507
rect 8113 16467 8171 16473
rect 7374 16396 7380 16448
rect 7432 16436 7438 16448
rect 9490 16436 9496 16448
rect 7432 16408 9496 16436
rect 7432 16396 7438 16408
rect 9490 16396 9496 16408
rect 9548 16436 9554 16448
rect 10137 16439 10195 16445
rect 10137 16436 10149 16439
rect 9548 16408 10149 16436
rect 9548 16396 9554 16408
rect 10137 16405 10149 16408
rect 10183 16436 10195 16439
rect 10410 16436 10416 16448
rect 10183 16408 10416 16436
rect 10183 16405 10195 16408
rect 10137 16399 10195 16405
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 11146 16396 11152 16448
rect 11204 16436 11210 16448
rect 11808 16445 11836 16544
rect 12621 16541 12633 16544
rect 12667 16541 12679 16575
rect 12621 16535 12679 16541
rect 12710 16532 12716 16584
rect 12768 16572 12774 16584
rect 13541 16575 13599 16581
rect 13541 16572 13553 16575
rect 12768 16544 13553 16572
rect 12768 16532 12774 16544
rect 13541 16541 13553 16544
rect 13587 16572 13599 16575
rect 13630 16572 13636 16584
rect 13587 16544 13636 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 13725 16575 13783 16581
rect 13725 16541 13737 16575
rect 13771 16572 13783 16575
rect 13906 16572 13912 16584
rect 13771 16544 13912 16572
rect 13771 16541 13783 16544
rect 13725 16535 13783 16541
rect 13906 16532 13912 16544
rect 13964 16532 13970 16584
rect 14829 16575 14887 16581
rect 14829 16541 14841 16575
rect 14875 16572 14887 16575
rect 15194 16572 15200 16584
rect 14875 16544 15200 16572
rect 14875 16541 14887 16544
rect 14829 16535 14887 16541
rect 15194 16532 15200 16544
rect 15252 16532 15258 16584
rect 15930 16532 15936 16584
rect 15988 16572 15994 16584
rect 16316 16572 16344 16612
rect 16393 16609 16405 16643
rect 16439 16609 16451 16643
rect 16574 16640 16580 16652
rect 16393 16603 16451 16609
rect 16500 16612 16580 16640
rect 16500 16572 16528 16612
rect 16574 16600 16580 16612
rect 16632 16600 16638 16652
rect 16942 16640 16948 16652
rect 16903 16612 16948 16640
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 17034 16600 17040 16652
rect 17092 16640 17098 16652
rect 17497 16643 17555 16649
rect 17497 16640 17509 16643
rect 17092 16612 17509 16640
rect 17092 16600 17098 16612
rect 17497 16609 17509 16612
rect 17543 16609 17555 16643
rect 17497 16603 17555 16609
rect 17773 16643 17831 16649
rect 17773 16609 17785 16643
rect 17819 16640 17831 16643
rect 18506 16640 18512 16652
rect 17819 16612 18512 16640
rect 17819 16609 17831 16612
rect 17773 16603 17831 16609
rect 18506 16600 18512 16612
rect 18564 16600 18570 16652
rect 18693 16643 18751 16649
rect 18693 16609 18705 16643
rect 18739 16640 18751 16643
rect 19150 16640 19156 16652
rect 18739 16612 19156 16640
rect 18739 16609 18751 16612
rect 18693 16603 18751 16609
rect 19150 16600 19156 16612
rect 19208 16600 19214 16652
rect 20257 16643 20315 16649
rect 20257 16640 20269 16643
rect 19536 16612 20269 16640
rect 15988 16544 16033 16572
rect 16316 16544 16528 16572
rect 18877 16575 18935 16581
rect 15988 16532 15994 16544
rect 18877 16541 18889 16575
rect 18923 16572 18935 16575
rect 19426 16572 19432 16584
rect 18923 16544 19432 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 19426 16532 19432 16544
rect 19484 16532 19490 16584
rect 15381 16507 15439 16513
rect 15381 16473 15393 16507
rect 15427 16504 15439 16507
rect 15654 16504 15660 16516
rect 15427 16476 15660 16504
rect 15427 16473 15439 16476
rect 15381 16467 15439 16473
rect 15654 16464 15660 16476
rect 15712 16464 15718 16516
rect 17586 16464 17592 16516
rect 17644 16504 17650 16516
rect 19536 16504 19564 16612
rect 20257 16609 20269 16612
rect 20303 16609 20315 16643
rect 21910 16640 21916 16652
rect 20257 16603 20315 16609
rect 20364 16612 21916 16640
rect 19702 16572 19708 16584
rect 19663 16544 19708 16572
rect 19702 16532 19708 16544
rect 19760 16532 19766 16584
rect 19794 16532 19800 16584
rect 19852 16572 19858 16584
rect 19852 16544 19897 16572
rect 19852 16532 19858 16544
rect 20364 16504 20392 16612
rect 21910 16600 21916 16612
rect 21968 16600 21974 16652
rect 17644 16476 19564 16504
rect 19904 16476 20392 16504
rect 17644 16464 17650 16476
rect 11793 16439 11851 16445
rect 11793 16436 11805 16439
rect 11204 16408 11805 16436
rect 11204 16396 11210 16408
rect 11793 16405 11805 16408
rect 11839 16405 11851 16439
rect 12066 16436 12072 16448
rect 12027 16408 12072 16436
rect 11793 16399 11851 16405
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 12158 16396 12164 16448
rect 12216 16436 12222 16448
rect 16482 16436 16488 16448
rect 12216 16408 16488 16436
rect 12216 16396 12222 16408
rect 16482 16396 16488 16408
rect 16540 16396 16546 16448
rect 17129 16439 17187 16445
rect 17129 16405 17141 16439
rect 17175 16436 17187 16439
rect 19904 16436 19932 16476
rect 20438 16436 20444 16448
rect 17175 16408 19932 16436
rect 20399 16408 20444 16436
rect 17175 16405 17187 16408
rect 17129 16399 17187 16405
rect 20438 16396 20444 16408
rect 20496 16396 20502 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 9674 16232 9680 16244
rect 8680 16204 9680 16232
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 6914 16028 6920 16040
rect 6871 16000 6920 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 6914 15988 6920 16000
rect 6972 16028 6978 16040
rect 7374 16028 7380 16040
rect 6972 16000 7380 16028
rect 6972 15988 6978 16000
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 8680 16037 8708 16204
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 10410 16192 10416 16244
rect 10468 16232 10474 16244
rect 10468 16204 12480 16232
rect 10468 16192 10474 16204
rect 12158 16164 12164 16176
rect 10704 16136 12164 16164
rect 8941 16099 8999 16105
rect 8941 16065 8953 16099
rect 8987 16096 8999 16099
rect 8987 16068 9628 16096
rect 8987 16065 8999 16068
rect 8941 16059 8999 16065
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 15997 8723 16031
rect 9490 16028 9496 16040
rect 9451 16000 9496 16028
rect 8665 15991 8723 15997
rect 9490 15988 9496 16000
rect 9548 15988 9554 16040
rect 9600 16028 9628 16068
rect 10704 16028 10732 16136
rect 12158 16124 12164 16136
rect 12216 16124 12222 16176
rect 11606 16096 11612 16108
rect 11567 16068 11612 16096
rect 11606 16056 11612 16068
rect 11664 16056 11670 16108
rect 12452 16105 12480 16204
rect 13464 16204 16436 16232
rect 11701 16099 11759 16105
rect 11701 16065 11713 16099
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 12437 16099 12495 16105
rect 12437 16065 12449 16099
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 11146 16028 11152 16040
rect 9600 16000 10732 16028
rect 10796 16000 11152 16028
rect 7092 15963 7150 15969
rect 7092 15929 7104 15963
rect 7138 15960 7150 15963
rect 9760 15963 9818 15969
rect 7138 15932 9720 15960
rect 7138 15929 7150 15932
rect 7092 15923 7150 15929
rect 8202 15892 8208 15904
rect 8163 15864 8208 15892
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 9692 15892 9720 15932
rect 9760 15929 9772 15963
rect 9806 15960 9818 15963
rect 10796 15960 10824 16000
rect 11146 15988 11152 16000
rect 11204 15988 11210 16040
rect 11514 16028 11520 16040
rect 11475 16000 11520 16028
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 11707 15960 11735 16059
rect 13464 16028 13492 16204
rect 15286 16124 15292 16176
rect 15344 16164 15350 16176
rect 15930 16164 15936 16176
rect 15344 16136 15936 16164
rect 15344 16124 15350 16136
rect 15930 16124 15936 16136
rect 15988 16124 15994 16176
rect 16408 16164 16436 16204
rect 16482 16192 16488 16244
rect 16540 16232 16546 16244
rect 19426 16232 19432 16244
rect 16540 16204 19104 16232
rect 19387 16204 19432 16232
rect 16540 16192 16546 16204
rect 16761 16167 16819 16173
rect 16761 16164 16773 16167
rect 16408 16136 16773 16164
rect 16761 16133 16773 16136
rect 16807 16133 16819 16167
rect 16761 16127 16819 16133
rect 16850 16124 16856 16176
rect 16908 16164 16914 16176
rect 16908 16136 16953 16164
rect 16908 16124 16914 16136
rect 16114 16056 16120 16108
rect 16172 16096 16178 16108
rect 16485 16099 16543 16105
rect 16485 16096 16497 16099
rect 16172 16068 16497 16096
rect 16172 16056 16178 16068
rect 16485 16065 16497 16068
rect 16531 16096 16543 16099
rect 17494 16096 17500 16108
rect 16531 16068 17500 16096
rect 16531 16065 16543 16068
rect 16485 16059 16543 16065
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 19076 16096 19104 16204
rect 19426 16192 19432 16204
rect 19484 16192 19490 16244
rect 19150 16124 19156 16176
rect 19208 16164 19214 16176
rect 19705 16167 19763 16173
rect 19705 16164 19717 16167
rect 19208 16136 19717 16164
rect 19208 16124 19214 16136
rect 19705 16133 19717 16136
rect 19751 16133 19763 16167
rect 19705 16127 19763 16133
rect 19886 16096 19892 16108
rect 19076 16068 19892 16096
rect 19886 16056 19892 16068
rect 19944 16056 19950 16108
rect 20257 16099 20315 16105
rect 20257 16065 20269 16099
rect 20303 16065 20315 16099
rect 20257 16059 20315 16065
rect 9806 15932 10824 15960
rect 10888 15932 11735 15960
rect 12176 16000 13492 16028
rect 9806 15929 9818 15932
rect 9760 15923 9818 15929
rect 10888 15901 10916 15932
rect 10873 15895 10931 15901
rect 10873 15892 10885 15895
rect 9692 15864 10885 15892
rect 10873 15861 10885 15864
rect 10919 15861 10931 15895
rect 11146 15892 11152 15904
rect 11107 15864 11152 15892
rect 10873 15855 10931 15861
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 11238 15852 11244 15904
rect 11296 15892 11302 15904
rect 12176 15892 12204 16000
rect 13538 15988 13544 16040
rect 13596 16028 13602 16040
rect 13722 16028 13728 16040
rect 13596 16000 13728 16028
rect 13596 15988 13602 16000
rect 13722 15988 13728 16000
rect 13780 16028 13786 16040
rect 14182 16028 14188 16040
rect 13780 16000 14188 16028
rect 13780 15988 13786 16000
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 14452 16031 14510 16037
rect 14452 15997 14464 16031
rect 14498 16028 14510 16031
rect 15194 16028 15200 16040
rect 14498 16000 15200 16028
rect 14498 15997 14510 16000
rect 14452 15991 14510 15997
rect 15194 15988 15200 16000
rect 15252 16028 15258 16040
rect 16132 16028 16160 16056
rect 16298 16028 16304 16040
rect 15252 16000 16160 16028
rect 16259 16000 16304 16028
rect 15252 15988 15258 16000
rect 16298 15988 16304 16000
rect 16356 15988 16362 16040
rect 16574 15988 16580 16040
rect 16632 16028 16638 16040
rect 18046 16028 18052 16040
rect 16632 16000 18052 16028
rect 16632 15988 16638 16000
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 18316 16031 18374 16037
rect 18316 15997 18328 16031
rect 18362 16028 18374 16031
rect 19794 16028 19800 16040
rect 18362 16000 19800 16028
rect 18362 15997 18374 16000
rect 18316 15991 18374 15997
rect 19794 15988 19800 16000
rect 19852 16028 19858 16040
rect 20272 16028 20300 16059
rect 19852 16000 20300 16028
rect 20717 16031 20775 16037
rect 19852 15988 19858 16000
rect 20717 15997 20729 16031
rect 20763 16028 20775 16031
rect 20898 16028 20904 16040
rect 20763 16000 20904 16028
rect 20763 15997 20775 16000
rect 20717 15991 20775 15997
rect 20898 15988 20904 16000
rect 20956 15988 20962 16040
rect 12704 15963 12762 15969
rect 12704 15929 12716 15963
rect 12750 15960 12762 15963
rect 13078 15960 13084 15972
rect 12750 15932 13084 15960
rect 12750 15929 12762 15932
rect 12704 15923 12762 15929
rect 13078 15920 13084 15932
rect 13136 15920 13142 15972
rect 16761 15963 16819 15969
rect 13464 15932 14504 15960
rect 11296 15864 12204 15892
rect 11296 15852 11302 15864
rect 12342 15852 12348 15904
rect 12400 15892 12406 15904
rect 13464 15892 13492 15932
rect 14476 15904 14504 15932
rect 16761 15929 16773 15963
rect 16807 15960 16819 15963
rect 17313 15963 17371 15969
rect 17313 15960 17325 15963
rect 16807 15932 17325 15960
rect 16807 15929 16819 15932
rect 16761 15923 16819 15929
rect 17313 15929 17325 15932
rect 17359 15960 17371 15963
rect 17402 15960 17408 15972
rect 17359 15932 17408 15960
rect 17359 15929 17371 15932
rect 17313 15923 17371 15929
rect 17402 15920 17408 15932
rect 17460 15920 17466 15972
rect 17678 15920 17684 15972
rect 17736 15960 17742 15972
rect 20165 15963 20223 15969
rect 20165 15960 20177 15963
rect 17736 15932 20177 15960
rect 17736 15920 17742 15932
rect 20165 15929 20177 15932
rect 20211 15929 20223 15963
rect 20165 15923 20223 15929
rect 12400 15864 13492 15892
rect 13817 15895 13875 15901
rect 12400 15852 12406 15864
rect 13817 15861 13829 15895
rect 13863 15892 13875 15895
rect 13906 15892 13912 15904
rect 13863 15864 13912 15892
rect 13863 15861 13875 15864
rect 13817 15855 13875 15861
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 14458 15852 14464 15904
rect 14516 15852 14522 15904
rect 15562 15892 15568 15904
rect 15523 15864 15568 15892
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 15838 15892 15844 15904
rect 15799 15864 15844 15892
rect 15838 15852 15844 15864
rect 15896 15852 15902 15904
rect 15930 15852 15936 15904
rect 15988 15892 15994 15904
rect 16209 15895 16267 15901
rect 16209 15892 16221 15895
rect 15988 15864 16221 15892
rect 15988 15852 15994 15864
rect 16209 15861 16221 15864
rect 16255 15861 16267 15895
rect 16209 15855 16267 15861
rect 16482 15852 16488 15904
rect 16540 15892 16546 15904
rect 17221 15895 17279 15901
rect 17221 15892 17233 15895
rect 16540 15864 17233 15892
rect 16540 15852 16546 15864
rect 17221 15861 17233 15864
rect 17267 15861 17279 15895
rect 17221 15855 17279 15861
rect 19150 15852 19156 15904
rect 19208 15892 19214 15904
rect 20073 15895 20131 15901
rect 20073 15892 20085 15895
rect 19208 15864 20085 15892
rect 19208 15852 19214 15864
rect 20073 15861 20085 15864
rect 20119 15861 20131 15895
rect 20073 15855 20131 15861
rect 20622 15852 20628 15904
rect 20680 15892 20686 15904
rect 20901 15895 20959 15901
rect 20901 15892 20913 15895
rect 20680 15864 20913 15892
rect 20680 15852 20686 15864
rect 20901 15861 20913 15864
rect 20947 15861 20959 15895
rect 20901 15855 20959 15861
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 7650 15648 7656 15700
rect 7708 15688 7714 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7708 15660 7849 15688
rect 7708 15648 7714 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 10689 15691 10747 15697
rect 10689 15657 10701 15691
rect 10735 15688 10747 15691
rect 11054 15688 11060 15700
rect 10735 15660 11060 15688
rect 10735 15657 10747 15660
rect 10689 15651 10747 15657
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 13906 15688 13912 15700
rect 13740 15660 13912 15688
rect 6914 15620 6920 15632
rect 6472 15592 6920 15620
rect 6472 15561 6500 15592
rect 6914 15580 6920 15592
rect 6972 15580 6978 15632
rect 9122 15580 9128 15632
rect 9180 15620 9186 15632
rect 11149 15623 11207 15629
rect 11149 15620 11161 15623
rect 9180 15592 11161 15620
rect 9180 15580 9186 15592
rect 11149 15589 11161 15592
rect 11195 15620 11207 15623
rect 11238 15620 11244 15632
rect 11195 15592 11244 15620
rect 11195 15589 11207 15592
rect 11149 15583 11207 15589
rect 11238 15580 11244 15592
rect 11296 15580 11302 15632
rect 11790 15580 11796 15632
rect 11848 15620 11854 15632
rect 13740 15620 13768 15660
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 14182 15648 14188 15700
rect 14240 15688 14246 15700
rect 15013 15691 15071 15697
rect 15013 15688 15025 15691
rect 14240 15660 15025 15688
rect 14240 15648 14246 15660
rect 15013 15657 15025 15660
rect 15059 15657 15071 15691
rect 15013 15651 15071 15657
rect 15657 15691 15715 15697
rect 15657 15657 15669 15691
rect 15703 15688 15715 15691
rect 16850 15688 16856 15700
rect 15703 15660 16856 15688
rect 15703 15657 15715 15660
rect 15657 15651 15715 15657
rect 16850 15648 16856 15660
rect 16908 15648 16914 15700
rect 17494 15648 17500 15700
rect 17552 15688 17558 15700
rect 17957 15691 18015 15697
rect 17957 15688 17969 15691
rect 17552 15660 17969 15688
rect 17552 15648 17558 15660
rect 17957 15657 17969 15660
rect 18003 15657 18015 15691
rect 17957 15651 18015 15657
rect 11848 15592 13768 15620
rect 13808 15623 13866 15629
rect 11848 15580 11854 15592
rect 13808 15589 13820 15623
rect 13854 15620 13866 15623
rect 15562 15620 15568 15632
rect 13854 15592 15568 15620
rect 13854 15589 13866 15592
rect 13808 15583 13866 15589
rect 15562 15580 15568 15592
rect 15620 15580 15626 15632
rect 15746 15620 15752 15632
rect 15707 15592 15752 15620
rect 15746 15580 15752 15592
rect 15804 15580 15810 15632
rect 18684 15623 18742 15629
rect 16316 15592 18644 15620
rect 6457 15555 6515 15561
rect 6457 15521 6469 15555
rect 6503 15521 6515 15555
rect 6457 15515 6515 15521
rect 6724 15555 6782 15561
rect 6724 15521 6736 15555
rect 6770 15552 6782 15555
rect 8110 15552 8116 15564
rect 6770 15524 8116 15552
rect 6770 15521 6782 15524
rect 6724 15515 6782 15521
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 9674 15552 9680 15564
rect 9635 15524 9680 15552
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15552 10011 15555
rect 10042 15552 10048 15564
rect 9999 15524 10048 15552
rect 9999 15521 10011 15524
rect 9953 15515 10011 15521
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15521 11115 15555
rect 11057 15515 11115 15521
rect 11072 15416 11100 15515
rect 11333 15487 11391 15493
rect 11333 15453 11345 15487
rect 11379 15484 11391 15487
rect 11808 15484 11836 15580
rect 12069 15555 12127 15561
rect 12069 15521 12081 15555
rect 12115 15552 12127 15555
rect 12434 15552 12440 15564
rect 12115 15524 12440 15552
rect 12115 15521 12127 15524
rect 12069 15515 12127 15521
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 12802 15552 12808 15564
rect 12763 15524 12808 15552
rect 12802 15512 12808 15524
rect 12860 15512 12866 15564
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15552 13139 15555
rect 16316 15552 16344 15592
rect 16482 15552 16488 15564
rect 13127 15524 16344 15552
rect 16443 15524 16488 15552
rect 13127 15521 13139 15524
rect 13081 15515 13139 15521
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 16844 15555 16902 15561
rect 16844 15521 16856 15555
rect 16890 15552 16902 15555
rect 17678 15552 17684 15564
rect 16890 15524 17684 15552
rect 16890 15521 16902 15524
rect 16844 15515 16902 15521
rect 17678 15512 17684 15524
rect 17736 15512 17742 15564
rect 18046 15512 18052 15564
rect 18104 15552 18110 15564
rect 18417 15555 18475 15561
rect 18417 15552 18429 15555
rect 18104 15524 18429 15552
rect 18104 15512 18110 15524
rect 18417 15521 18429 15524
rect 18463 15521 18475 15555
rect 18616 15552 18644 15592
rect 18684 15589 18696 15623
rect 18730 15620 18742 15623
rect 19426 15620 19432 15632
rect 18730 15592 19432 15620
rect 18730 15589 18742 15592
rect 18684 15583 18742 15589
rect 19426 15580 19432 15592
rect 19484 15580 19490 15632
rect 20070 15552 20076 15564
rect 18616 15524 19932 15552
rect 20031 15524 20076 15552
rect 18417 15515 18475 15521
rect 11379 15456 11836 15484
rect 11379 15453 11391 15456
rect 11333 15447 11391 15453
rect 11882 15444 11888 15496
rect 11940 15484 11946 15496
rect 12161 15487 12219 15493
rect 12161 15484 12173 15487
rect 11940 15456 12173 15484
rect 11940 15444 11946 15456
rect 12161 15453 12173 15456
rect 12207 15453 12219 15487
rect 12161 15447 12219 15453
rect 12342 15444 12348 15496
rect 12400 15484 12406 15496
rect 13538 15484 13544 15496
rect 12400 15456 13124 15484
rect 13499 15456 13544 15484
rect 12400 15444 12406 15456
rect 12894 15416 12900 15428
rect 11072 15388 12900 15416
rect 12894 15376 12900 15388
rect 12952 15376 12958 15428
rect 11698 15348 11704 15360
rect 11659 15320 11704 15348
rect 11698 15308 11704 15320
rect 11756 15308 11762 15360
rect 13096 15348 13124 15456
rect 13538 15444 13544 15456
rect 13596 15444 13602 15496
rect 15562 15444 15568 15496
rect 15620 15484 15626 15496
rect 15841 15487 15899 15493
rect 15841 15484 15853 15487
rect 15620 15456 15853 15484
rect 15620 15444 15626 15456
rect 15841 15453 15853 15456
rect 15887 15453 15899 15487
rect 15841 15447 15899 15453
rect 16209 15487 16267 15493
rect 16209 15453 16221 15487
rect 16255 15484 16267 15487
rect 16574 15484 16580 15496
rect 16255 15456 16580 15484
rect 16255 15453 16267 15456
rect 16209 15447 16267 15453
rect 16574 15444 16580 15456
rect 16632 15444 16638 15496
rect 15289 15419 15347 15425
rect 15289 15385 15301 15419
rect 15335 15416 15347 15419
rect 19904 15416 19932 15524
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 20254 15484 20260 15496
rect 20215 15456 20260 15484
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 20714 15416 20720 15428
rect 15335 15388 16611 15416
rect 19904 15388 20720 15416
rect 15335 15385 15347 15388
rect 15289 15379 15347 15385
rect 13722 15348 13728 15360
rect 13096 15320 13728 15348
rect 13722 15308 13728 15320
rect 13780 15308 13786 15360
rect 14918 15348 14924 15360
rect 14879 15320 14924 15348
rect 14918 15308 14924 15320
rect 14976 15308 14982 15360
rect 15013 15351 15071 15357
rect 15013 15317 15025 15351
rect 15059 15348 15071 15351
rect 16209 15351 16267 15357
rect 16209 15348 16221 15351
rect 15059 15320 16221 15348
rect 15059 15317 15071 15320
rect 15013 15311 15071 15317
rect 16209 15317 16221 15320
rect 16255 15348 16267 15351
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 16255 15320 16313 15348
rect 16255 15317 16267 15320
rect 16209 15311 16267 15317
rect 16301 15317 16313 15320
rect 16347 15317 16359 15351
rect 16583 15348 16611 15388
rect 20714 15376 20720 15388
rect 20772 15376 20778 15428
rect 16850 15348 16856 15360
rect 16583 15320 16856 15348
rect 16301 15311 16359 15317
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 19794 15348 19800 15360
rect 19755 15320 19800 15348
rect 19794 15308 19800 15320
rect 19852 15308 19858 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 8110 15104 8116 15156
rect 8168 15144 8174 15156
rect 9125 15147 9183 15153
rect 9125 15144 9137 15147
rect 8168 15116 9137 15144
rect 8168 15104 8174 15116
rect 9125 15113 9137 15116
rect 9171 15113 9183 15147
rect 9125 15107 9183 15113
rect 9401 15147 9459 15153
rect 9401 15113 9413 15147
rect 9447 15144 9459 15147
rect 9674 15144 9680 15156
rect 9447 15116 9680 15144
rect 9447 15113 9459 15116
rect 9401 15107 9459 15113
rect 6178 15008 6184 15020
rect 6139 14980 6184 15008
rect 6178 14968 6184 14980
rect 6236 14968 6242 15020
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 15008 6423 15011
rect 6914 15008 6920 15020
rect 6411 14980 6920 15008
rect 6411 14977 6423 14980
rect 6365 14971 6423 14977
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 7374 14968 7380 15020
rect 7432 15008 7438 15020
rect 7745 15011 7803 15017
rect 7745 15008 7757 15011
rect 7432 14980 7757 15008
rect 7432 14968 7438 14980
rect 7745 14977 7757 14980
rect 7791 14977 7803 15011
rect 9140 15008 9168 15107
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 12437 15147 12495 15153
rect 12437 15113 12449 15147
rect 12483 15144 12495 15147
rect 12802 15144 12808 15156
rect 12483 15116 12808 15144
rect 12483 15113 12495 15116
rect 12437 15107 12495 15113
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 16209 15147 16267 15153
rect 16209 15144 16221 15147
rect 13648 15116 16221 15144
rect 13648 15076 13676 15116
rect 16209 15113 16221 15116
rect 16255 15113 16267 15147
rect 16209 15107 16267 15113
rect 16393 15147 16451 15153
rect 16393 15113 16405 15147
rect 16439 15144 16451 15147
rect 20070 15144 20076 15156
rect 16439 15116 20076 15144
rect 16439 15113 16451 15116
rect 16393 15107 16451 15113
rect 20070 15104 20076 15116
rect 20128 15104 20134 15156
rect 10888 15048 13676 15076
rect 10888 15017 10916 15048
rect 14918 15036 14924 15088
rect 14976 15076 14982 15088
rect 19429 15079 19487 15085
rect 14976 15048 17080 15076
rect 14976 15036 14982 15048
rect 9953 15011 10011 15017
rect 9953 15008 9965 15011
rect 9140 14980 9965 15008
rect 7745 14971 7803 14977
rect 9953 14977 9965 14980
rect 9999 14977 10011 15011
rect 9953 14971 10011 14977
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 11698 14968 11704 15020
rect 11756 15008 11762 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11756 14980 11805 15008
rect 11756 14968 11762 14980
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 11793 14971 11851 14977
rect 11977 15011 12035 15017
rect 11977 14977 11989 15011
rect 12023 15008 12035 15011
rect 12434 15008 12440 15020
rect 12023 14980 12440 15008
rect 12023 14977 12035 14980
rect 11977 14971 12035 14977
rect 12434 14968 12440 14980
rect 12492 14968 12498 15020
rect 13078 15008 13084 15020
rect 13039 14980 13084 15008
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 13538 14968 13544 15020
rect 13596 15008 13602 15020
rect 13633 15011 13691 15017
rect 13633 15008 13645 15011
rect 13596 14980 13645 15008
rect 13596 14968 13602 14980
rect 13633 14977 13645 14980
rect 13679 14977 13691 15011
rect 13633 14971 13691 14977
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 6086 14940 6092 14952
rect 5592 14912 6092 14940
rect 5592 14900 5598 14912
rect 6086 14900 6092 14912
rect 6144 14900 6150 14952
rect 10597 14943 10655 14949
rect 10597 14909 10609 14943
rect 10643 14940 10655 14943
rect 11146 14940 11152 14952
rect 10643 14912 11152 14940
rect 10643 14909 10655 14912
rect 10597 14903 10655 14909
rect 11146 14900 11152 14912
rect 11204 14900 11210 14952
rect 13900 14943 13958 14949
rect 13900 14909 13912 14943
rect 13946 14940 13958 14943
rect 14936 14940 14964 15036
rect 15470 14968 15476 15020
rect 15528 15008 15534 15020
rect 15841 15011 15899 15017
rect 15841 15008 15853 15011
rect 15528 14980 15853 15008
rect 15528 14968 15534 14980
rect 15841 14977 15853 14980
rect 15887 15008 15899 15011
rect 15930 15008 15936 15020
rect 15887 14980 15936 15008
rect 15887 14977 15899 14980
rect 15841 14971 15899 14977
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 16025 15011 16083 15017
rect 16025 14977 16037 15011
rect 16071 15008 16083 15011
rect 16114 15008 16120 15020
rect 16071 14980 16120 15008
rect 16071 14977 16083 14980
rect 16025 14971 16083 14977
rect 16114 14968 16120 14980
rect 16172 14968 16178 15020
rect 16850 14968 16856 15020
rect 16908 15008 16914 15020
rect 17052 15017 17080 15048
rect 19429 15045 19441 15079
rect 19475 15076 19487 15079
rect 20530 15076 20536 15088
rect 19475 15048 20536 15076
rect 19475 15045 19487 15048
rect 19429 15039 19487 15045
rect 20530 15036 20536 15048
rect 20588 15036 20594 15088
rect 17037 15011 17095 15017
rect 16908 14980 16953 15008
rect 16908 14968 16914 14980
rect 17037 14977 17049 15011
rect 17083 14977 17095 15011
rect 17037 14971 17095 14977
rect 17770 14968 17776 15020
rect 17828 15008 17834 15020
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 17828 14980 18889 15008
rect 17828 14968 17834 14980
rect 18877 14977 18889 14980
rect 18923 14977 18935 15011
rect 18877 14971 18935 14977
rect 19061 15011 19119 15017
rect 19061 14977 19073 15011
rect 19107 15008 19119 15011
rect 19794 15008 19800 15020
rect 19107 14980 19800 15008
rect 19107 14977 19119 14980
rect 19061 14971 19119 14977
rect 19794 14968 19800 14980
rect 19852 14968 19858 15020
rect 19978 15008 19984 15020
rect 19939 14980 19984 15008
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20717 15011 20775 15017
rect 20717 14977 20729 15011
rect 20763 15008 20775 15011
rect 20990 15008 20996 15020
rect 20763 14980 20996 15008
rect 20763 14977 20775 14980
rect 20717 14971 20775 14977
rect 20990 14968 20996 14980
rect 21048 14968 21054 15020
rect 13946 14912 14964 14940
rect 13946 14909 13958 14912
rect 13900 14903 13958 14909
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 16761 14943 16819 14949
rect 16761 14940 16773 14943
rect 15344 14912 16773 14940
rect 15344 14900 15350 14912
rect 16761 14909 16773 14912
rect 16807 14909 16819 14943
rect 16761 14903 16819 14909
rect 17512 14912 20024 14940
rect 8012 14875 8070 14881
rect 8012 14841 8024 14875
rect 8058 14872 8070 14875
rect 8294 14872 8300 14884
rect 8058 14844 8300 14872
rect 8058 14841 8070 14844
rect 8012 14835 8070 14841
rect 8294 14832 8300 14844
rect 8352 14832 8358 14884
rect 8570 14832 8576 14884
rect 8628 14872 8634 14884
rect 9861 14875 9919 14881
rect 9861 14872 9873 14875
rect 8628 14844 9873 14872
rect 8628 14832 8634 14844
rect 9861 14841 9873 14844
rect 9907 14841 9919 14875
rect 12897 14875 12955 14881
rect 12897 14872 12909 14875
rect 9861 14835 9919 14841
rect 11348 14844 12909 14872
rect 5721 14807 5779 14813
rect 5721 14773 5733 14807
rect 5767 14804 5779 14807
rect 9030 14804 9036 14816
rect 5767 14776 9036 14804
rect 5767 14773 5779 14776
rect 5721 14767 5779 14773
rect 9030 14764 9036 14776
rect 9088 14764 9094 14816
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 11348 14813 11376 14844
rect 12897 14841 12909 14844
rect 12943 14841 12955 14875
rect 12897 14835 12955 14841
rect 15749 14875 15807 14881
rect 15749 14841 15761 14875
rect 15795 14872 15807 14875
rect 17405 14875 17463 14881
rect 17405 14872 17417 14875
rect 15795 14844 17417 14872
rect 15795 14841 15807 14844
rect 15749 14835 15807 14841
rect 17405 14841 17417 14844
rect 17451 14841 17463 14875
rect 17405 14835 17463 14841
rect 9769 14807 9827 14813
rect 9769 14804 9781 14807
rect 9732 14776 9781 14804
rect 9732 14764 9738 14776
rect 9769 14773 9781 14776
rect 9815 14773 9827 14807
rect 9769 14767 9827 14773
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14773 11391 14807
rect 11698 14804 11704 14816
rect 11659 14776 11704 14804
rect 11333 14767 11391 14773
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 12710 14764 12716 14816
rect 12768 14804 12774 14816
rect 12805 14807 12863 14813
rect 12805 14804 12817 14807
rect 12768 14776 12817 14804
rect 12768 14764 12774 14776
rect 12805 14773 12817 14776
rect 12851 14773 12863 14807
rect 15010 14804 15016 14816
rect 14971 14776 15016 14804
rect 12805 14767 12863 14773
rect 15010 14764 15016 14776
rect 15068 14764 15074 14816
rect 15381 14807 15439 14813
rect 15381 14773 15393 14807
rect 15427 14804 15439 14807
rect 15654 14804 15660 14816
rect 15427 14776 15660 14804
rect 15427 14773 15439 14776
rect 15381 14767 15439 14773
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 16209 14807 16267 14813
rect 16209 14773 16221 14807
rect 16255 14804 16267 14807
rect 17512 14804 17540 14912
rect 19889 14875 19947 14881
rect 19889 14872 19901 14875
rect 18432 14844 19901 14872
rect 18432 14813 18460 14844
rect 19889 14841 19901 14844
rect 19935 14841 19947 14875
rect 19996 14872 20024 14912
rect 20162 14900 20168 14952
rect 20220 14940 20226 14952
rect 20441 14943 20499 14949
rect 20441 14940 20453 14943
rect 20220 14912 20453 14940
rect 20220 14900 20226 14912
rect 20441 14909 20453 14912
rect 20487 14909 20499 14943
rect 20441 14903 20499 14909
rect 20898 14872 20904 14884
rect 19996 14844 20904 14872
rect 19889 14835 19947 14841
rect 20898 14832 20904 14844
rect 20956 14832 20962 14884
rect 16255 14776 17540 14804
rect 18417 14807 18475 14813
rect 16255 14773 16267 14776
rect 16209 14767 16267 14773
rect 18417 14773 18429 14807
rect 18463 14773 18475 14807
rect 18417 14767 18475 14773
rect 18785 14807 18843 14813
rect 18785 14773 18797 14807
rect 18831 14804 18843 14807
rect 19242 14804 19248 14816
rect 18831 14776 19248 14804
rect 18831 14773 18843 14776
rect 18785 14767 18843 14773
rect 19242 14764 19248 14776
rect 19300 14764 19306 14816
rect 19702 14764 19708 14816
rect 19760 14804 19766 14816
rect 19797 14807 19855 14813
rect 19797 14804 19809 14807
rect 19760 14776 19809 14804
rect 19760 14764 19766 14776
rect 19797 14773 19809 14776
rect 19843 14773 19855 14807
rect 19797 14767 19855 14773
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 8570 14600 8576 14612
rect 8531 14572 8576 14600
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 9030 14600 9036 14612
rect 8991 14572 9036 14600
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 9674 14600 9680 14612
rect 9635 14572 9680 14600
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 12434 14560 12440 14612
rect 12492 14600 12498 14612
rect 12492 14572 12537 14600
rect 12492 14560 12498 14572
rect 13078 14560 13084 14612
rect 13136 14600 13142 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13136 14572 14105 14600
rect 13136 14560 13142 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 15286 14600 15292 14612
rect 15247 14572 15292 14600
rect 14093 14563 14151 14569
rect 15286 14560 15292 14572
rect 15344 14560 15350 14612
rect 15654 14600 15660 14612
rect 15615 14572 15660 14600
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 15749 14603 15807 14609
rect 15749 14569 15761 14603
rect 15795 14600 15807 14603
rect 15838 14600 15844 14612
rect 15795 14572 15844 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 15838 14560 15844 14572
rect 15896 14560 15902 14612
rect 17678 14600 17684 14612
rect 17639 14572 17684 14600
rect 17678 14560 17684 14572
rect 17736 14560 17742 14612
rect 6914 14492 6920 14544
rect 6972 14532 6978 14544
rect 7184 14535 7242 14541
rect 7184 14532 7196 14535
rect 6972 14504 7196 14532
rect 6972 14492 6978 14504
rect 7184 14501 7196 14504
rect 7230 14532 7242 14535
rect 8202 14532 8208 14544
rect 7230 14504 8208 14532
rect 7230 14501 7242 14504
rect 7184 14495 7242 14501
rect 8202 14492 8208 14504
rect 8260 14492 8266 14544
rect 8941 14535 8999 14541
rect 8941 14501 8953 14535
rect 8987 14532 8999 14535
rect 11054 14532 11060 14544
rect 8987 14504 11060 14532
rect 8987 14501 8999 14504
rect 8941 14495 8999 14501
rect 11054 14492 11060 14504
rect 11112 14492 11118 14544
rect 11324 14535 11382 14541
rect 11324 14501 11336 14535
rect 11370 14532 11382 14535
rect 12342 14532 12348 14544
rect 11370 14504 12348 14532
rect 11370 14501 11382 14504
rect 11324 14495 11382 14501
rect 12342 14492 12348 14504
rect 12400 14492 12406 14544
rect 12452 14532 12480 14560
rect 12958 14535 13016 14541
rect 12958 14532 12970 14535
rect 12452 14504 12970 14532
rect 12958 14501 12970 14504
rect 13004 14532 13016 14535
rect 13630 14532 13636 14544
rect 13004 14504 13636 14532
rect 13004 14501 13016 14504
rect 12958 14495 13016 14501
rect 13630 14492 13636 14504
rect 13688 14492 13694 14544
rect 14550 14492 14556 14544
rect 14608 14532 14614 14544
rect 14645 14535 14703 14541
rect 14645 14532 14657 14535
rect 14608 14504 14657 14532
rect 14608 14492 14614 14504
rect 14645 14501 14657 14504
rect 14691 14501 14703 14535
rect 18868 14535 18926 14541
rect 14645 14495 14703 14501
rect 16316 14504 18644 14532
rect 10042 14464 10048 14476
rect 10003 14436 10048 14464
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 12066 14464 12072 14476
rect 11011 14436 12072 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 12066 14424 12072 14436
rect 12124 14424 12130 14476
rect 12713 14467 12771 14473
rect 12713 14433 12725 14467
rect 12759 14464 12771 14467
rect 13538 14464 13544 14476
rect 12759 14436 13544 14464
rect 12759 14433 12771 14436
rect 12713 14427 12771 14433
rect 13538 14424 13544 14436
rect 13596 14424 13602 14476
rect 14366 14464 14372 14476
rect 14327 14436 14372 14464
rect 14366 14424 14372 14436
rect 14424 14424 14430 14476
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14365 6975 14399
rect 6917 14359 6975 14365
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14365 9275 14399
rect 10134 14396 10140 14408
rect 10095 14368 10140 14396
rect 9217 14359 9275 14365
rect 6932 14260 6960 14359
rect 8294 14328 8300 14340
rect 8207 14300 8300 14328
rect 8294 14288 8300 14300
rect 8352 14328 8358 14340
rect 9232 14328 9260 14359
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 11057 14399 11115 14405
rect 11057 14396 11069 14399
rect 10229 14359 10287 14365
rect 10336 14368 11069 14396
rect 10244 14328 10272 14359
rect 8352 14300 10272 14328
rect 8352 14288 8358 14300
rect 9214 14260 9220 14272
rect 6932 14232 9220 14260
rect 9214 14220 9220 14232
rect 9272 14260 9278 14272
rect 10336 14260 10364 14368
rect 11057 14365 11069 14368
rect 11103 14365 11115 14399
rect 11057 14359 11115 14365
rect 15562 14356 15568 14408
rect 15620 14396 15626 14408
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15620 14368 15853 14396
rect 15620 14356 15626 14368
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 16206 14356 16212 14408
rect 16264 14396 16270 14408
rect 16316 14405 16344 14504
rect 16568 14467 16626 14473
rect 16568 14433 16580 14467
rect 16614 14464 16626 14467
rect 17586 14464 17592 14476
rect 16614 14436 17592 14464
rect 16614 14433 16626 14436
rect 16568 14427 16626 14433
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 18616 14473 18644 14504
rect 18868 14501 18880 14535
rect 18914 14532 18926 14535
rect 19794 14532 19800 14544
rect 18914 14504 19800 14532
rect 18914 14501 18926 14504
rect 18868 14495 18926 14501
rect 19794 14492 19800 14504
rect 19852 14492 19858 14544
rect 18601 14467 18659 14473
rect 18601 14433 18613 14467
rect 18647 14433 18659 14467
rect 20254 14464 20260 14476
rect 20215 14436 20260 14464
rect 18601 14427 18659 14433
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 16301 14399 16359 14405
rect 16301 14396 16313 14399
rect 16264 14368 16313 14396
rect 16264 14356 16270 14368
rect 16301 14365 16313 14368
rect 16347 14365 16359 14399
rect 17954 14396 17960 14408
rect 17915 14368 17960 14396
rect 16301 14359 16359 14365
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 20070 14356 20076 14408
rect 20128 14396 20134 14408
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20128 14368 20913 14396
rect 20128 14356 20134 14368
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 9272 14232 10364 14260
rect 9272 14220 9278 14232
rect 10502 14220 10508 14272
rect 10560 14260 10566 14272
rect 10781 14263 10839 14269
rect 10781 14260 10793 14263
rect 10560 14232 10793 14260
rect 10560 14220 10566 14232
rect 10781 14229 10793 14232
rect 10827 14229 10839 14263
rect 10781 14223 10839 14229
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 19978 14260 19984 14272
rect 13688 14232 19984 14260
rect 13688 14220 13694 14232
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 20438 14260 20444 14272
rect 20399 14232 20444 14260
rect 20438 14220 20444 14232
rect 20496 14220 20502 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 11698 14056 11704 14068
rect 11379 14028 11704 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 12710 14056 12716 14068
rect 12671 14028 12716 14056
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 13541 14059 13599 14065
rect 13541 14025 13553 14059
rect 13587 14056 13599 14059
rect 13725 14059 13783 14065
rect 13725 14056 13737 14059
rect 13587 14028 13737 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 13725 14025 13737 14028
rect 13771 14025 13783 14059
rect 13725 14019 13783 14025
rect 15933 14059 15991 14065
rect 15933 14025 15945 14059
rect 15979 14056 15991 14059
rect 16482 14056 16488 14068
rect 15979 14028 16488 14056
rect 15979 14025 15991 14028
rect 15933 14019 15991 14025
rect 16482 14016 16488 14028
rect 16540 14016 16546 14068
rect 16942 14016 16948 14068
rect 17000 14056 17006 14068
rect 17586 14056 17592 14068
rect 17000 14028 17448 14056
rect 17547 14028 17592 14056
rect 17000 14016 17006 14028
rect 15746 13988 15752 14000
rect 11808 13960 15752 13988
rect 11808 13932 11836 13960
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 17420 13988 17448 14028
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 19702 14056 19708 14068
rect 19663 14028 19708 14056
rect 19702 14016 19708 14028
rect 19760 14016 19766 14068
rect 20898 14056 20904 14068
rect 20859 14028 20904 14056
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 17420 13960 19187 13988
rect 9214 13920 9220 13932
rect 9175 13892 9220 13920
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 11790 13920 11796 13932
rect 11703 13892 11796 13920
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13920 12035 13923
rect 12342 13920 12348 13932
rect 12023 13892 12348 13920
rect 12023 13889 12035 13892
rect 11977 13883 12035 13889
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 13170 13920 13176 13932
rect 13131 13892 13176 13920
rect 13170 13880 13176 13892
rect 13228 13880 13234 13932
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13920 13415 13923
rect 13538 13920 13544 13932
rect 13403 13892 13544 13920
rect 13403 13889 13415 13892
rect 13357 13883 13415 13889
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 14182 13920 14188 13932
rect 14143 13892 14188 13920
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13920 14427 13923
rect 15010 13920 15016 13932
rect 14415 13892 15016 13920
rect 14415 13889 14427 13892
rect 14369 13883 14427 13889
rect 9484 13855 9542 13861
rect 9484 13821 9496 13855
rect 9530 13852 9542 13855
rect 13630 13852 13636 13864
rect 9530 13824 13636 13852
rect 9530 13821 9542 13824
rect 9484 13815 9542 13821
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 14384 13852 14412 13883
rect 15010 13880 15016 13892
rect 15068 13880 15074 13932
rect 15562 13920 15568 13932
rect 15523 13892 15568 13920
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 13780 13824 14412 13852
rect 15381 13855 15439 13861
rect 13780 13812 13786 13824
rect 15381 13821 15393 13855
rect 15427 13852 15439 13855
rect 15427 13824 15516 13852
rect 15427 13821 15439 13824
rect 15381 13815 15439 13821
rect 15488 13796 15516 13824
rect 15838 13812 15844 13864
rect 15896 13852 15902 13864
rect 16109 13855 16167 13861
rect 16109 13852 16121 13855
rect 15896 13824 16121 13852
rect 15896 13812 15902 13824
rect 16109 13821 16121 13824
rect 16155 13821 16167 13855
rect 16109 13815 16167 13821
rect 16209 13855 16267 13861
rect 16209 13821 16221 13855
rect 16255 13852 16267 13855
rect 16298 13852 16304 13864
rect 16255 13824 16304 13852
rect 16255 13821 16267 13824
rect 16209 13815 16267 13821
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 16476 13855 16534 13861
rect 16476 13821 16488 13855
rect 16522 13852 16534 13855
rect 16850 13852 16856 13864
rect 16522 13824 16856 13852
rect 16522 13821 16534 13824
rect 16476 13815 16534 13821
rect 16850 13812 16856 13824
rect 16908 13852 16914 13864
rect 18616 13852 18644 13883
rect 19058 13852 19064 13864
rect 16908 13824 19064 13852
rect 16908 13812 16914 13824
rect 19058 13812 19064 13824
rect 19116 13812 19122 13864
rect 19159 13852 19187 13960
rect 19794 13880 19800 13932
rect 19852 13920 19858 13932
rect 20257 13923 20315 13929
rect 20257 13920 20269 13923
rect 19852 13892 20269 13920
rect 19852 13880 19858 13892
rect 20257 13889 20269 13892
rect 20303 13889 20315 13923
rect 20257 13883 20315 13889
rect 20165 13855 20223 13861
rect 20165 13852 20177 13855
rect 19159 13824 20177 13852
rect 20165 13821 20177 13824
rect 20211 13821 20223 13855
rect 20714 13852 20720 13864
rect 20675 13824 20720 13852
rect 20165 13815 20223 13821
rect 20714 13812 20720 13824
rect 20772 13812 20778 13864
rect 8757 13787 8815 13793
rect 8757 13753 8769 13787
rect 8803 13784 8815 13787
rect 10042 13784 10048 13796
rect 8803 13756 10048 13784
rect 8803 13753 8815 13756
rect 8757 13747 8815 13753
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 13081 13787 13139 13793
rect 10428 13756 11744 13784
rect 9582 13676 9588 13728
rect 9640 13716 9646 13728
rect 10428 13716 10456 13756
rect 10594 13716 10600 13728
rect 9640 13688 10456 13716
rect 10555 13688 10600 13716
rect 9640 13676 9646 13688
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 11716 13725 11744 13756
rect 13081 13753 13093 13787
rect 13127 13784 13139 13787
rect 13541 13787 13599 13793
rect 13541 13784 13553 13787
rect 13127 13756 13553 13784
rect 13127 13753 13139 13756
rect 13081 13747 13139 13753
rect 13541 13753 13553 13756
rect 13587 13753 13599 13787
rect 13541 13747 13599 13753
rect 13648 13756 15424 13784
rect 11701 13719 11759 13725
rect 11701 13685 11713 13719
rect 11747 13716 11759 13719
rect 13648 13716 13676 13756
rect 14090 13716 14096 13728
rect 11747 13688 13676 13716
rect 14051 13688 14096 13716
rect 11747 13685 11759 13688
rect 11701 13679 11759 13685
rect 14090 13676 14096 13688
rect 14148 13676 14154 13728
rect 14550 13676 14556 13728
rect 14608 13716 14614 13728
rect 14921 13719 14979 13725
rect 14921 13716 14933 13719
rect 14608 13688 14933 13716
rect 14608 13676 14614 13688
rect 14921 13685 14933 13688
rect 14967 13685 14979 13719
rect 15286 13716 15292 13728
rect 15247 13688 15292 13716
rect 14921 13679 14979 13685
rect 15286 13676 15292 13688
rect 15344 13676 15350 13728
rect 15396 13716 15424 13756
rect 15470 13744 15476 13796
rect 15528 13744 15534 13796
rect 15654 13744 15660 13796
rect 15712 13784 15718 13796
rect 16666 13784 16672 13796
rect 15712 13756 16672 13784
rect 15712 13744 15718 13756
rect 16666 13744 16672 13756
rect 16724 13744 16730 13796
rect 18509 13787 18567 13793
rect 18509 13784 18521 13787
rect 16776 13756 18521 13784
rect 16776 13716 16804 13756
rect 18509 13753 18521 13756
rect 18555 13784 18567 13787
rect 18782 13784 18788 13796
rect 18555 13756 18788 13784
rect 18555 13753 18567 13756
rect 18509 13747 18567 13753
rect 18782 13744 18788 13756
rect 18840 13744 18846 13796
rect 20070 13784 20076 13796
rect 20031 13756 20076 13784
rect 20070 13744 20076 13756
rect 20128 13744 20134 13796
rect 18046 13716 18052 13728
rect 15396 13688 16804 13716
rect 18007 13688 18052 13716
rect 18046 13676 18052 13688
rect 18104 13676 18110 13728
rect 18414 13716 18420 13728
rect 18375 13688 18420 13716
rect 18414 13676 18420 13688
rect 18472 13676 18478 13728
rect 18690 13676 18696 13728
rect 18748 13716 18754 13728
rect 18966 13716 18972 13728
rect 18748 13688 18972 13716
rect 18748 13676 18754 13688
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 9769 13515 9827 13521
rect 9769 13481 9781 13515
rect 9815 13512 9827 13515
rect 10962 13512 10968 13524
rect 9815 13484 10968 13512
rect 9815 13481 9827 13484
rect 9769 13475 9827 13481
rect 10962 13472 10968 13484
rect 11020 13472 11026 13524
rect 11241 13515 11299 13521
rect 11241 13481 11253 13515
rect 11287 13512 11299 13515
rect 11606 13512 11612 13524
rect 11287 13484 11612 13512
rect 11287 13481 11299 13484
rect 11241 13475 11299 13481
rect 11606 13472 11612 13484
rect 11664 13512 11670 13524
rect 11974 13512 11980 13524
rect 11664 13484 11980 13512
rect 11664 13472 11670 13484
rect 11974 13472 11980 13484
rect 12032 13472 12038 13524
rect 13170 13512 13176 13524
rect 13131 13484 13176 13512
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 14550 13512 14556 13524
rect 14511 13484 14556 13512
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 16761 13515 16819 13521
rect 16761 13481 16773 13515
rect 16807 13512 16819 13515
rect 17034 13512 17040 13524
rect 16807 13484 17040 13512
rect 16807 13481 16819 13484
rect 16761 13475 16819 13481
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 17221 13515 17279 13521
rect 17221 13481 17233 13515
rect 17267 13512 17279 13515
rect 17773 13515 17831 13521
rect 17773 13512 17785 13515
rect 17267 13484 17785 13512
rect 17267 13481 17279 13484
rect 17221 13475 17279 13481
rect 17773 13481 17785 13484
rect 17819 13481 17831 13515
rect 17773 13475 17831 13481
rect 18046 13472 18052 13524
rect 18104 13512 18110 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 18104 13484 18153 13512
rect 18104 13472 18110 13484
rect 18141 13481 18153 13484
rect 18187 13481 18199 13515
rect 18141 13475 18199 13481
rect 18233 13515 18291 13521
rect 18233 13481 18245 13515
rect 18279 13512 18291 13515
rect 18785 13515 18843 13521
rect 18785 13512 18797 13515
rect 18279 13484 18797 13512
rect 18279 13481 18291 13484
rect 18233 13475 18291 13481
rect 18785 13481 18797 13484
rect 18831 13481 18843 13515
rect 18785 13475 18843 13481
rect 19797 13515 19855 13521
rect 19797 13481 19809 13515
rect 19843 13512 19855 13515
rect 20162 13512 20168 13524
rect 19843 13484 20168 13512
rect 19843 13481 19855 13484
rect 19797 13475 19855 13481
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 11054 13404 11060 13456
rect 11112 13444 11118 13456
rect 11149 13447 11207 13453
rect 11149 13444 11161 13447
rect 11112 13416 11161 13444
rect 11112 13404 11118 13416
rect 11149 13413 11161 13416
rect 11195 13444 11207 13447
rect 11790 13444 11796 13456
rect 11195 13416 11796 13444
rect 11195 13413 11207 13416
rect 11149 13407 11207 13413
rect 11790 13404 11796 13416
rect 11848 13404 11854 13456
rect 13541 13447 13599 13453
rect 13541 13413 13553 13447
rect 13587 13444 13599 13447
rect 13630 13444 13636 13456
rect 13587 13416 13636 13444
rect 13587 13413 13599 13416
rect 13541 13407 13599 13413
rect 13630 13404 13636 13416
rect 13688 13404 13694 13456
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 13998 13444 14004 13456
rect 13872 13416 14004 13444
rect 13872 13404 13878 13416
rect 13998 13404 14004 13416
rect 14056 13404 14062 13456
rect 14090 13404 14096 13456
rect 14148 13444 14154 13456
rect 15289 13447 15347 13453
rect 15289 13444 15301 13447
rect 14148 13416 15301 13444
rect 14148 13404 14154 13416
rect 15289 13413 15301 13416
rect 15335 13413 15347 13447
rect 15289 13407 15347 13413
rect 15746 13404 15752 13456
rect 15804 13444 15810 13456
rect 15804 13416 19012 13444
rect 15804 13404 15810 13416
rect 10134 13376 10140 13388
rect 10095 13348 10140 13376
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 12342 13376 12348 13388
rect 12303 13348 12348 13376
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 12526 13336 12532 13388
rect 12584 13376 12590 13388
rect 13170 13376 13176 13388
rect 12584 13348 13176 13376
rect 12584 13336 12590 13348
rect 13170 13336 13176 13348
rect 13228 13336 13234 13388
rect 13722 13336 13728 13388
rect 13780 13336 13786 13388
rect 14016 13376 14044 13404
rect 18984 13388 19012 13416
rect 16117 13379 16175 13385
rect 16117 13376 16129 13379
rect 14016 13348 16129 13376
rect 16117 13345 16129 13348
rect 16163 13345 16175 13379
rect 16117 13339 16175 13345
rect 16209 13379 16267 13385
rect 16209 13345 16221 13379
rect 16255 13376 16267 13379
rect 16390 13376 16396 13388
rect 16255 13348 16396 13376
rect 16255 13345 16267 13348
rect 16209 13339 16267 13345
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 16574 13336 16580 13388
rect 16632 13376 16638 13388
rect 17129 13379 17187 13385
rect 17129 13376 17141 13379
rect 16632 13348 17141 13376
rect 16632 13336 16638 13348
rect 17129 13345 17141 13348
rect 17175 13345 17187 13379
rect 17129 13339 17187 13345
rect 17586 13336 17592 13388
rect 17644 13376 17650 13388
rect 17644 13348 18368 13376
rect 17644 13336 17650 13348
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 10244 13240 10272 13271
rect 10318 13268 10324 13320
rect 10376 13308 10382 13320
rect 10376 13280 10421 13308
rect 10376 13268 10382 13280
rect 10594 13268 10600 13320
rect 10652 13308 10658 13320
rect 11333 13311 11391 13317
rect 10652 13280 11192 13308
rect 10652 13268 10658 13280
rect 11054 13240 11060 13252
rect 10244 13212 11060 13240
rect 11054 13200 11060 13212
rect 11112 13200 11118 13252
rect 11164 13240 11192 13280
rect 11333 13277 11345 13311
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 12437 13311 12495 13317
rect 12437 13277 12449 13311
rect 12483 13277 12495 13311
rect 12618 13308 12624 13320
rect 12579 13280 12624 13308
rect 12437 13271 12495 13277
rect 11348 13240 11376 13271
rect 11164 13212 11376 13240
rect 12452 13240 12480 13271
rect 12618 13268 12624 13280
rect 12676 13268 12682 13320
rect 13633 13311 13691 13317
rect 13633 13277 13645 13311
rect 13679 13277 13691 13311
rect 13740 13308 13768 13336
rect 13817 13311 13875 13317
rect 13817 13308 13829 13311
rect 13740 13280 13829 13308
rect 13633 13271 13691 13277
rect 13817 13277 13829 13280
rect 13863 13277 13875 13311
rect 13817 13271 13875 13277
rect 13538 13240 13544 13252
rect 12452 13212 13544 13240
rect 13538 13200 13544 13212
rect 13596 13200 13602 13252
rect 13648 13240 13676 13271
rect 13998 13268 14004 13320
rect 14056 13308 14062 13320
rect 14645 13311 14703 13317
rect 14645 13308 14657 13311
rect 14056 13280 14657 13308
rect 14056 13268 14062 13280
rect 14645 13277 14657 13280
rect 14691 13277 14703 13311
rect 14645 13271 14703 13277
rect 14734 13268 14740 13320
rect 14792 13308 14798 13320
rect 16301 13311 16359 13317
rect 14792 13280 14837 13308
rect 14792 13268 14798 13280
rect 16301 13277 16313 13311
rect 16347 13308 16359 13311
rect 16850 13308 16856 13320
rect 16347 13280 16856 13308
rect 16347 13277 16359 13280
rect 16301 13271 16359 13277
rect 16850 13268 16856 13280
rect 16908 13268 16914 13320
rect 17405 13311 17463 13317
rect 17405 13277 17417 13311
rect 17451 13308 17463 13311
rect 17678 13308 17684 13320
rect 17451 13280 17684 13308
rect 17451 13277 17463 13280
rect 17405 13271 17463 13277
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 18340 13317 18368 13348
rect 18966 13336 18972 13388
rect 19024 13376 19030 13388
rect 19153 13379 19211 13385
rect 19153 13376 19165 13379
rect 19024 13348 19165 13376
rect 19024 13336 19030 13348
rect 19153 13345 19165 13348
rect 19199 13345 19211 13379
rect 19153 13339 19211 13345
rect 19426 13336 19432 13388
rect 19484 13376 19490 13388
rect 20165 13379 20223 13385
rect 20165 13376 20177 13379
rect 19484 13348 20177 13376
rect 19484 13336 19490 13348
rect 20165 13345 20177 13348
rect 20211 13345 20223 13379
rect 20165 13339 20223 13345
rect 18325 13311 18383 13317
rect 18325 13277 18337 13311
rect 18371 13277 18383 13311
rect 19242 13308 19248 13320
rect 19203 13280 19248 13308
rect 18325 13271 18383 13277
rect 19242 13268 19248 13280
rect 19300 13268 19306 13320
rect 19337 13311 19395 13317
rect 19337 13277 19349 13311
rect 19383 13277 19395 13311
rect 20254 13308 20260 13320
rect 20215 13280 20260 13308
rect 19337 13271 19395 13277
rect 16666 13240 16672 13252
rect 13648 13212 16672 13240
rect 16666 13200 16672 13212
rect 16724 13240 16730 13252
rect 17218 13240 17224 13252
rect 16724 13212 17224 13240
rect 16724 13200 16730 13212
rect 17218 13200 17224 13212
rect 17276 13240 17282 13252
rect 18414 13240 18420 13252
rect 17276 13212 18420 13240
rect 17276 13200 17282 13212
rect 18414 13200 18420 13212
rect 18472 13200 18478 13252
rect 19058 13200 19064 13252
rect 19116 13240 19122 13252
rect 19352 13240 19380 13271
rect 20254 13268 20260 13280
rect 20312 13268 20318 13320
rect 20349 13311 20407 13317
rect 20349 13277 20361 13311
rect 20395 13277 20407 13311
rect 20349 13271 20407 13277
rect 19116 13212 19380 13240
rect 19116 13200 19122 13212
rect 19978 13200 19984 13252
rect 20036 13240 20042 13252
rect 20364 13240 20392 13271
rect 20036 13212 20392 13240
rect 20036 13200 20042 13212
rect 10778 13172 10784 13184
rect 10739 13144 10784 13172
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 11977 13175 12035 13181
rect 11977 13141 11989 13175
rect 12023 13172 12035 13175
rect 12434 13172 12440 13184
rect 12023 13144 12440 13172
rect 12023 13141 12035 13144
rect 11977 13135 12035 13141
rect 12434 13132 12440 13144
rect 12492 13132 12498 13184
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 14185 13175 14243 13181
rect 14185 13172 14197 13175
rect 13872 13144 14197 13172
rect 13872 13132 13878 13144
rect 14185 13141 14197 13144
rect 14231 13141 14243 13175
rect 15746 13172 15752 13184
rect 15707 13144 15752 13172
rect 14185 13135 14243 13141
rect 15746 13132 15752 13144
rect 15804 13132 15810 13184
rect 16298 13132 16304 13184
rect 16356 13172 16362 13184
rect 17770 13172 17776 13184
rect 16356 13144 17776 13172
rect 16356 13132 16362 13144
rect 17770 13132 17776 13144
rect 17828 13132 17834 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 9125 12971 9183 12977
rect 9125 12937 9137 12971
rect 9171 12968 9183 12971
rect 9214 12968 9220 12980
rect 9171 12940 9220 12968
rect 9171 12937 9183 12940
rect 9125 12931 9183 12937
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12937 10839 12971
rect 11054 12968 11060 12980
rect 11015 12940 11060 12968
rect 10781 12931 10839 12937
rect 8478 12792 8484 12844
rect 8536 12832 8542 12844
rect 9232 12832 9260 12928
rect 10796 12900 10824 12931
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 13357 12971 13415 12977
rect 13357 12937 13369 12971
rect 13403 12968 13415 12971
rect 14274 12968 14280 12980
rect 13403 12940 14280 12968
rect 13403 12937 13415 12940
rect 13357 12931 13415 12937
rect 14274 12928 14280 12940
rect 14332 12928 14338 12980
rect 15838 12968 15844 12980
rect 14384 12940 15844 12968
rect 10870 12900 10876 12912
rect 10783 12872 10876 12900
rect 10870 12860 10876 12872
rect 10928 12900 10934 12912
rect 12066 12900 12072 12912
rect 10928 12872 11652 12900
rect 11979 12872 12072 12900
rect 10928 12860 10934 12872
rect 9401 12835 9459 12841
rect 9401 12832 9413 12835
rect 8536 12804 9413 12832
rect 8536 12792 8542 12804
rect 9401 12801 9413 12804
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 10778 12792 10784 12844
rect 10836 12832 10842 12844
rect 11624 12841 11652 12872
rect 12066 12860 12072 12872
rect 12124 12900 12130 12912
rect 14384 12900 14412 12940
rect 15838 12928 15844 12940
rect 15896 12928 15902 12980
rect 16574 12968 16580 12980
rect 16535 12940 16580 12968
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 18325 12971 18383 12977
rect 18325 12937 18337 12971
rect 18371 12968 18383 12971
rect 18598 12968 18604 12980
rect 18371 12940 18604 12968
rect 18371 12937 18383 12940
rect 18325 12931 18383 12937
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 19058 12928 19064 12980
rect 19116 12968 19122 12980
rect 20073 12971 20131 12977
rect 20073 12968 20085 12971
rect 19116 12940 20085 12968
rect 19116 12928 19122 12940
rect 20073 12937 20085 12940
rect 20119 12937 20131 12971
rect 20073 12931 20131 12937
rect 12124 12872 14412 12900
rect 12124 12860 12130 12872
rect 16206 12860 16212 12912
rect 16264 12900 16270 12912
rect 16264 12872 18736 12900
rect 16264 12860 16270 12872
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 10836 12804 11529 12832
rect 10836 12792 10842 12804
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 11609 12835 11667 12841
rect 11609 12801 11621 12835
rect 11655 12801 11667 12835
rect 11609 12795 11667 12801
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12832 12771 12835
rect 12986 12832 12992 12844
rect 12759 12804 12992 12832
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13814 12832 13820 12844
rect 13775 12804 13820 12832
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12832 14059 12835
rect 14047 12804 14504 12832
rect 14047 12801 14059 12804
rect 14001 12795 14059 12801
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 9668 12767 9726 12773
rect 9668 12733 9680 12767
rect 9714 12764 9726 12767
rect 10594 12764 10600 12776
rect 9714 12736 10600 12764
rect 9714 12733 9726 12736
rect 9668 12727 9726 12733
rect 9324 12696 9352 12727
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 11882 12724 11888 12776
rect 11940 12764 11946 12776
rect 12158 12764 12164 12776
rect 11940 12736 12164 12764
rect 11940 12724 11946 12736
rect 12158 12724 12164 12736
rect 12216 12724 12222 12776
rect 12253 12767 12311 12773
rect 12253 12733 12265 12767
rect 12299 12733 12311 12767
rect 12253 12727 12311 12733
rect 10502 12696 10508 12708
rect 9324 12668 10508 12696
rect 10502 12656 10508 12668
rect 10560 12656 10566 12708
rect 11422 12696 11428 12708
rect 11383 12668 11428 12696
rect 11422 12656 11428 12668
rect 11480 12656 11486 12708
rect 12268 12696 12296 12727
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 14182 12764 14188 12776
rect 12492 12736 12537 12764
rect 12636 12736 14188 12764
rect 12492 12724 12498 12736
rect 12636 12696 12664 12736
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 14369 12767 14427 12773
rect 14369 12733 14381 12767
rect 14415 12733 14427 12767
rect 14369 12727 14427 12733
rect 12268 12668 12664 12696
rect 13354 12656 13360 12708
rect 13412 12696 13418 12708
rect 14384 12696 14412 12727
rect 13412 12668 14412 12696
rect 13412 12656 13418 12668
rect 13725 12631 13783 12637
rect 13725 12597 13737 12631
rect 13771 12628 13783 12631
rect 14366 12628 14372 12640
rect 13771 12600 14372 12628
rect 13771 12597 13783 12600
rect 13725 12591 13783 12597
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 14476 12628 14504 12804
rect 15746 12792 15752 12844
rect 15804 12832 15810 12844
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 15804 12804 17049 12832
rect 15804 12792 15810 12804
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12832 17279 12835
rect 17586 12832 17592 12844
rect 17267 12804 17592 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 17586 12792 17592 12804
rect 17644 12792 17650 12844
rect 18598 12792 18604 12844
rect 18656 12832 18662 12844
rect 18708 12841 18736 12872
rect 18693 12835 18751 12841
rect 18693 12832 18705 12835
rect 18656 12804 18705 12832
rect 18656 12792 18662 12804
rect 18693 12801 18705 12804
rect 18739 12801 18751 12835
rect 18693 12795 18751 12801
rect 19794 12792 19800 12844
rect 19852 12832 19858 12844
rect 20901 12835 20959 12841
rect 20901 12832 20913 12835
rect 19852 12804 20913 12832
rect 19852 12792 19858 12804
rect 20901 12801 20913 12804
rect 20947 12801 20959 12835
rect 20901 12795 20959 12801
rect 16393 12767 16451 12773
rect 16393 12733 16405 12767
rect 16439 12764 16451 12767
rect 16482 12764 16488 12776
rect 16439 12736 16488 12764
rect 16439 12733 16451 12736
rect 16393 12727 16451 12733
rect 16482 12724 16488 12736
rect 16540 12724 16546 12776
rect 16945 12767 17003 12773
rect 16945 12733 16957 12767
rect 16991 12764 17003 12767
rect 17954 12764 17960 12776
rect 16991 12736 17960 12764
rect 16991 12733 17003 12736
rect 16945 12727 17003 12733
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 18138 12764 18144 12776
rect 18099 12736 18144 12764
rect 18138 12724 18144 12736
rect 18196 12724 18202 12776
rect 18960 12767 19018 12773
rect 18960 12733 18972 12767
rect 19006 12764 19018 12767
rect 19978 12764 19984 12776
rect 19006 12736 19984 12764
rect 19006 12733 19018 12736
rect 18960 12727 19018 12733
rect 19978 12724 19984 12736
rect 20036 12724 20042 12776
rect 14550 12656 14556 12708
rect 14608 12705 14614 12708
rect 14608 12699 14672 12705
rect 14608 12665 14626 12699
rect 14660 12696 14672 12699
rect 14734 12696 14740 12708
rect 14660 12668 14740 12696
rect 14660 12665 14672 12668
rect 14608 12659 14672 12665
rect 14608 12656 14614 12659
rect 14734 12656 14740 12668
rect 14792 12656 14798 12708
rect 17586 12656 17592 12708
rect 17644 12696 17650 12708
rect 17644 12668 20392 12696
rect 17644 12656 17650 12668
rect 15746 12628 15752 12640
rect 14476 12600 15752 12628
rect 15746 12588 15752 12600
rect 15804 12588 15810 12640
rect 15838 12588 15844 12640
rect 15896 12628 15902 12640
rect 16206 12628 16212 12640
rect 15896 12600 16212 12628
rect 15896 12588 15902 12600
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 20364 12637 20392 12668
rect 20622 12656 20628 12708
rect 20680 12696 20686 12708
rect 20809 12699 20867 12705
rect 20809 12696 20821 12699
rect 20680 12668 20821 12696
rect 20680 12656 20686 12668
rect 20809 12665 20821 12668
rect 20855 12665 20867 12699
rect 20809 12659 20867 12665
rect 20349 12631 20407 12637
rect 20349 12597 20361 12631
rect 20395 12597 20407 12631
rect 20349 12591 20407 12597
rect 20530 12588 20536 12640
rect 20588 12628 20594 12640
rect 20717 12631 20775 12637
rect 20717 12628 20729 12631
rect 20588 12600 20729 12628
rect 20588 12588 20594 12600
rect 20717 12597 20729 12600
rect 20763 12597 20775 12631
rect 20717 12591 20775 12597
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 11057 12427 11115 12433
rect 11057 12393 11069 12427
rect 11103 12393 11115 12427
rect 11057 12387 11115 12393
rect 7736 12359 7794 12365
rect 7736 12325 7748 12359
rect 7782 12356 7794 12359
rect 10318 12356 10324 12368
rect 7782 12328 10324 12356
rect 7782 12325 7794 12328
rect 7736 12319 7794 12325
rect 10318 12316 10324 12328
rect 10376 12356 10382 12368
rect 11072 12356 11100 12387
rect 12618 12384 12624 12436
rect 12676 12424 12682 12436
rect 12805 12427 12863 12433
rect 12805 12424 12817 12427
rect 12676 12396 12817 12424
rect 12676 12384 12682 12396
rect 12805 12393 12817 12396
rect 12851 12393 12863 12427
rect 12805 12387 12863 12393
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17862 12424 17868 12436
rect 17000 12396 17868 12424
rect 17000 12384 17006 12396
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 19978 12424 19984 12436
rect 19939 12396 19984 12424
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 20438 12424 20444 12436
rect 20399 12396 20444 12424
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 10376 12328 11100 12356
rect 13716 12359 13774 12365
rect 10376 12316 10382 12328
rect 13716 12325 13728 12359
rect 13762 12356 13774 12359
rect 13814 12356 13820 12368
rect 13762 12328 13820 12356
rect 13762 12325 13774 12328
rect 13716 12319 13774 12325
rect 13814 12316 13820 12328
rect 13872 12316 13878 12368
rect 15746 12316 15752 12368
rect 15804 12356 15810 12368
rect 15994 12359 16052 12365
rect 15994 12356 16006 12359
rect 15804 12328 16006 12356
rect 15804 12316 15810 12328
rect 15994 12325 16006 12328
rect 16040 12325 16052 12359
rect 15994 12319 16052 12325
rect 17773 12359 17831 12365
rect 17773 12325 17785 12359
rect 17819 12356 17831 12359
rect 17954 12356 17960 12368
rect 17819 12328 17960 12356
rect 17819 12325 17831 12328
rect 17773 12319 17831 12325
rect 17954 12316 17960 12328
rect 18012 12316 18018 12368
rect 18414 12316 18420 12368
rect 18472 12356 18478 12368
rect 18472 12328 20300 12356
rect 18472 12316 18478 12328
rect 8478 12288 8484 12300
rect 7484 12260 8484 12288
rect 7484 12232 7512 12260
rect 8478 12248 8484 12260
rect 8536 12288 8542 12300
rect 9677 12291 9735 12297
rect 9677 12288 9689 12291
rect 8536 12260 9689 12288
rect 8536 12248 8542 12260
rect 7466 12220 7472 12232
rect 7427 12192 7472 12220
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12220 9183 12223
rect 9490 12220 9496 12232
rect 9171 12192 9496 12220
rect 9171 12189 9183 12192
rect 9125 12183 9183 12189
rect 9490 12180 9496 12192
rect 9548 12180 9554 12232
rect 9398 12112 9404 12164
rect 9456 12152 9462 12164
rect 9600 12152 9628 12260
rect 9677 12257 9689 12260
rect 9723 12257 9735 12291
rect 9677 12251 9735 12257
rect 9944 12291 10002 12297
rect 9944 12257 9956 12291
rect 9990 12288 10002 12291
rect 10870 12288 10876 12300
rect 9990 12260 10876 12288
rect 9990 12257 10002 12260
rect 9944 12251 10002 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 11692 12291 11750 12297
rect 11692 12257 11704 12291
rect 11738 12288 11750 12291
rect 12250 12288 12256 12300
rect 11738 12260 12256 12288
rect 11738 12257 11750 12260
rect 11692 12251 11750 12257
rect 12250 12248 12256 12260
rect 12308 12248 12314 12300
rect 12526 12248 12532 12300
rect 12584 12288 12590 12300
rect 18138 12288 18144 12300
rect 12584 12260 18144 12288
rect 12584 12248 12590 12260
rect 18138 12248 18144 12260
rect 18196 12248 18202 12300
rect 18868 12291 18926 12297
rect 18868 12257 18880 12291
rect 18914 12288 18926 12291
rect 19242 12288 19248 12300
rect 18914 12260 19248 12288
rect 18914 12257 18926 12260
rect 18868 12251 18926 12257
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 20272 12297 20300 12328
rect 20257 12291 20315 12297
rect 20257 12257 20269 12291
rect 20303 12257 20315 12291
rect 20257 12251 20315 12257
rect 11425 12223 11483 12229
rect 11425 12220 11437 12223
rect 9456 12124 9628 12152
rect 9456 12112 9462 12124
rect 8849 12087 8907 12093
rect 8849 12053 8861 12087
rect 8895 12084 8907 12087
rect 9030 12084 9036 12096
rect 8895 12056 9036 12084
rect 8895 12053 8907 12056
rect 8849 12047 8907 12053
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 9600 12084 9628 12124
rect 10704 12192 11437 12220
rect 10704 12084 10732 12192
rect 11425 12189 11437 12192
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 9600 12056 10732 12084
rect 11440 12084 11468 12183
rect 13354 12180 13360 12232
rect 13412 12220 13418 12232
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 13412 12192 13461 12220
rect 13412 12180 13418 12192
rect 13449 12189 13461 12192
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 11790 12084 11796 12096
rect 11440 12056 11796 12084
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 13464 12084 13492 12183
rect 15102 12180 15108 12232
rect 15160 12220 15166 12232
rect 15289 12223 15347 12229
rect 15289 12220 15301 12223
rect 15160 12192 15301 12220
rect 15160 12180 15166 12192
rect 15289 12189 15301 12192
rect 15335 12189 15347 12223
rect 15746 12220 15752 12232
rect 15659 12192 15752 12220
rect 15289 12183 15347 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12189 18015 12223
rect 18598 12220 18604 12232
rect 18559 12192 18604 12220
rect 17957 12183 18015 12189
rect 15764 12152 15792 12180
rect 14476 12124 15792 12152
rect 14476 12084 14504 12124
rect 13464 12056 14504 12084
rect 14550 12044 14556 12096
rect 14608 12084 14614 12096
rect 14829 12087 14887 12093
rect 14829 12084 14841 12087
rect 14608 12056 14841 12084
rect 14608 12044 14614 12056
rect 14829 12053 14841 12056
rect 14875 12053 14887 12087
rect 17126 12084 17132 12096
rect 17087 12056 17132 12084
rect 14829 12047 14887 12053
rect 17126 12044 17132 12056
rect 17184 12044 17190 12096
rect 17218 12044 17224 12096
rect 17276 12084 17282 12096
rect 17405 12087 17463 12093
rect 17405 12084 17417 12087
rect 17276 12056 17417 12084
rect 17276 12044 17282 12056
rect 17405 12053 17417 12056
rect 17451 12053 17463 12087
rect 17405 12047 17463 12053
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 17972 12084 18000 12183
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 19610 12180 19616 12232
rect 19668 12220 19674 12232
rect 20901 12223 20959 12229
rect 20901 12220 20913 12223
rect 19668 12192 20913 12220
rect 19668 12180 19674 12192
rect 20901 12189 20913 12192
rect 20947 12189 20959 12223
rect 20901 12183 20959 12189
rect 17920 12056 18000 12084
rect 17920 12044 17926 12056
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 10229 11883 10287 11889
rect 10229 11880 10241 11883
rect 10192 11852 10241 11880
rect 10192 11840 10198 11852
rect 10229 11849 10241 11852
rect 10275 11849 10287 11883
rect 10229 11843 10287 11849
rect 11333 11883 11391 11889
rect 11333 11849 11345 11883
rect 11379 11880 11391 11883
rect 12342 11880 12348 11892
rect 11379 11852 12348 11880
rect 11379 11849 11391 11852
rect 11333 11843 11391 11849
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 13909 11883 13967 11889
rect 13909 11880 13921 11883
rect 13596 11852 13921 11880
rect 13596 11840 13602 11852
rect 13909 11849 13921 11852
rect 13955 11849 13967 11883
rect 13909 11843 13967 11849
rect 15838 11840 15844 11892
rect 15896 11880 15902 11892
rect 18693 11883 18751 11889
rect 15896 11852 18276 11880
rect 15896 11840 15902 11852
rect 18248 11824 18276 11852
rect 18693 11849 18705 11883
rect 18739 11880 18751 11883
rect 19426 11880 19432 11892
rect 18739 11852 19432 11880
rect 18739 11849 18751 11852
rect 18693 11843 18751 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 8297 11815 8355 11821
rect 8297 11781 8309 11815
rect 8343 11812 8355 11815
rect 8343 11784 9352 11812
rect 8343 11781 8355 11784
rect 8297 11775 8355 11781
rect 8846 11744 8852 11756
rect 8807 11716 8852 11744
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 9324 11685 9352 11784
rect 14090 11772 14096 11824
rect 14148 11812 14154 11824
rect 14148 11784 18184 11812
rect 14148 11772 14154 11784
rect 10870 11744 10876 11756
rect 10831 11716 10876 11744
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 12250 11744 12256 11756
rect 12023 11716 12256 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 12250 11704 12256 11716
rect 12308 11744 12314 11756
rect 14553 11747 14611 11753
rect 12308 11716 12572 11744
rect 12308 11704 12314 11716
rect 9309 11679 9367 11685
rect 9309 11645 9321 11679
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9490 11636 9496 11688
rect 9548 11676 9554 11688
rect 10597 11679 10655 11685
rect 10597 11676 10609 11679
rect 9548 11648 10609 11676
rect 9548 11636 9554 11648
rect 10597 11645 10609 11648
rect 10643 11645 10655 11679
rect 10597 11639 10655 11645
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 11848 11648 12449 11676
rect 11848 11636 11854 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12544 11676 12572 11716
rect 14553 11713 14565 11747
rect 14599 11713 14611 11747
rect 14553 11707 14611 11713
rect 12544 11648 14495 11676
rect 12437 11639 12495 11645
rect 9585 11611 9643 11617
rect 9585 11577 9597 11611
rect 9631 11608 9643 11611
rect 12526 11608 12532 11620
rect 9631 11580 12532 11608
rect 9631 11577 9643 11580
rect 9585 11571 9643 11577
rect 12526 11568 12532 11580
rect 12584 11568 12590 11620
rect 12618 11568 12624 11620
rect 12676 11617 12682 11620
rect 12676 11611 12740 11617
rect 12676 11577 12694 11611
rect 12728 11577 12740 11611
rect 12676 11571 12740 11577
rect 12676 11568 12682 11571
rect 13354 11568 13360 11620
rect 13412 11608 13418 11620
rect 14369 11611 14427 11617
rect 14369 11608 14381 11611
rect 13412 11580 14381 11608
rect 13412 11568 13418 11580
rect 14369 11577 14381 11580
rect 14415 11577 14427 11611
rect 14467 11608 14495 11648
rect 14568 11608 14596 11707
rect 15562 11704 15568 11756
rect 15620 11744 15626 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15620 11716 15945 11744
rect 15620 11704 15626 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 17497 11747 17555 11753
rect 17497 11713 17509 11747
rect 17543 11744 17555 11747
rect 17678 11744 17684 11756
rect 17543 11716 17684 11744
rect 17543 11713 17555 11716
rect 17497 11707 17555 11713
rect 17678 11704 17684 11716
rect 17736 11704 17742 11756
rect 17218 11676 17224 11688
rect 17179 11648 17224 11676
rect 17218 11636 17224 11648
rect 17276 11636 17282 11688
rect 18156 11685 18184 11784
rect 18230 11772 18236 11824
rect 18288 11772 18294 11824
rect 18325 11815 18383 11821
rect 18325 11781 18337 11815
rect 18371 11781 18383 11815
rect 18325 11775 18383 11781
rect 18340 11744 18368 11775
rect 18598 11772 18604 11824
rect 18656 11812 18662 11824
rect 18656 11784 19748 11812
rect 18656 11772 18662 11784
rect 18690 11744 18696 11756
rect 18340 11716 18696 11744
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 19242 11744 19248 11756
rect 19203 11716 19248 11744
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 19720 11753 19748 11784
rect 19705 11747 19763 11753
rect 19705 11713 19717 11747
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 18141 11679 18199 11685
rect 18141 11645 18153 11679
rect 18187 11645 18199 11679
rect 18141 11639 18199 11645
rect 19061 11679 19119 11685
rect 19061 11645 19073 11679
rect 19107 11676 19119 11679
rect 19610 11676 19616 11688
rect 19107 11648 19616 11676
rect 19107 11645 19119 11648
rect 19061 11639 19119 11645
rect 19610 11636 19616 11648
rect 19668 11636 19674 11688
rect 14467 11580 14596 11608
rect 14369 11571 14427 11577
rect 15286 11568 15292 11620
rect 15344 11608 15350 11620
rect 15470 11608 15476 11620
rect 15344 11580 15476 11608
rect 15344 11568 15350 11580
rect 15470 11568 15476 11580
rect 15528 11608 15534 11620
rect 18506 11608 18512 11620
rect 15528 11580 18512 11608
rect 15528 11568 15534 11580
rect 18506 11568 18512 11580
rect 18564 11568 18570 11620
rect 18690 11568 18696 11620
rect 18748 11608 18754 11620
rect 18874 11608 18880 11620
rect 18748 11580 18880 11608
rect 18748 11568 18754 11580
rect 18874 11568 18880 11580
rect 18932 11568 18938 11620
rect 19978 11617 19984 11620
rect 19972 11608 19984 11617
rect 19939 11580 19984 11608
rect 19972 11571 19984 11580
rect 19978 11568 19984 11571
rect 20036 11568 20042 11620
rect 8662 11540 8668 11552
rect 8623 11512 8668 11540
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 10689 11543 10747 11549
rect 8812 11512 8857 11540
rect 8812 11500 8818 11512
rect 10689 11509 10701 11543
rect 10735 11540 10747 11543
rect 11422 11540 11428 11552
rect 10735 11512 11428 11540
rect 10735 11509 10747 11512
rect 10689 11503 10747 11509
rect 11422 11500 11428 11512
rect 11480 11500 11486 11552
rect 11698 11540 11704 11552
rect 11659 11512 11704 11540
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 11793 11543 11851 11549
rect 11793 11509 11805 11543
rect 11839 11540 11851 11543
rect 12434 11540 12440 11552
rect 11839 11512 12440 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 13814 11540 13820 11552
rect 13775 11512 13820 11540
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 14274 11540 14280 11552
rect 14235 11512 14280 11540
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 15010 11500 15016 11552
rect 15068 11540 15074 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 15068 11512 15393 11540
rect 15068 11500 15074 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 15746 11540 15752 11552
rect 15707 11512 15752 11540
rect 15381 11503 15439 11509
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 15841 11543 15899 11549
rect 15841 11509 15853 11543
rect 15887 11540 15899 11543
rect 16206 11540 16212 11552
rect 15887 11512 16212 11540
rect 15887 11509 15899 11512
rect 15841 11503 15899 11509
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 16850 11500 16856 11552
rect 16908 11540 16914 11552
rect 17310 11540 17316 11552
rect 16908 11512 16953 11540
rect 17271 11512 17316 11540
rect 16908 11500 16914 11512
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 18598 11500 18604 11552
rect 18656 11540 18662 11552
rect 19153 11543 19211 11549
rect 19153 11540 19165 11543
rect 18656 11512 19165 11540
rect 18656 11500 18662 11512
rect 19153 11509 19165 11512
rect 19199 11509 19211 11543
rect 19153 11503 19211 11509
rect 19242 11500 19248 11552
rect 19300 11540 19306 11552
rect 21085 11543 21143 11549
rect 21085 11540 21097 11543
rect 19300 11512 21097 11540
rect 19300 11500 19306 11512
rect 21085 11509 21097 11512
rect 21131 11509 21143 11543
rect 21085 11503 21143 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 9033 11339 9091 11345
rect 9033 11336 9045 11339
rect 8720 11308 9045 11336
rect 8720 11296 8726 11308
rect 9033 11305 9045 11308
rect 9079 11305 9091 11339
rect 9033 11299 9091 11305
rect 9769 11339 9827 11345
rect 9769 11305 9781 11339
rect 9815 11336 9827 11339
rect 9815 11308 11376 11336
rect 9815 11305 9827 11308
rect 9769 11299 9827 11305
rect 10134 11268 10140 11280
rect 10095 11240 10140 11268
rect 10134 11228 10140 11240
rect 10192 11228 10198 11280
rect 10226 11228 10232 11280
rect 10284 11268 10290 11280
rect 10594 11268 10600 11280
rect 10284 11240 10600 11268
rect 10284 11228 10290 11240
rect 10594 11228 10600 11240
rect 10652 11228 10658 11280
rect 11348 11268 11376 11308
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 12437 11339 12495 11345
rect 12437 11336 12449 11339
rect 11756 11308 12449 11336
rect 11756 11296 11762 11308
rect 12437 11305 12449 11308
rect 12483 11305 12495 11339
rect 13998 11336 14004 11348
rect 12437 11299 12495 11305
rect 13004 11308 14004 11336
rect 13004 11268 13032 11308
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 14182 11296 14188 11348
rect 14240 11336 14246 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 14240 11308 14381 11336
rect 14240 11296 14246 11308
rect 14369 11305 14381 11308
rect 14415 11305 14427 11339
rect 14369 11299 14427 11305
rect 15654 11296 15660 11348
rect 15712 11336 15718 11348
rect 15933 11339 15991 11345
rect 15933 11336 15945 11339
rect 15712 11308 15945 11336
rect 15712 11296 15718 11308
rect 15933 11305 15945 11308
rect 15979 11305 15991 11339
rect 15933 11299 15991 11305
rect 16574 11296 16580 11348
rect 16632 11336 16638 11348
rect 17862 11336 17868 11348
rect 16632 11308 17868 11336
rect 16632 11296 16638 11308
rect 17862 11296 17868 11308
rect 17920 11336 17926 11348
rect 17957 11339 18015 11345
rect 17957 11336 17969 11339
rect 17920 11308 17969 11336
rect 17920 11296 17926 11308
rect 17957 11305 17969 11308
rect 18003 11305 18015 11339
rect 17957 11299 18015 11305
rect 19797 11339 19855 11345
rect 19797 11305 19809 11339
rect 19843 11336 19855 11339
rect 20254 11336 20260 11348
rect 19843 11308 20260 11336
rect 19843 11305 19855 11308
rect 19797 11299 19855 11305
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 10888 11240 11284 11268
rect 11348 11240 13032 11268
rect 13081 11271 13139 11277
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11200 7435 11203
rect 7466 11200 7472 11212
rect 7423 11172 7472 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 7466 11160 7472 11172
rect 7524 11160 7530 11212
rect 7644 11203 7702 11209
rect 7644 11169 7656 11203
rect 7690 11200 7702 11203
rect 9030 11200 9036 11212
rect 7690 11172 9036 11200
rect 7690 11169 7702 11172
rect 7644 11163 7702 11169
rect 9030 11160 9036 11172
rect 9088 11160 9094 11212
rect 9398 11160 9404 11212
rect 9456 11200 9462 11212
rect 10781 11203 10839 11209
rect 10781 11200 10793 11203
rect 9456 11172 10793 11200
rect 9456 11160 9462 11172
rect 10781 11169 10793 11172
rect 10827 11169 10839 11203
rect 10781 11163 10839 11169
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11132 10471 11135
rect 10888 11132 10916 11240
rect 11054 11209 11060 11212
rect 11048 11163 11060 11209
rect 11112 11200 11118 11212
rect 11256 11200 11284 11240
rect 13081 11237 13093 11271
rect 13127 11268 13139 11271
rect 13262 11268 13268 11280
rect 13127 11240 13268 11268
rect 13127 11237 13139 11240
rect 13081 11231 13139 11237
rect 13262 11228 13268 11240
rect 13320 11228 13326 11280
rect 16025 11271 16083 11277
rect 16025 11237 16037 11271
rect 16071 11268 16083 11271
rect 18598 11268 18604 11280
rect 16071 11240 18604 11268
rect 16071 11237 16083 11240
rect 16025 11231 16083 11237
rect 18598 11228 18604 11240
rect 18656 11228 18662 11280
rect 19153 11271 19211 11277
rect 19153 11237 19165 11271
rect 19199 11268 19211 11271
rect 19242 11268 19248 11280
rect 19199 11240 19248 11268
rect 19199 11237 19211 11240
rect 19153 11231 19211 11237
rect 19242 11228 19248 11240
rect 19300 11228 19306 11280
rect 19334 11228 19340 11280
rect 19392 11268 19398 11280
rect 19392 11240 20300 11268
rect 19392 11228 19398 11240
rect 13814 11200 13820 11212
rect 11112 11172 11148 11200
rect 11256 11172 13820 11200
rect 11054 11160 11060 11163
rect 11112 11160 11118 11172
rect 13814 11160 13820 11172
rect 13872 11200 13878 11212
rect 15562 11200 15568 11212
rect 13872 11172 15568 11200
rect 13872 11160 13878 11172
rect 15562 11160 15568 11172
rect 15620 11160 15626 11212
rect 16844 11203 16902 11209
rect 16844 11200 16856 11203
rect 16500 11172 16856 11200
rect 10459 11104 10916 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 13998 11132 14004 11144
rect 13780 11104 14004 11132
rect 13780 11092 13786 11104
rect 13998 11092 14004 11104
rect 14056 11092 14062 11144
rect 16209 11135 16267 11141
rect 16209 11101 16221 11135
rect 16255 11132 16267 11135
rect 16500 11132 16528 11172
rect 16844 11169 16856 11172
rect 16890 11200 16902 11203
rect 17218 11200 17224 11212
rect 16890 11172 17224 11200
rect 16890 11169 16902 11172
rect 16844 11163 16902 11169
rect 17218 11160 17224 11172
rect 17276 11160 17282 11212
rect 17402 11160 17408 11212
rect 17460 11200 17466 11212
rect 17460 11172 19288 11200
rect 17460 11160 17466 11172
rect 16255 11104 16528 11132
rect 16577 11135 16635 11141
rect 16255 11101 16267 11104
rect 16209 11095 16267 11101
rect 16577 11101 16589 11135
rect 16623 11101 16635 11135
rect 16577 11095 16635 11101
rect 8662 11024 8668 11076
rect 8720 11064 8726 11076
rect 8757 11067 8815 11073
rect 8757 11064 8769 11067
rect 8720 11036 8769 11064
rect 8720 11024 8726 11036
rect 8757 11033 8769 11036
rect 8803 11064 8815 11067
rect 8846 11064 8852 11076
rect 8803 11036 8852 11064
rect 8803 11033 8815 11036
rect 8757 11027 8815 11033
rect 8846 11024 8852 11036
rect 8904 11024 8910 11076
rect 13814 11024 13820 11076
rect 13872 11064 13878 11076
rect 15838 11064 15844 11076
rect 13872 11036 15844 11064
rect 13872 11024 13878 11036
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 12161 10999 12219 11005
rect 12161 10965 12173 10999
rect 12207 10996 12219 10999
rect 12250 10996 12256 11008
rect 12207 10968 12256 10996
rect 12207 10965 12219 10968
rect 12161 10959 12219 10965
rect 12250 10956 12256 10968
rect 12308 10956 12314 11008
rect 15562 10996 15568 11008
rect 15523 10968 15568 10996
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 16592 10996 16620 11095
rect 18598 11092 18604 11144
rect 18656 11132 18662 11144
rect 18966 11132 18972 11144
rect 18656 11104 18972 11132
rect 18656 11092 18662 11104
rect 18966 11092 18972 11104
rect 19024 11092 19030 11144
rect 19260 11141 19288 11172
rect 19702 11160 19708 11212
rect 19760 11200 19766 11212
rect 20165 11203 20223 11209
rect 20165 11200 20177 11203
rect 19760 11172 20177 11200
rect 19760 11160 19766 11172
rect 20165 11169 20177 11172
rect 20211 11169 20223 11203
rect 20272 11200 20300 11240
rect 20272 11172 20392 11200
rect 20165 11163 20223 11169
rect 19245 11135 19303 11141
rect 19245 11101 19257 11135
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19337 11135 19395 11141
rect 19337 11101 19349 11135
rect 19383 11101 19395 11135
rect 20254 11132 20260 11144
rect 20215 11104 20260 11132
rect 19337 11095 19395 11101
rect 19058 11024 19064 11076
rect 19116 11064 19122 11076
rect 19352 11064 19380 11095
rect 20254 11092 20260 11104
rect 20312 11092 20318 11144
rect 20364 11141 20392 11172
rect 20349 11135 20407 11141
rect 20349 11101 20361 11135
rect 20395 11101 20407 11135
rect 20349 11095 20407 11101
rect 19116 11036 19380 11064
rect 19116 11024 19122 11036
rect 16942 10996 16948 11008
rect 16592 10968 16948 10996
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 18782 10996 18788 11008
rect 18743 10968 18788 10996
rect 18782 10956 18788 10968
rect 18840 10956 18846 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 8481 10795 8539 10801
rect 8481 10761 8493 10795
rect 8527 10792 8539 10795
rect 8754 10792 8760 10804
rect 8527 10764 8760 10792
rect 8527 10761 8539 10764
rect 8481 10755 8539 10761
rect 8754 10752 8760 10764
rect 8812 10752 8818 10804
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 12342 10792 12348 10804
rect 12032 10764 12348 10792
rect 12032 10752 12038 10764
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 13265 10795 13323 10801
rect 12492 10764 12537 10792
rect 12492 10752 12498 10764
rect 13265 10761 13277 10795
rect 13311 10792 13323 10795
rect 14274 10792 14280 10804
rect 13311 10764 14280 10792
rect 13311 10761 13323 10764
rect 13265 10755 13323 10761
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 15289 10795 15347 10801
rect 15289 10761 15301 10795
rect 15335 10792 15347 10795
rect 17310 10792 17316 10804
rect 15335 10764 17316 10792
rect 15335 10761 15347 10764
rect 15289 10755 15347 10761
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 10597 10727 10655 10733
rect 10597 10693 10609 10727
rect 10643 10693 10655 10727
rect 10597 10687 10655 10693
rect 9030 10656 9036 10668
rect 8991 10628 9036 10656
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 8941 10591 8999 10597
rect 8941 10557 8953 10591
rect 8987 10588 8999 10591
rect 9122 10588 9128 10600
rect 8987 10560 9128 10588
rect 8987 10557 8999 10560
rect 8941 10551 8999 10557
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9493 10591 9551 10597
rect 9493 10557 9505 10591
rect 9539 10557 9551 10591
rect 10612 10588 10640 10687
rect 12618 10684 12624 10736
rect 12676 10724 12682 10736
rect 15194 10724 15200 10736
rect 12676 10696 15200 10724
rect 12676 10684 12682 10696
rect 15194 10684 15200 10696
rect 15252 10684 15258 10736
rect 11146 10656 11152 10668
rect 11107 10628 11152 10656
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 11882 10656 11888 10668
rect 11843 10628 11888 10656
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 12308 10628 13093 10656
rect 12308 10616 12314 10628
rect 13081 10625 13093 10628
rect 13127 10656 13139 10659
rect 13817 10659 13875 10665
rect 13817 10656 13829 10659
rect 13127 10628 13829 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13817 10625 13829 10628
rect 13863 10625 13875 10659
rect 13817 10619 13875 10625
rect 14921 10659 14979 10665
rect 14921 10625 14933 10659
rect 14967 10656 14979 10659
rect 15286 10656 15292 10668
rect 14967 10628 15292 10656
rect 14967 10625 14979 10628
rect 14921 10619 14979 10625
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 15979 10628 16436 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 11609 10591 11667 10597
rect 11609 10588 11621 10591
rect 10612 10560 11621 10588
rect 9493 10551 9551 10557
rect 11609 10557 11621 10560
rect 11655 10557 11667 10591
rect 11609 10551 11667 10557
rect 13725 10591 13783 10597
rect 13725 10557 13737 10591
rect 13771 10588 13783 10591
rect 14274 10588 14280 10600
rect 13771 10560 14280 10588
rect 13771 10557 13783 10560
rect 13725 10551 13783 10557
rect 8570 10480 8576 10532
rect 8628 10520 8634 10532
rect 9508 10520 9536 10551
rect 14274 10548 14280 10560
rect 14332 10548 14338 10600
rect 14737 10591 14795 10597
rect 14737 10557 14749 10591
rect 14783 10588 14795 10591
rect 14783 10560 15516 10588
rect 14783 10557 14795 10560
rect 14737 10551 14795 10557
rect 8628 10492 9536 10520
rect 9769 10523 9827 10529
rect 8628 10480 8634 10492
rect 9769 10489 9781 10523
rect 9815 10520 9827 10523
rect 14090 10520 14096 10532
rect 9815 10492 14096 10520
rect 9815 10489 9827 10492
rect 9769 10483 9827 10489
rect 14090 10480 14096 10492
rect 14148 10480 14154 10532
rect 14645 10523 14703 10529
rect 14645 10489 14657 10523
rect 14691 10520 14703 10523
rect 15194 10520 15200 10532
rect 14691 10492 15200 10520
rect 14691 10489 14703 10492
rect 14645 10483 14703 10489
rect 15194 10480 15200 10492
rect 15252 10480 15258 10532
rect 15488 10520 15516 10560
rect 15562 10548 15568 10600
rect 15620 10588 15626 10600
rect 15657 10591 15715 10597
rect 15657 10588 15669 10591
rect 15620 10560 15669 10588
rect 15620 10548 15626 10560
rect 15657 10557 15669 10560
rect 15703 10557 15715 10591
rect 15657 10551 15715 10557
rect 16301 10591 16359 10597
rect 16301 10557 16313 10591
rect 16347 10557 16359 10591
rect 16408 10588 16436 10628
rect 17954 10616 17960 10668
rect 18012 10656 18018 10668
rect 18049 10659 18107 10665
rect 18049 10656 18061 10659
rect 18012 10628 18061 10656
rect 18012 10616 18018 10628
rect 18049 10625 18061 10628
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10656 19303 10659
rect 19291 10628 19748 10656
rect 19291 10625 19303 10628
rect 19245 10619 19303 10625
rect 16574 10597 16580 10600
rect 16568 10588 16580 10597
rect 16408 10560 16580 10588
rect 16301 10551 16359 10557
rect 16568 10551 16580 10560
rect 16206 10520 16212 10532
rect 15488 10492 16212 10520
rect 16206 10480 16212 10492
rect 16264 10480 16270 10532
rect 16316 10520 16344 10551
rect 16574 10548 16580 10551
rect 16632 10548 16638 10600
rect 17862 10588 17868 10600
rect 17052 10560 17868 10588
rect 16666 10520 16672 10532
rect 16316 10492 16672 10520
rect 16666 10480 16672 10492
rect 16724 10520 16730 10532
rect 16942 10520 16948 10532
rect 16724 10492 16948 10520
rect 16724 10480 16730 10492
rect 16942 10480 16948 10492
rect 17000 10480 17006 10532
rect 8849 10455 8907 10461
rect 8849 10421 8861 10455
rect 8895 10452 8907 10455
rect 8938 10452 8944 10464
rect 8895 10424 8944 10452
rect 8895 10421 8907 10424
rect 8849 10415 8907 10421
rect 8938 10412 8944 10424
rect 8996 10412 9002 10464
rect 10962 10452 10968 10464
rect 10923 10424 10968 10452
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11112 10424 11157 10452
rect 11112 10412 11118 10424
rect 12618 10412 12624 10464
rect 12676 10452 12682 10464
rect 12805 10455 12863 10461
rect 12805 10452 12817 10455
rect 12676 10424 12817 10452
rect 12676 10412 12682 10424
rect 12805 10421 12817 10424
rect 12851 10421 12863 10455
rect 12805 10415 12863 10421
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13262 10452 13268 10464
rect 12943 10424 13268 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13262 10412 13268 10424
rect 13320 10452 13326 10464
rect 13538 10452 13544 10464
rect 13320 10424 13544 10452
rect 13320 10412 13326 10424
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 13633 10455 13691 10461
rect 13633 10421 13645 10455
rect 13679 10452 13691 10455
rect 13722 10452 13728 10464
rect 13679 10424 13728 10452
rect 13679 10421 13691 10424
rect 13633 10415 13691 10421
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 14277 10455 14335 10461
rect 14277 10452 14289 10455
rect 13872 10424 14289 10452
rect 13872 10412 13878 10424
rect 14277 10421 14289 10424
rect 14323 10421 14335 10455
rect 14277 10415 14335 10421
rect 15749 10455 15807 10461
rect 15749 10421 15761 10455
rect 15795 10452 15807 10455
rect 17052 10452 17080 10560
rect 17862 10548 17868 10560
rect 17920 10548 17926 10600
rect 18782 10548 18788 10600
rect 18840 10588 18846 10600
rect 18969 10591 19027 10597
rect 18969 10588 18981 10591
rect 18840 10560 18981 10588
rect 18840 10548 18846 10560
rect 18969 10557 18981 10560
rect 19015 10557 19027 10591
rect 18969 10551 19027 10557
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 19613 10591 19671 10597
rect 19613 10588 19625 10591
rect 19392 10560 19625 10588
rect 19392 10548 19398 10560
rect 19613 10557 19625 10560
rect 19659 10557 19671 10591
rect 19613 10551 19671 10557
rect 17126 10480 17132 10532
rect 17184 10520 17190 10532
rect 19061 10523 19119 10529
rect 19061 10520 19073 10523
rect 17184 10492 19073 10520
rect 17184 10480 17190 10492
rect 19061 10489 19073 10492
rect 19107 10489 19119 10523
rect 19720 10520 19748 10628
rect 19880 10523 19938 10529
rect 19880 10520 19892 10523
rect 19720 10492 19892 10520
rect 19061 10483 19119 10489
rect 19880 10489 19892 10492
rect 19926 10520 19938 10523
rect 20530 10520 20536 10532
rect 19926 10492 20536 10520
rect 19926 10489 19938 10492
rect 19880 10483 19938 10489
rect 20530 10480 20536 10492
rect 20588 10480 20594 10532
rect 17678 10452 17684 10464
rect 15795 10424 17080 10452
rect 17639 10424 17684 10452
rect 15795 10421 15807 10424
rect 15749 10415 15807 10421
rect 17678 10412 17684 10424
rect 17736 10412 17742 10464
rect 18601 10455 18659 10461
rect 18601 10421 18613 10455
rect 18647 10452 18659 10455
rect 18966 10452 18972 10464
rect 18647 10424 18972 10452
rect 18647 10421 18659 10424
rect 18601 10415 18659 10421
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 20622 10412 20628 10464
rect 20680 10452 20686 10464
rect 20993 10455 21051 10461
rect 20993 10452 21005 10455
rect 20680 10424 21005 10452
rect 20680 10412 20686 10424
rect 20993 10421 21005 10424
rect 21039 10421 21051 10455
rect 20993 10415 21051 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 10594 10208 10600 10260
rect 10652 10208 10658 10260
rect 11238 10208 11244 10260
rect 11296 10248 11302 10260
rect 11793 10251 11851 10257
rect 11793 10248 11805 10251
rect 11296 10220 11805 10248
rect 11296 10208 11302 10220
rect 11793 10217 11805 10220
rect 11839 10217 11851 10251
rect 11793 10211 11851 10217
rect 12345 10251 12403 10257
rect 12345 10217 12357 10251
rect 12391 10248 12403 10251
rect 13354 10248 13360 10260
rect 12391 10220 13360 10248
rect 12391 10217 12403 10220
rect 12345 10211 12403 10217
rect 7920 10183 7978 10189
rect 7920 10149 7932 10183
rect 7966 10180 7978 10183
rect 8662 10180 8668 10192
rect 7966 10152 8668 10180
rect 7966 10149 7978 10152
rect 7920 10143 7978 10149
rect 8662 10140 8668 10152
rect 8720 10140 8726 10192
rect 10612 10112 10640 10208
rect 10680 10183 10738 10189
rect 10680 10149 10692 10183
rect 10726 10180 10738 10183
rect 11146 10180 11152 10192
rect 10726 10152 11152 10180
rect 10726 10149 10738 10152
rect 10680 10143 10738 10149
rect 11146 10140 11152 10152
rect 11204 10140 11210 10192
rect 11808 10180 11836 10211
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 13814 10248 13820 10260
rect 13775 10220 13820 10248
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 14366 10248 14372 10260
rect 14327 10220 14372 10248
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 14829 10251 14887 10257
rect 14829 10217 14841 10251
rect 14875 10248 14887 10251
rect 15010 10248 15016 10260
rect 14875 10220 15016 10248
rect 14875 10217 14887 10220
rect 14829 10211 14887 10217
rect 15010 10208 15016 10220
rect 15068 10208 15074 10260
rect 15470 10208 15476 10260
rect 15528 10248 15534 10260
rect 15749 10251 15807 10257
rect 15749 10248 15761 10251
rect 15528 10220 15761 10248
rect 15528 10208 15534 10220
rect 15749 10217 15761 10220
rect 15795 10217 15807 10251
rect 17126 10248 17132 10260
rect 17087 10220 17132 10248
rect 15749 10211 15807 10217
rect 17126 10208 17132 10220
rect 17184 10208 17190 10260
rect 17586 10248 17592 10260
rect 17547 10220 17592 10248
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 18141 10251 18199 10257
rect 18141 10217 18153 10251
rect 18187 10248 18199 10251
rect 20254 10248 20260 10260
rect 18187 10220 20260 10248
rect 18187 10217 18199 10220
rect 18141 10211 18199 10217
rect 20254 10208 20260 10220
rect 20312 10208 20318 10260
rect 20530 10248 20536 10260
rect 20491 10220 20536 10248
rect 20530 10208 20536 10220
rect 20588 10208 20594 10260
rect 12250 10180 12256 10192
rect 11808 10152 12256 10180
rect 12250 10140 12256 10152
rect 12308 10180 12314 10192
rect 13173 10183 13231 10189
rect 13173 10180 13185 10183
rect 12308 10152 13185 10180
rect 12308 10140 12314 10152
rect 13173 10149 13185 10152
rect 13219 10149 13231 10183
rect 13173 10143 13231 10149
rect 14737 10183 14795 10189
rect 14737 10149 14749 10183
rect 14783 10180 14795 10183
rect 15102 10180 15108 10192
rect 14783 10152 15108 10180
rect 14783 10149 14795 10152
rect 14737 10143 14795 10149
rect 15102 10140 15108 10152
rect 15160 10140 15166 10192
rect 16669 10183 16727 10189
rect 16669 10149 16681 10183
rect 16715 10180 16727 10183
rect 16758 10180 16764 10192
rect 16715 10152 16764 10180
rect 16715 10149 16727 10152
rect 16669 10143 16727 10149
rect 16758 10140 16764 10152
rect 16816 10140 16822 10192
rect 18782 10140 18788 10192
rect 18840 10180 18846 10192
rect 19978 10180 19984 10192
rect 18840 10152 19984 10180
rect 18840 10140 18846 10152
rect 19978 10140 19984 10152
rect 20036 10180 20042 10192
rect 20622 10180 20628 10192
rect 20036 10152 20628 10180
rect 20036 10140 20042 10152
rect 20622 10140 20628 10152
rect 20680 10140 20686 10192
rect 12713 10115 12771 10121
rect 10612 10084 12296 10112
rect 7650 10044 7656 10056
rect 7611 10016 7656 10044
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 10410 10044 10416 10056
rect 10371 10016 10416 10044
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 12268 10044 12296 10084
rect 12713 10081 12725 10115
rect 12759 10112 12771 10115
rect 13725 10115 13783 10121
rect 12759 10084 13584 10112
rect 12759 10081 12771 10084
rect 12713 10075 12771 10081
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12268 10016 12817 10044
rect 12805 10013 12817 10016
rect 12851 10013 12863 10047
rect 12805 10007 12863 10013
rect 12989 10047 13047 10053
rect 12989 10013 13001 10047
rect 13035 10044 13047 10047
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 13035 10016 13185 10044
rect 13035 10013 13047 10016
rect 12989 10007 13047 10013
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 8754 9936 8760 9988
rect 8812 9976 8818 9988
rect 9214 9976 9220 9988
rect 8812 9948 9220 9976
rect 8812 9936 8818 9948
rect 9214 9936 9220 9948
rect 9272 9976 9278 9988
rect 13556 9976 13584 10084
rect 13725 10081 13737 10115
rect 13771 10112 13783 10115
rect 15657 10115 15715 10121
rect 13771 10084 15332 10112
rect 13771 10081 13783 10084
rect 13725 10075 13783 10081
rect 13630 10004 13636 10056
rect 13688 10044 13694 10056
rect 13909 10047 13967 10053
rect 13909 10044 13921 10047
rect 13688 10016 13921 10044
rect 13688 10004 13694 10016
rect 13909 10013 13921 10016
rect 13955 10013 13967 10047
rect 13909 10007 13967 10013
rect 14550 10004 14556 10056
rect 14608 10044 14614 10056
rect 14921 10047 14979 10053
rect 14921 10044 14933 10047
rect 14608 10016 14933 10044
rect 14608 10004 14614 10016
rect 14921 10013 14933 10016
rect 14967 10013 14979 10047
rect 14921 10007 14979 10013
rect 14366 9976 14372 9988
rect 9272 9948 10456 9976
rect 9272 9936 9278 9948
rect 9033 9911 9091 9917
rect 9033 9877 9045 9911
rect 9079 9908 9091 9911
rect 9122 9908 9128 9920
rect 9079 9880 9128 9908
rect 9079 9877 9091 9880
rect 9033 9871 9091 9877
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 10428 9908 10456 9948
rect 11339 9948 13492 9976
rect 13556 9948 14372 9976
rect 11339 9908 11367 9948
rect 10428 9880 11367 9908
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 13357 9911 13415 9917
rect 13357 9908 13369 9911
rect 12768 9880 13369 9908
rect 12768 9868 12774 9880
rect 13357 9877 13369 9880
rect 13403 9877 13415 9911
rect 13464 9908 13492 9948
rect 14366 9936 14372 9948
rect 14424 9936 14430 9988
rect 15304 9985 15332 10084
rect 15657 10081 15669 10115
rect 15703 10112 15715 10115
rect 16117 10115 16175 10121
rect 16117 10112 16129 10115
rect 15703 10084 16129 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 16117 10081 16129 10084
rect 16163 10081 16175 10115
rect 16117 10075 16175 10081
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10112 16451 10115
rect 16850 10112 16856 10124
rect 16439 10084 16856 10112
rect 16439 10081 16451 10084
rect 16393 10075 16451 10081
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 17497 10115 17555 10121
rect 17497 10081 17509 10115
rect 17543 10081 17555 10115
rect 18506 10112 18512 10124
rect 18467 10084 18512 10112
rect 17497 10075 17555 10081
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10013 15899 10047
rect 15841 10007 15899 10013
rect 15289 9979 15347 9985
rect 15289 9945 15301 9979
rect 15335 9945 15347 9979
rect 15289 9939 15347 9945
rect 15378 9936 15384 9988
rect 15436 9976 15442 9988
rect 15856 9976 15884 10007
rect 15436 9948 15884 9976
rect 15436 9936 15442 9948
rect 17512 9908 17540 10075
rect 18506 10072 18512 10084
rect 18564 10072 18570 10124
rect 19409 10115 19467 10121
rect 19409 10112 19421 10115
rect 19076 10084 19421 10112
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10013 17831 10047
rect 17773 10007 17831 10013
rect 17788 9976 17816 10007
rect 18414 10004 18420 10056
rect 18472 10044 18478 10056
rect 18601 10047 18659 10053
rect 18601 10044 18613 10047
rect 18472 10016 18613 10044
rect 18472 10004 18478 10016
rect 18601 10013 18613 10016
rect 18647 10013 18659 10047
rect 18782 10044 18788 10056
rect 18743 10016 18788 10044
rect 18601 10007 18659 10013
rect 18782 10004 18788 10016
rect 18840 10004 18846 10056
rect 19076 9988 19104 10084
rect 19409 10081 19421 10084
rect 19455 10081 19467 10115
rect 19409 10075 19467 10081
rect 19153 10047 19211 10053
rect 19153 10013 19165 10047
rect 19199 10013 19211 10047
rect 19153 10007 19211 10013
rect 19058 9976 19064 9988
rect 17788 9948 19064 9976
rect 19058 9936 19064 9948
rect 19116 9936 19122 9988
rect 13464 9880 17540 9908
rect 19168 9908 19196 10007
rect 19334 9908 19340 9920
rect 19168 9880 19340 9908
rect 13357 9871 13415 9877
rect 19334 9868 19340 9880
rect 19392 9868 19398 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 15933 9707 15991 9713
rect 15933 9704 15945 9707
rect 15344 9676 15945 9704
rect 15344 9664 15350 9676
rect 15933 9673 15945 9676
rect 15979 9673 15991 9707
rect 15933 9667 15991 9673
rect 17126 9664 17132 9716
rect 17184 9704 17190 9716
rect 17770 9704 17776 9716
rect 17184 9676 17776 9704
rect 17184 9664 17190 9676
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 18506 9664 18512 9716
rect 18564 9704 18570 9716
rect 18782 9704 18788 9716
rect 18564 9676 18788 9704
rect 18564 9664 18570 9676
rect 18782 9664 18788 9676
rect 18840 9664 18846 9716
rect 19334 9704 19340 9716
rect 18892 9676 19340 9704
rect 11146 9636 11152 9648
rect 11107 9608 11152 9636
rect 11146 9596 11152 9608
rect 11204 9596 11210 9648
rect 16206 9636 16212 9648
rect 16167 9608 16212 9636
rect 16206 9596 16212 9608
rect 16264 9596 16270 9648
rect 17954 9596 17960 9648
rect 18012 9636 18018 9648
rect 18049 9639 18107 9645
rect 18049 9636 18061 9639
rect 18012 9608 18061 9636
rect 18012 9596 18018 9608
rect 18049 9605 18061 9608
rect 18095 9605 18107 9639
rect 18049 9599 18107 9605
rect 18322 9596 18328 9648
rect 18380 9636 18386 9648
rect 18892 9636 18920 9676
rect 19334 9664 19340 9676
rect 19392 9664 19398 9716
rect 18380 9608 18920 9636
rect 18380 9596 18386 9608
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 8021 9571 8079 9577
rect 8021 9568 8033 9571
rect 7708 9540 8033 9568
rect 7708 9528 7714 9540
rect 8021 9537 8033 9540
rect 8067 9537 8079 9571
rect 16761 9571 16819 9577
rect 16761 9568 16773 9571
rect 8021 9531 8079 9537
rect 13464 9540 14688 9568
rect 8036 9500 8064 9531
rect 9769 9503 9827 9509
rect 9769 9500 9781 9503
rect 8036 9472 9781 9500
rect 9769 9469 9781 9472
rect 9815 9500 9827 9503
rect 10410 9500 10416 9512
rect 9815 9472 10416 9500
rect 9815 9469 9827 9472
rect 9769 9463 9827 9469
rect 10410 9460 10416 9472
rect 10468 9500 10474 9512
rect 12342 9500 12348 9512
rect 10468 9472 12348 9500
rect 10468 9460 10474 9472
rect 12342 9460 12348 9472
rect 12400 9500 12406 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12400 9472 12449 9500
rect 12400 9460 12406 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 12526 9460 12532 9512
rect 12584 9500 12590 9512
rect 13464 9500 13492 9540
rect 14660 9512 14688 9540
rect 15856 9540 16773 9568
rect 12584 9472 13492 9500
rect 12584 9460 12590 9472
rect 14182 9460 14188 9512
rect 14240 9500 14246 9512
rect 14277 9503 14335 9509
rect 14277 9500 14289 9503
rect 14240 9472 14289 9500
rect 14240 9460 14246 9472
rect 14277 9469 14289 9472
rect 14323 9469 14335 9503
rect 14277 9463 14335 9469
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9500 14519 9503
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 14507 9472 14565 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 14553 9469 14565 9472
rect 14599 9469 14611 9503
rect 14553 9463 14611 9469
rect 14642 9460 14648 9512
rect 14700 9460 14706 9512
rect 15286 9500 15292 9512
rect 14752 9472 15292 9500
rect 8288 9435 8346 9441
rect 8288 9401 8300 9435
rect 8334 9432 8346 9435
rect 9122 9432 9128 9444
rect 8334 9404 9128 9432
rect 8334 9401 8346 9404
rect 8288 9395 8346 9401
rect 9122 9392 9128 9404
rect 9180 9392 9186 9444
rect 10036 9435 10094 9441
rect 10036 9401 10048 9435
rect 10082 9432 10094 9435
rect 11238 9432 11244 9444
rect 10082 9404 11244 9432
rect 10082 9401 10094 9404
rect 10036 9395 10094 9401
rect 11238 9392 11244 9404
rect 11296 9392 11302 9444
rect 12704 9435 12762 9441
rect 12704 9401 12716 9435
rect 12750 9432 12762 9435
rect 14752 9432 14780 9472
rect 15286 9460 15292 9472
rect 15344 9460 15350 9512
rect 15856 9444 15884 9540
rect 16761 9537 16773 9540
rect 16807 9537 16819 9571
rect 16761 9531 16819 9537
rect 17218 9528 17224 9580
rect 17276 9568 17282 9580
rect 18601 9571 18659 9577
rect 18601 9568 18613 9571
rect 17276 9540 18613 9568
rect 17276 9528 17282 9540
rect 18601 9537 18613 9540
rect 18647 9537 18659 9571
rect 19337 9571 19395 9577
rect 19337 9568 19349 9571
rect 18601 9531 18659 9537
rect 18708 9540 19349 9568
rect 16022 9460 16028 9512
rect 16080 9500 16086 9512
rect 18708 9500 18736 9540
rect 19337 9537 19349 9540
rect 19383 9537 19395 9571
rect 20438 9568 20444 9580
rect 20399 9540 20444 9568
rect 19337 9531 19395 9537
rect 20438 9528 20444 9540
rect 20496 9528 20502 9580
rect 20622 9568 20628 9580
rect 20583 9540 20628 9568
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 16080 9472 18736 9500
rect 16080 9460 16086 9472
rect 18966 9460 18972 9512
rect 19024 9500 19030 9512
rect 19061 9503 19119 9509
rect 19061 9500 19073 9503
rect 19024 9472 19073 9500
rect 19024 9460 19030 9472
rect 19061 9469 19073 9472
rect 19107 9469 19119 9503
rect 19061 9463 19119 9469
rect 12750 9404 14780 9432
rect 14820 9435 14878 9441
rect 12750 9401 12762 9404
rect 12704 9395 12762 9401
rect 14820 9401 14832 9435
rect 14866 9432 14878 9435
rect 15838 9432 15844 9444
rect 14866 9404 15844 9432
rect 14866 9401 14878 9404
rect 14820 9395 14878 9401
rect 15838 9392 15844 9404
rect 15896 9392 15902 9444
rect 16482 9392 16488 9444
rect 16540 9432 16546 9444
rect 16669 9435 16727 9441
rect 16669 9432 16681 9435
rect 16540 9404 16681 9432
rect 16540 9392 16546 9404
rect 16669 9401 16681 9404
rect 16715 9401 16727 9435
rect 18414 9432 18420 9444
rect 18375 9404 18420 9432
rect 16669 9395 16727 9401
rect 18414 9392 18420 9404
rect 18472 9392 18478 9444
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 9272 9336 9413 9364
rect 9272 9324 9278 9336
rect 9401 9333 9413 9336
rect 9447 9333 9459 9367
rect 11422 9364 11428 9376
rect 11383 9336 11428 9364
rect 9401 9327 9459 9333
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 12066 9324 12072 9376
rect 12124 9364 12130 9376
rect 13538 9364 13544 9376
rect 12124 9336 13544 9364
rect 12124 9324 12130 9336
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 13630 9324 13636 9376
rect 13688 9364 13694 9376
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 13688 9336 13829 9364
rect 13688 9324 13694 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 14090 9364 14096 9376
rect 14051 9336 14096 9364
rect 13817 9327 13875 9333
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14461 9367 14519 9373
rect 14461 9333 14473 9367
rect 14507 9364 14519 9367
rect 15562 9364 15568 9376
rect 14507 9336 15568 9364
rect 14507 9333 14519 9336
rect 14461 9327 14519 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 16577 9367 16635 9373
rect 16577 9333 16589 9367
rect 16623 9364 16635 9367
rect 17402 9364 17408 9376
rect 16623 9336 17408 9364
rect 16623 9333 16635 9336
rect 16577 9327 16635 9333
rect 17402 9324 17408 9336
rect 17460 9364 17466 9376
rect 17586 9364 17592 9376
rect 17460 9336 17592 9364
rect 17460 9324 17466 9336
rect 17586 9324 17592 9336
rect 17644 9324 17650 9376
rect 18506 9364 18512 9376
rect 18467 9336 18512 9364
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 19886 9324 19892 9376
rect 19944 9364 19950 9376
rect 19981 9367 20039 9373
rect 19981 9364 19993 9367
rect 19944 9336 19993 9364
rect 19944 9324 19950 9336
rect 19981 9333 19993 9336
rect 20027 9333 20039 9367
rect 20346 9364 20352 9376
rect 20307 9336 20352 9364
rect 19981 9327 20039 9333
rect 20346 9324 20352 9336
rect 20404 9324 20410 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 8570 9160 8576 9172
rect 8531 9132 8576 9160
rect 8570 9120 8576 9132
rect 8628 9120 8634 9172
rect 8941 9163 8999 9169
rect 8941 9129 8953 9163
rect 8987 9160 8999 9163
rect 9674 9160 9680 9172
rect 8987 9132 9680 9160
rect 8987 9129 8999 9132
rect 8941 9123 8999 9129
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10410 9160 10416 9172
rect 10371 9132 10416 9160
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 10689 9163 10747 9169
rect 10689 9129 10701 9163
rect 10735 9160 10747 9163
rect 10962 9160 10968 9172
rect 10735 9132 10968 9160
rect 10735 9129 10747 9132
rect 10689 9123 10747 9129
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 11057 9163 11115 9169
rect 11057 9129 11069 9163
rect 11103 9160 11115 9163
rect 11422 9160 11428 9172
rect 11103 9132 11428 9160
rect 11103 9129 11115 9132
rect 11057 9123 11115 9129
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 11532 9132 15148 9160
rect 3418 9052 3424 9104
rect 3476 9092 3482 9104
rect 11532 9092 11560 9132
rect 3476 9064 11560 9092
rect 12161 9095 12219 9101
rect 3476 9052 3482 9064
rect 12161 9061 12173 9095
rect 12207 9092 12219 9095
rect 12526 9092 12532 9104
rect 12207 9064 12532 9092
rect 12207 9061 12219 9064
rect 12161 9055 12219 9061
rect 12526 9052 12532 9064
rect 12584 9052 12590 9104
rect 13072 9095 13130 9101
rect 13072 9061 13084 9095
rect 13118 9092 13130 9095
rect 13630 9092 13636 9104
rect 13118 9064 13636 9092
rect 13118 9061 13130 9064
rect 13072 9055 13130 9061
rect 13630 9052 13636 9064
rect 13688 9052 13694 9104
rect 15120 9092 15148 9132
rect 15194 9120 15200 9172
rect 15252 9160 15258 9172
rect 15289 9163 15347 9169
rect 15289 9160 15301 9163
rect 15252 9132 15301 9160
rect 15252 9120 15258 9132
rect 15289 9129 15301 9132
rect 15335 9129 15347 9163
rect 15289 9123 15347 9129
rect 15470 9120 15476 9172
rect 15528 9160 15534 9172
rect 15657 9163 15715 9169
rect 15657 9160 15669 9163
rect 15528 9132 15669 9160
rect 15528 9120 15534 9132
rect 15657 9129 15669 9132
rect 15703 9160 15715 9163
rect 17954 9160 17960 9172
rect 15703 9132 17960 9160
rect 15703 9129 15715 9132
rect 15657 9123 15715 9129
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 18417 9163 18475 9169
rect 18417 9129 18429 9163
rect 18463 9129 18475 9163
rect 18417 9123 18475 9129
rect 17304 9095 17362 9101
rect 15120 9064 17264 9092
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 9024 10655 9027
rect 10962 9024 10968 9036
rect 10643 8996 10968 9024
rect 10643 8993 10655 8996
rect 10597 8987 10655 8993
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 11146 9024 11152 9036
rect 11072 8996 11152 9024
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 9033 8959 9091 8965
rect 9033 8956 9045 8959
rect 8628 8928 9045 8956
rect 8628 8916 8634 8928
rect 9033 8925 9045 8928
rect 9079 8925 9091 8959
rect 9214 8956 9220 8968
rect 9175 8928 9220 8956
rect 9033 8919 9091 8925
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 11072 8956 11100 8996
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 12066 9024 12072 9036
rect 12027 8996 12072 9024
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 12342 8984 12348 9036
rect 12400 9024 12406 9036
rect 12805 9027 12863 9033
rect 12805 9024 12817 9027
rect 12400 8996 12817 9024
rect 12400 8984 12406 8996
rect 12805 8993 12817 8996
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 13538 8984 13544 9036
rect 13596 9024 13602 9036
rect 15930 9024 15936 9036
rect 13596 8996 15936 9024
rect 13596 8984 13602 8996
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 16942 9024 16948 9036
rect 16903 8996 16948 9024
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17236 9024 17264 9064
rect 17304 9061 17316 9095
rect 17350 9092 17362 9095
rect 17678 9092 17684 9104
rect 17350 9064 17684 9092
rect 17350 9061 17362 9064
rect 17304 9055 17362 9061
rect 17678 9052 17684 9064
rect 17736 9052 17742 9104
rect 18432 9092 18460 9123
rect 19242 9120 19248 9172
rect 19300 9160 19306 9172
rect 20349 9163 20407 9169
rect 20349 9160 20361 9163
rect 19300 9132 20361 9160
rect 19300 9120 19306 9132
rect 20349 9129 20361 9132
rect 20395 9129 20407 9163
rect 20349 9123 20407 9129
rect 18960 9095 19018 9101
rect 18960 9092 18972 9095
rect 18432 9064 18972 9092
rect 18960 9061 18972 9064
rect 19006 9092 19018 9095
rect 19794 9092 19800 9104
rect 19006 9064 19800 9092
rect 19006 9061 19018 9064
rect 18960 9055 19018 9061
rect 19794 9052 19800 9064
rect 19852 9052 19858 9104
rect 20070 9024 20076 9036
rect 17236 8996 20076 9024
rect 20070 8984 20076 8996
rect 20128 8984 20134 9036
rect 10704 8928 11100 8956
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 10704 8888 10732 8928
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 12253 8959 12311 8965
rect 11296 8928 11341 8956
rect 11296 8916 11302 8928
rect 12253 8925 12265 8959
rect 12299 8925 12311 8959
rect 12253 8919 12311 8925
rect 8260 8860 10732 8888
rect 8260 8848 8266 8860
rect 10778 8848 10784 8900
rect 10836 8888 10842 8900
rect 12268 8888 12296 8919
rect 15654 8916 15660 8968
rect 15712 8956 15718 8968
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 15712 8928 15761 8956
rect 15712 8916 15718 8928
rect 15749 8925 15761 8928
rect 15795 8925 15807 8959
rect 15749 8919 15807 8925
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 17037 8959 17095 8965
rect 15896 8928 15941 8956
rect 15896 8916 15902 8928
rect 17037 8925 17049 8959
rect 17083 8925 17095 8959
rect 17037 8919 17095 8925
rect 10836 8860 12296 8888
rect 10836 8848 10842 8860
rect 15562 8848 15568 8900
rect 15620 8888 15626 8900
rect 16666 8888 16672 8900
rect 15620 8860 16672 8888
rect 15620 8848 15626 8860
rect 16666 8848 16672 8860
rect 16724 8888 16730 8900
rect 16761 8891 16819 8897
rect 16761 8888 16773 8891
rect 16724 8860 16773 8888
rect 16724 8848 16730 8860
rect 16761 8857 16773 8860
rect 16807 8888 16819 8891
rect 17052 8888 17080 8919
rect 18322 8916 18328 8968
rect 18380 8956 18386 8968
rect 18693 8959 18751 8965
rect 18693 8956 18705 8959
rect 18380 8928 18705 8956
rect 18380 8916 18386 8928
rect 18693 8925 18705 8928
rect 18739 8925 18751 8959
rect 18693 8919 18751 8925
rect 16807 8860 17080 8888
rect 16807 8857 16819 8860
rect 16761 8851 16819 8857
rect 11698 8820 11704 8832
rect 11659 8792 11704 8820
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 14182 8820 14188 8832
rect 14095 8792 14188 8820
rect 14182 8780 14188 8792
rect 14240 8820 14246 8832
rect 14734 8820 14740 8832
rect 14240 8792 14740 8820
rect 14240 8780 14246 8792
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 15102 8780 15108 8832
rect 15160 8820 15166 8832
rect 16482 8820 16488 8832
rect 15160 8792 16488 8820
rect 15160 8780 15166 8792
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 17052 8820 17080 8860
rect 17770 8820 17776 8832
rect 17052 8792 17776 8820
rect 17770 8780 17776 8792
rect 17828 8820 17834 8832
rect 18340 8820 18368 8916
rect 17828 8792 18368 8820
rect 17828 8780 17834 8792
rect 19058 8780 19064 8832
rect 19116 8820 19122 8832
rect 20073 8823 20131 8829
rect 20073 8820 20085 8823
rect 19116 8792 20085 8820
rect 19116 8780 19122 8792
rect 20073 8789 20085 8792
rect 20119 8789 20131 8823
rect 20073 8783 20131 8789
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 8570 8616 8576 8628
rect 8531 8588 8576 8616
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 11333 8619 11391 8625
rect 11333 8616 11345 8619
rect 11112 8588 11345 8616
rect 11112 8576 11118 8588
rect 11333 8585 11345 8588
rect 11379 8585 11391 8619
rect 11333 8579 11391 8585
rect 14108 8588 15424 8616
rect 14108 8560 14136 8588
rect 10962 8508 10968 8560
rect 11020 8548 11026 8560
rect 12621 8551 12679 8557
rect 12621 8548 12633 8551
rect 11020 8520 12633 8548
rect 11020 8508 11026 8520
rect 12621 8517 12633 8520
rect 12667 8517 12679 8551
rect 14090 8548 14096 8560
rect 12621 8511 12679 8517
rect 12820 8520 14096 8548
rect 9122 8480 9128 8492
rect 9083 8452 9128 8480
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11164 8452 11897 8480
rect 11164 8424 11192 8452
rect 11885 8449 11897 8452
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8412 9091 8415
rect 9582 8412 9588 8424
rect 9079 8384 9588 8412
rect 9079 8381 9091 8384
rect 9033 8375 9091 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 10410 8412 10416 8424
rect 9723 8384 10416 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 10410 8372 10416 8384
rect 10468 8412 10474 8424
rect 10870 8412 10876 8424
rect 10468 8384 10876 8412
rect 10468 8372 10474 8384
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11146 8372 11152 8424
rect 11204 8372 11210 8424
rect 11698 8412 11704 8424
rect 11659 8384 11704 8412
rect 11698 8372 11704 8384
rect 11756 8372 11762 8424
rect 12820 8421 12848 8520
rect 14090 8508 14096 8520
rect 14148 8508 14154 8560
rect 14185 8551 14243 8557
rect 14185 8517 14197 8551
rect 14231 8517 14243 8551
rect 14185 8511 14243 8517
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 13725 8483 13783 8489
rect 13725 8480 13737 8483
rect 13688 8452 13737 8480
rect 13688 8440 13694 8452
rect 13725 8449 13737 8452
rect 13771 8449 13783 8483
rect 13725 8443 13783 8449
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8412 13599 8415
rect 14200 8412 14228 8511
rect 14734 8480 14740 8492
rect 14695 8452 14740 8480
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 13587 8384 14228 8412
rect 13587 8381 13599 8384
rect 13541 8375 13599 8381
rect 14274 8372 14280 8424
rect 14332 8412 14338 8424
rect 14553 8415 14611 8421
rect 14553 8412 14565 8415
rect 14332 8384 14565 8412
rect 14332 8372 14338 8384
rect 14553 8381 14565 8384
rect 14599 8412 14611 8415
rect 15286 8412 15292 8424
rect 14599 8384 15292 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 15286 8372 15292 8384
rect 15344 8372 15350 8424
rect 15396 8421 15424 8588
rect 15838 8576 15844 8628
rect 15896 8616 15902 8628
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 15896 8588 16957 8616
rect 15896 8576 15902 8588
rect 16945 8585 16957 8588
rect 16991 8585 17003 8619
rect 18598 8616 18604 8628
rect 16945 8579 17003 8585
rect 18432 8588 18604 8616
rect 15562 8480 15568 8492
rect 15523 8452 15568 8480
rect 15562 8440 15568 8452
rect 15620 8440 15626 8492
rect 16574 8440 16580 8492
rect 16632 8480 16638 8492
rect 16632 8452 18276 8480
rect 16632 8440 16638 8452
rect 15381 8415 15439 8421
rect 15381 8381 15393 8415
rect 15427 8381 15439 8415
rect 16942 8412 16948 8424
rect 15381 8375 15439 8381
rect 15764 8384 16948 8412
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 8941 8347 8999 8353
rect 8941 8344 8953 8347
rect 6972 8316 8953 8344
rect 6972 8304 6978 8316
rect 8941 8313 8953 8316
rect 8987 8313 8999 8347
rect 8941 8307 8999 8313
rect 9944 8347 10002 8353
rect 9944 8313 9956 8347
rect 9990 8344 10002 8347
rect 10778 8344 10784 8356
rect 9990 8316 10784 8344
rect 9990 8313 10002 8316
rect 9944 8307 10002 8313
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 11164 8344 11192 8372
rect 11072 8316 11192 8344
rect 11072 8285 11100 8316
rect 11238 8304 11244 8356
rect 11296 8344 11302 8356
rect 12066 8344 12072 8356
rect 11296 8316 12072 8344
rect 11296 8304 11302 8316
rect 12066 8304 12072 8316
rect 12124 8304 12130 8356
rect 13633 8347 13691 8353
rect 13633 8313 13645 8347
rect 13679 8344 13691 8347
rect 13722 8344 13728 8356
rect 13679 8316 13728 8344
rect 13679 8313 13691 8316
rect 13633 8307 13691 8313
rect 13722 8304 13728 8316
rect 13780 8304 13786 8356
rect 14366 8304 14372 8356
rect 14424 8344 14430 8356
rect 14645 8347 14703 8353
rect 14645 8344 14657 8347
rect 14424 8316 14657 8344
rect 14424 8304 14430 8316
rect 14645 8313 14657 8316
rect 14691 8344 14703 8347
rect 15010 8344 15016 8356
rect 14691 8316 15016 8344
rect 14691 8313 14703 8316
rect 14645 8307 14703 8313
rect 15010 8304 15016 8316
rect 15068 8304 15074 8356
rect 15764 8344 15792 8384
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 15212 8316 15792 8344
rect 15832 8347 15890 8353
rect 11057 8279 11115 8285
rect 11057 8245 11069 8279
rect 11103 8245 11115 8279
rect 11057 8239 11115 8245
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 11793 8279 11851 8285
rect 11793 8276 11805 8279
rect 11204 8248 11805 8276
rect 11204 8236 11210 8248
rect 11793 8245 11805 8248
rect 11839 8245 11851 8279
rect 13170 8276 13176 8288
rect 13131 8248 13176 8276
rect 11793 8239 11851 8245
rect 13170 8236 13176 8248
rect 13228 8236 13234 8288
rect 13262 8236 13268 8288
rect 13320 8276 13326 8288
rect 14274 8276 14280 8288
rect 13320 8248 14280 8276
rect 13320 8236 13326 8248
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 15212 8285 15240 8316
rect 15832 8313 15844 8347
rect 15878 8344 15890 8347
rect 16298 8344 16304 8356
rect 15878 8316 16304 8344
rect 15878 8313 15890 8316
rect 15832 8307 15890 8313
rect 16298 8304 16304 8316
rect 16356 8304 16362 8356
rect 18138 8344 18144 8356
rect 16408 8316 18144 8344
rect 15197 8279 15255 8285
rect 15197 8245 15209 8279
rect 15243 8245 15255 8279
rect 15197 8239 15255 8245
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 16408 8276 16436 8316
rect 18138 8304 18144 8316
rect 18196 8304 18202 8356
rect 18248 8344 18276 8452
rect 18432 8412 18460 8588
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 19521 8551 19579 8557
rect 19521 8517 19533 8551
rect 19567 8548 19579 8551
rect 19794 8548 19800 8560
rect 19567 8520 19800 8548
rect 19567 8517 19579 8520
rect 19521 8511 19579 8517
rect 19794 8508 19800 8520
rect 19852 8508 19858 8560
rect 18598 8480 18604 8492
rect 18559 8452 18604 8480
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 20070 8480 20076 8492
rect 20031 8452 20076 8480
rect 20070 8440 20076 8452
rect 20128 8440 20134 8492
rect 18509 8415 18567 8421
rect 18509 8412 18521 8415
rect 18432 8384 18521 8412
rect 18509 8381 18521 8384
rect 18555 8381 18567 8415
rect 19886 8412 19892 8424
rect 19847 8384 19892 8412
rect 18509 8375 18567 8381
rect 19886 8372 19892 8384
rect 19944 8372 19950 8424
rect 18417 8347 18475 8353
rect 18417 8344 18429 8347
rect 18248 8316 18429 8344
rect 18417 8313 18429 8316
rect 18463 8313 18475 8347
rect 18417 8307 18475 8313
rect 17218 8276 17224 8288
rect 15344 8248 16436 8276
rect 17179 8248 17224 8276
rect 15344 8236 15350 8248
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 17954 8236 17960 8288
rect 18012 8276 18018 8288
rect 18049 8279 18107 8285
rect 18049 8276 18061 8279
rect 18012 8248 18061 8276
rect 18012 8236 18018 8248
rect 18049 8245 18061 8248
rect 18095 8245 18107 8279
rect 18049 8239 18107 8245
rect 19978 8236 19984 8288
rect 20036 8276 20042 8288
rect 20036 8248 20081 8276
rect 20036 8236 20042 8248
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 10137 8075 10195 8081
rect 10137 8041 10149 8075
rect 10183 8072 10195 8075
rect 11146 8072 11152 8084
rect 10183 8044 11152 8072
rect 10183 8041 10195 8044
rect 10137 8035 10195 8041
rect 11146 8032 11152 8044
rect 11204 8032 11210 8084
rect 14921 8075 14979 8081
rect 14921 8072 14933 8075
rect 13648 8044 14933 8072
rect 13648 8016 13676 8044
rect 14921 8041 14933 8044
rect 14967 8041 14979 8075
rect 18046 8072 18052 8084
rect 14921 8035 14979 8041
rect 15948 8044 18052 8072
rect 10505 8007 10563 8013
rect 10505 7973 10517 8007
rect 10551 8004 10563 8007
rect 11416 8007 11474 8013
rect 10551 7976 11284 8004
rect 10551 7973 10563 7976
rect 10505 7967 10563 7973
rect 8849 7939 8907 7945
rect 8849 7905 8861 7939
rect 8895 7936 8907 7939
rect 9674 7936 9680 7948
rect 8895 7908 9680 7936
rect 8895 7905 8907 7908
rect 8849 7899 8907 7905
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 10597 7939 10655 7945
rect 10597 7905 10609 7939
rect 10643 7936 10655 7939
rect 11054 7936 11060 7948
rect 10643 7908 11060 7936
rect 10643 7905 10655 7908
rect 10597 7899 10655 7905
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 11256 7936 11284 7976
rect 11416 7973 11428 8007
rect 11462 8004 11474 8007
rect 13630 8004 13636 8016
rect 11462 7976 13636 8004
rect 11462 7973 11474 7976
rect 11416 7967 11474 7973
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 13808 8007 13866 8013
rect 13808 7973 13820 8007
rect 13854 8004 13866 8007
rect 14182 8004 14188 8016
rect 13854 7976 14188 8004
rect 13854 7973 13866 7976
rect 13808 7967 13866 7973
rect 14182 7964 14188 7976
rect 14240 7964 14246 8016
rect 14090 7936 14096 7948
rect 11256 7908 14096 7936
rect 14090 7896 14096 7908
rect 14148 7936 14154 7948
rect 15948 7936 15976 8044
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 20070 8032 20076 8084
rect 20128 8072 20134 8084
rect 20257 8075 20315 8081
rect 20257 8072 20269 8075
rect 20128 8044 20269 8072
rect 20128 8032 20134 8044
rect 20257 8041 20269 8044
rect 20303 8041 20315 8075
rect 20257 8035 20315 8041
rect 20346 8032 20352 8084
rect 20404 8072 20410 8084
rect 20901 8075 20959 8081
rect 20901 8072 20913 8075
rect 20404 8044 20913 8072
rect 20404 8032 20410 8044
rect 20901 8041 20913 8044
rect 20947 8041 20959 8075
rect 20901 8035 20959 8041
rect 16936 8007 16994 8013
rect 16936 7973 16948 8007
rect 16982 8004 16994 8007
rect 18598 8004 18604 8016
rect 16982 7976 18604 8004
rect 16982 7973 16994 7976
rect 16936 7967 16994 7973
rect 18598 7964 18604 7976
rect 18656 7964 18662 8016
rect 14148 7908 15976 7936
rect 16025 7939 16083 7945
rect 14148 7896 14154 7908
rect 16025 7905 16037 7939
rect 16071 7936 16083 7939
rect 16758 7936 16764 7948
rect 16071 7908 16764 7936
rect 16071 7905 16083 7908
rect 16025 7899 16083 7905
rect 16758 7896 16764 7908
rect 16816 7896 16822 7948
rect 17770 7896 17776 7948
rect 17828 7936 17834 7948
rect 18877 7939 18935 7945
rect 18877 7936 18889 7939
rect 17828 7908 18889 7936
rect 17828 7896 17834 7908
rect 18877 7905 18889 7908
rect 18923 7905 18935 7939
rect 18877 7899 18935 7905
rect 19144 7939 19202 7945
rect 19144 7905 19156 7939
rect 19190 7936 19202 7939
rect 20622 7936 20628 7948
rect 19190 7908 20628 7936
rect 19190 7905 19202 7908
rect 19144 7899 19202 7905
rect 20622 7896 20628 7908
rect 20680 7896 20686 7948
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7868 9183 7871
rect 10778 7868 10784 7880
rect 9171 7840 10088 7868
rect 10739 7840 10784 7868
rect 9171 7837 9183 7840
rect 9125 7831 9183 7837
rect 10060 7732 10088 7840
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 10870 7828 10876 7880
rect 10928 7868 10934 7880
rect 11149 7871 11207 7877
rect 11149 7868 11161 7871
rect 10928 7840 11161 7868
rect 10928 7828 10934 7840
rect 11149 7837 11161 7840
rect 11195 7837 11207 7871
rect 13538 7868 13544 7880
rect 13499 7840 13544 7868
rect 11149 7831 11207 7837
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 16117 7871 16175 7877
rect 16117 7837 16129 7871
rect 16163 7837 16175 7871
rect 16298 7868 16304 7880
rect 16259 7840 16304 7868
rect 16117 7831 16175 7837
rect 11790 7732 11796 7744
rect 10060 7704 11796 7732
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 12066 7692 12072 7744
rect 12124 7732 12130 7744
rect 12529 7735 12587 7741
rect 12529 7732 12541 7735
rect 12124 7704 12541 7732
rect 12124 7692 12130 7704
rect 12529 7701 12541 7704
rect 12575 7701 12587 7735
rect 12529 7695 12587 7701
rect 13262 7692 13268 7744
rect 13320 7732 13326 7744
rect 15657 7735 15715 7741
rect 15657 7732 15669 7735
rect 13320 7704 15669 7732
rect 13320 7692 13326 7704
rect 15657 7701 15669 7704
rect 15703 7701 15715 7735
rect 16132 7732 16160 7831
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 16666 7868 16672 7880
rect 16627 7840 16672 7868
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 17770 7732 17776 7744
rect 16132 7704 17776 7732
rect 15657 7695 15715 7701
rect 17770 7692 17776 7704
rect 17828 7692 17834 7744
rect 17862 7692 17868 7744
rect 17920 7732 17926 7744
rect 18049 7735 18107 7741
rect 18049 7732 18061 7735
rect 17920 7704 18061 7732
rect 17920 7692 17926 7704
rect 18049 7701 18061 7704
rect 18095 7701 18107 7735
rect 18049 7695 18107 7701
rect 18782 7692 18788 7744
rect 18840 7732 18846 7744
rect 19058 7732 19064 7744
rect 18840 7704 19064 7732
rect 18840 7692 18846 7704
rect 19058 7692 19064 7704
rect 19116 7692 19122 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 9306 7488 9312 7540
rect 9364 7528 9370 7540
rect 10505 7531 10563 7537
rect 9364 7500 10456 7528
rect 9364 7488 9370 7500
rect 10428 7460 10456 7500
rect 10505 7497 10517 7531
rect 10551 7528 10563 7531
rect 10778 7528 10784 7540
rect 10551 7500 10784 7528
rect 10551 7497 10563 7500
rect 10505 7491 10563 7497
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 13464 7500 16243 7528
rect 10428 7432 12296 7460
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12066 7392 12072 7404
rect 12023 7364 12072 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12268 7392 12296 7432
rect 13464 7392 13492 7500
rect 13538 7420 13544 7472
rect 13596 7460 13602 7472
rect 15194 7460 15200 7472
rect 13596 7432 15200 7460
rect 13596 7420 13602 7432
rect 15194 7420 15200 7432
rect 15252 7460 15258 7472
rect 16215 7460 16243 7500
rect 16298 7488 16304 7540
rect 16356 7528 16362 7540
rect 16669 7531 16727 7537
rect 16669 7528 16681 7531
rect 16356 7500 16681 7528
rect 16356 7488 16362 7500
rect 16669 7497 16681 7500
rect 16715 7497 16727 7531
rect 16669 7491 16727 7497
rect 16758 7488 16764 7540
rect 16816 7528 16822 7540
rect 16945 7531 17003 7537
rect 16945 7528 16957 7531
rect 16816 7500 16957 7528
rect 16816 7488 16822 7500
rect 16945 7497 16957 7500
rect 16991 7497 17003 7531
rect 16945 7491 17003 7497
rect 17770 7488 17776 7540
rect 17828 7528 17834 7540
rect 18049 7531 18107 7537
rect 18049 7528 18061 7531
rect 17828 7500 18061 7528
rect 17828 7488 17834 7500
rect 18049 7497 18061 7500
rect 18095 7497 18107 7531
rect 18049 7491 18107 7497
rect 19978 7488 19984 7540
rect 20036 7528 20042 7540
rect 20073 7531 20131 7537
rect 20073 7528 20085 7531
rect 20036 7500 20085 7528
rect 20036 7488 20042 7500
rect 20073 7497 20085 7500
rect 20119 7497 20131 7531
rect 20073 7491 20131 7497
rect 17402 7460 17408 7472
rect 15252 7432 15332 7460
rect 16215 7432 17408 7460
rect 15252 7420 15258 7432
rect 12268 7364 13492 7392
rect 13630 7352 13636 7404
rect 13688 7392 13694 7404
rect 13725 7395 13783 7401
rect 13725 7392 13737 7395
rect 13688 7364 13737 7392
rect 13688 7352 13694 7364
rect 13725 7361 13737 7364
rect 13771 7361 13783 7395
rect 13725 7355 13783 7361
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 15304 7401 15332 7432
rect 17402 7420 17408 7432
rect 17460 7460 17466 7472
rect 17460 7432 19748 7460
rect 17460 7420 17466 7432
rect 14737 7395 14795 7401
rect 14737 7392 14749 7395
rect 14240 7364 14749 7392
rect 14240 7352 14246 7364
rect 14737 7361 14749 7364
rect 14783 7361 14795 7395
rect 14737 7355 14795 7361
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7361 15347 7395
rect 17497 7395 17555 7401
rect 17497 7392 17509 7395
rect 15289 7355 15347 7361
rect 17144 7364 17509 7392
rect 9122 7324 9128 7336
rect 9083 7296 9128 7324
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 11793 7327 11851 7333
rect 11793 7293 11805 7327
rect 11839 7324 11851 7327
rect 13170 7324 13176 7336
rect 11839 7296 13176 7324
rect 11839 7293 11851 7296
rect 11793 7287 11851 7293
rect 13170 7284 13176 7296
rect 13228 7284 13234 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 13872 7296 14657 7324
rect 13872 7284 13878 7296
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 14645 7287 14703 7293
rect 15556 7327 15614 7333
rect 15556 7293 15568 7327
rect 15602 7324 15614 7327
rect 17144 7324 17172 7364
rect 17497 7361 17509 7364
rect 17543 7392 17555 7395
rect 17862 7392 17868 7404
rect 17543 7364 17868 7392
rect 17543 7361 17555 7364
rect 17497 7355 17555 7361
rect 17862 7352 17868 7364
rect 17920 7392 17926 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 17920 7364 18613 7392
rect 17920 7352 17926 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 18690 7352 18696 7404
rect 18748 7392 18754 7404
rect 19613 7395 19671 7401
rect 19613 7392 19625 7395
rect 18748 7364 19625 7392
rect 18748 7352 18754 7364
rect 19613 7361 19625 7364
rect 19659 7361 19671 7395
rect 19613 7355 19671 7361
rect 15602 7296 17172 7324
rect 15602 7293 15614 7296
rect 15556 7287 15614 7293
rect 17218 7284 17224 7336
rect 17276 7324 17282 7336
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 17276 7296 17325 7324
rect 17276 7284 17282 7296
rect 17313 7293 17325 7296
rect 17359 7293 17371 7327
rect 17313 7287 17371 7293
rect 17405 7327 17463 7333
rect 17405 7293 17417 7327
rect 17451 7324 17463 7327
rect 17954 7324 17960 7336
rect 17451 7296 17960 7324
rect 17451 7293 17463 7296
rect 17405 7287 17463 7293
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 18506 7284 18512 7336
rect 18564 7324 18570 7336
rect 19426 7324 19432 7336
rect 18564 7296 19288 7324
rect 19387 7296 19432 7324
rect 18564 7284 18570 7296
rect 9398 7265 9404 7268
rect 9392 7256 9404 7265
rect 9359 7228 9404 7256
rect 9392 7219 9404 7228
rect 9398 7216 9404 7219
rect 9456 7216 9462 7268
rect 11701 7259 11759 7265
rect 11701 7225 11713 7259
rect 11747 7256 11759 7259
rect 12713 7259 12771 7265
rect 11747 7228 12480 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7188 11391 7191
rect 12250 7188 12256 7200
rect 11379 7160 12256 7188
rect 11379 7157 11391 7160
rect 11333 7151 11391 7157
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 12452 7188 12480 7228
rect 12713 7225 12725 7259
rect 12759 7256 12771 7259
rect 13541 7259 13599 7265
rect 13541 7256 13553 7259
rect 12759 7228 13553 7256
rect 12759 7225 12771 7228
rect 12713 7219 12771 7225
rect 13541 7225 13553 7228
rect 13587 7225 13599 7259
rect 13541 7219 13599 7225
rect 13906 7216 13912 7268
rect 13964 7256 13970 7268
rect 14553 7259 14611 7265
rect 14553 7256 14565 7259
rect 13964 7228 14565 7256
rect 13964 7216 13970 7228
rect 14553 7225 14565 7228
rect 14599 7256 14611 7259
rect 16574 7256 16580 7268
rect 14599 7228 16580 7256
rect 14599 7225 14611 7228
rect 14553 7219 14611 7225
rect 16574 7216 16580 7228
rect 16632 7216 16638 7268
rect 18417 7259 18475 7265
rect 18417 7225 18429 7259
rect 18463 7256 18475 7259
rect 18463 7228 19104 7256
rect 18463 7225 18475 7228
rect 18417 7219 18475 7225
rect 13173 7191 13231 7197
rect 13173 7188 13185 7191
rect 12452 7160 13185 7188
rect 13173 7157 13185 7160
rect 13219 7157 13231 7191
rect 13173 7151 13231 7157
rect 13633 7191 13691 7197
rect 13633 7157 13645 7191
rect 13679 7188 13691 7191
rect 14185 7191 14243 7197
rect 14185 7188 14197 7191
rect 13679 7160 14197 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 14185 7157 14197 7160
rect 14231 7157 14243 7191
rect 18506 7188 18512 7200
rect 18467 7160 18512 7188
rect 14185 7151 14243 7157
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 19076 7197 19104 7228
rect 19260 7200 19288 7296
rect 19426 7284 19432 7296
rect 19484 7284 19490 7336
rect 19720 7324 19748 7432
rect 20622 7392 20628 7404
rect 20583 7364 20628 7392
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 20533 7327 20591 7333
rect 20533 7324 20545 7327
rect 19720 7296 20545 7324
rect 20533 7293 20545 7296
rect 20579 7293 20591 7327
rect 20533 7287 20591 7293
rect 19061 7191 19119 7197
rect 19061 7157 19073 7191
rect 19107 7157 19119 7191
rect 19061 7151 19119 7157
rect 19242 7148 19248 7200
rect 19300 7188 19306 7200
rect 19521 7191 19579 7197
rect 19521 7188 19533 7191
rect 19300 7160 19533 7188
rect 19300 7148 19306 7160
rect 19521 7157 19533 7160
rect 19567 7157 19579 7191
rect 20438 7188 20444 7200
rect 20399 7160 20444 7188
rect 19521 7151 19579 7157
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 9674 6984 9680 6996
rect 9635 6956 9680 6984
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 14093 6987 14151 6993
rect 14093 6953 14105 6987
rect 14139 6984 14151 6987
rect 14366 6984 14372 6996
rect 14139 6956 14372 6984
rect 14139 6953 14151 6956
rect 14093 6947 14151 6953
rect 14366 6944 14372 6956
rect 14424 6984 14430 6996
rect 18509 6987 18567 6993
rect 14424 6956 15792 6984
rect 14424 6944 14430 6956
rect 9122 6916 9128 6928
rect 8128 6888 9128 6916
rect 8128 6848 8156 6888
rect 9122 6876 9128 6888
rect 9180 6876 9186 6928
rect 11784 6919 11842 6925
rect 10796 6888 11100 6916
rect 7944 6820 8156 6848
rect 8196 6851 8254 6857
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 7944 6789 7972 6820
rect 8196 6817 8208 6851
rect 8242 6848 8254 6851
rect 9030 6848 9036 6860
rect 8242 6820 9036 6848
rect 8242 6817 8254 6820
rect 8196 6811 8254 6817
rect 9030 6808 9036 6820
rect 9088 6808 9094 6860
rect 10042 6848 10048 6860
rect 10003 6820 10048 6848
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10796 6848 10824 6888
rect 10962 6848 10968 6860
rect 10376 6820 10824 6848
rect 10923 6820 10968 6848
rect 10376 6808 10382 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11072 6848 11100 6888
rect 11784 6885 11796 6919
rect 11830 6916 11842 6919
rect 12066 6916 12072 6928
rect 11830 6888 12072 6916
rect 11830 6885 11842 6888
rect 11784 6879 11842 6885
rect 12066 6876 12072 6888
rect 12124 6876 12130 6928
rect 15378 6876 15384 6928
rect 15436 6916 15442 6928
rect 15657 6919 15715 6925
rect 15657 6916 15669 6919
rect 15436 6888 15669 6916
rect 15436 6876 15442 6888
rect 15657 6885 15669 6888
rect 15703 6885 15715 6919
rect 15764 6916 15792 6956
rect 18509 6953 18521 6987
rect 18555 6984 18567 6987
rect 18598 6984 18604 6996
rect 18555 6956 18604 6984
rect 18555 6953 18567 6956
rect 18509 6947 18567 6953
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 20533 6987 20591 6993
rect 20533 6953 20545 6987
rect 20579 6984 20591 6987
rect 20622 6984 20628 6996
rect 20579 6956 20628 6984
rect 20579 6953 20591 6956
rect 20533 6947 20591 6953
rect 20622 6944 20628 6956
rect 20680 6944 20686 6996
rect 19886 6916 19892 6928
rect 15764 6888 19892 6916
rect 15657 6879 15715 6885
rect 19886 6876 19892 6888
rect 19944 6876 19950 6928
rect 13446 6848 13452 6860
rect 11072 6820 13452 6848
rect 13446 6808 13452 6820
rect 13504 6808 13510 6860
rect 13998 6808 14004 6860
rect 14056 6808 14062 6860
rect 14185 6851 14243 6857
rect 14185 6817 14197 6851
rect 14231 6848 14243 6851
rect 14458 6848 14464 6860
rect 14231 6820 14464 6848
rect 14231 6817 14243 6820
rect 14185 6811 14243 6817
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 16942 6848 16948 6860
rect 16903 6820 16948 6848
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 17396 6851 17454 6857
rect 17396 6817 17408 6851
rect 17442 6848 17454 6851
rect 18690 6848 18696 6860
rect 17442 6820 18696 6848
rect 17442 6817 17454 6820
rect 17396 6811 17454 6817
rect 18690 6808 18696 6820
rect 18748 6808 18754 6860
rect 19426 6857 19432 6860
rect 19420 6848 19432 6857
rect 19387 6820 19432 6848
rect 19420 6811 19432 6820
rect 19426 6808 19432 6811
rect 19484 6808 19490 6860
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7708 6752 7941 6780
rect 7708 6740 7714 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 7929 6743 7987 6749
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 10229 6743 10287 6749
rect 10888 6752 11529 6780
rect 9309 6715 9367 6721
rect 9309 6681 9321 6715
rect 9355 6712 9367 6715
rect 9398 6712 9404 6724
rect 9355 6684 9404 6712
rect 9355 6681 9367 6684
rect 9309 6675 9367 6681
rect 9398 6672 9404 6684
rect 9456 6712 9462 6724
rect 10244 6712 10272 6743
rect 9456 6684 10272 6712
rect 9456 6672 9462 6684
rect 10888 6656 10916 6752
rect 11517 6749 11529 6752
rect 11563 6749 11575 6783
rect 14016 6780 14044 6808
rect 11517 6743 11575 6749
rect 12820 6752 14044 6780
rect 9122 6604 9128 6656
rect 9180 6644 9186 6656
rect 10781 6647 10839 6653
rect 10781 6644 10793 6647
rect 9180 6616 10793 6644
rect 9180 6604 9186 6616
rect 10781 6613 10793 6616
rect 10827 6644 10839 6647
rect 10870 6644 10876 6656
rect 10827 6616 10876 6644
rect 10827 6613 10839 6616
rect 10781 6607 10839 6613
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 12820 6644 12848 6752
rect 14274 6740 14280 6792
rect 14332 6780 14338 6792
rect 14332 6752 14377 6780
rect 14332 6740 14338 6752
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 15344 6752 15761 6780
rect 15344 6740 15350 6752
rect 15749 6749 15761 6752
rect 15795 6749 15807 6783
rect 15930 6780 15936 6792
rect 15891 6752 15936 6780
rect 15749 6743 15807 6749
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 16298 6780 16304 6792
rect 16259 6752 16304 6780
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 17129 6783 17187 6789
rect 17129 6749 17141 6783
rect 17175 6749 17187 6783
rect 19153 6783 19211 6789
rect 19153 6780 19165 6783
rect 17129 6743 17187 6749
rect 18524 6752 19165 6780
rect 13722 6712 13728 6724
rect 13683 6684 13728 6712
rect 13722 6672 13728 6684
rect 13780 6672 13786 6724
rect 15194 6672 15200 6724
rect 15252 6712 15258 6724
rect 16761 6715 16819 6721
rect 16761 6712 16773 6715
rect 15252 6684 16773 6712
rect 15252 6672 15258 6684
rect 16761 6681 16773 6684
rect 16807 6712 16819 6715
rect 17144 6712 17172 6743
rect 16807 6684 17172 6712
rect 16807 6681 16819 6684
rect 16761 6675 16819 6681
rect 11020 6616 12848 6644
rect 12897 6647 12955 6653
rect 11020 6604 11026 6616
rect 12897 6613 12909 6647
rect 12943 6644 12955 6647
rect 14090 6644 14096 6656
rect 12943 6616 14096 6644
rect 12943 6613 12955 6616
rect 12897 6607 12955 6613
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 15289 6647 15347 6653
rect 15289 6613 15301 6647
rect 15335 6644 15347 6647
rect 16114 6644 16120 6656
rect 15335 6616 16120 6644
rect 15335 6613 15347 6616
rect 15289 6607 15347 6613
rect 16114 6604 16120 6616
rect 16172 6604 16178 6656
rect 17144 6644 17172 6684
rect 18524 6644 18552 6752
rect 19153 6749 19165 6752
rect 19199 6749 19211 6783
rect 19153 6743 19211 6749
rect 17144 6616 18552 6644
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 9030 6440 9036 6452
rect 8991 6412 9036 6440
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 10042 6440 10048 6452
rect 9355 6412 10048 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 10192 6412 10333 6440
rect 10192 6400 10198 6412
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 10321 6403 10379 6409
rect 10962 6400 10968 6452
rect 11020 6400 11026 6452
rect 11054 6400 11060 6452
rect 11112 6440 11118 6452
rect 13538 6440 13544 6452
rect 11112 6412 13544 6440
rect 11112 6400 11118 6412
rect 13538 6400 13544 6412
rect 13596 6400 13602 6452
rect 15286 6440 15292 6452
rect 15247 6412 15292 6440
rect 15286 6400 15292 6412
rect 15344 6400 15350 6452
rect 16390 6400 16396 6452
rect 16448 6440 16454 6452
rect 18049 6443 18107 6449
rect 16448 6412 17172 6440
rect 16448 6400 16454 6412
rect 6086 6264 6092 6316
rect 6144 6304 6150 6316
rect 9048 6304 9076 6400
rect 10226 6332 10232 6384
rect 10284 6372 10290 6384
rect 10980 6372 11008 6400
rect 10284 6344 11008 6372
rect 10284 6332 10290 6344
rect 12066 6332 12072 6384
rect 12124 6372 12130 6384
rect 12434 6372 12440 6384
rect 12124 6344 12440 6372
rect 12124 6332 12130 6344
rect 12434 6332 12440 6344
rect 12492 6372 12498 6384
rect 17144 6372 17172 6412
rect 18049 6409 18061 6443
rect 18095 6440 18107 6443
rect 18506 6440 18512 6452
rect 18095 6412 18512 6440
rect 18095 6409 18107 6412
rect 18049 6403 18107 6409
rect 18506 6400 18512 6412
rect 18564 6400 18570 6452
rect 20714 6372 20720 6384
rect 12492 6344 16979 6372
rect 17144 6344 20720 6372
rect 12492 6332 12498 6344
rect 9861 6307 9919 6313
rect 9861 6304 9873 6307
rect 6144 6276 7788 6304
rect 9048 6276 9873 6304
rect 6144 6264 6150 6276
rect 7650 6236 7656 6248
rect 7611 6208 7656 6236
rect 7650 6196 7656 6208
rect 7708 6196 7714 6248
rect 7760 6236 7788 6276
rect 9861 6273 9873 6276
rect 9907 6304 9919 6307
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 9907 6276 10885 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11020 6276 11897 6304
rect 11020 6264 11026 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 12986 6304 12992 6316
rect 12947 6276 12992 6304
rect 11885 6267 11943 6273
rect 12986 6264 12992 6276
rect 13044 6264 13050 6316
rect 14090 6304 14096 6316
rect 14051 6276 14096 6304
rect 14090 6264 14096 6276
rect 14148 6264 14154 6316
rect 15470 6264 15476 6316
rect 15528 6304 15534 6316
rect 15841 6307 15899 6313
rect 15841 6304 15853 6307
rect 15528 6276 15853 6304
rect 15528 6264 15534 6276
rect 15841 6273 15853 6276
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 15930 6264 15936 6316
rect 15988 6304 15994 6316
rect 16482 6304 16488 6316
rect 15988 6276 16488 6304
rect 15988 6264 15994 6276
rect 16482 6264 16488 6276
rect 16540 6304 16546 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16540 6276 16865 6304
rect 16540 6264 16546 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 11701 6239 11759 6245
rect 7760 6208 11468 6236
rect 7742 6128 7748 6180
rect 7800 6168 7806 6180
rect 7898 6171 7956 6177
rect 7898 6168 7910 6171
rect 7800 6140 7910 6168
rect 7800 6128 7806 6140
rect 7898 6137 7910 6140
rect 7944 6137 7956 6171
rect 7898 6131 7956 6137
rect 9122 6128 9128 6180
rect 9180 6168 9186 6180
rect 9677 6171 9735 6177
rect 9677 6168 9689 6171
rect 9180 6140 9689 6168
rect 9180 6128 9186 6140
rect 9677 6137 9689 6140
rect 9723 6137 9735 6171
rect 9677 6131 9735 6137
rect 10689 6171 10747 6177
rect 10689 6137 10701 6171
rect 10735 6168 10747 6171
rect 10735 6140 11376 6168
rect 10735 6137 10747 6140
rect 10689 6131 10747 6137
rect 9766 6100 9772 6112
rect 9727 6072 9772 6100
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10778 6100 10784 6112
rect 10739 6072 10784 6100
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 11348 6109 11376 6140
rect 11333 6103 11391 6109
rect 11333 6069 11345 6103
rect 11379 6069 11391 6103
rect 11440 6100 11468 6208
rect 11701 6205 11713 6239
rect 11747 6236 11759 6239
rect 12158 6236 12164 6248
rect 11747 6208 12164 6236
rect 11747 6205 11759 6208
rect 11701 6199 11759 6205
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 15654 6236 15660 6248
rect 12728 6208 15660 6236
rect 11793 6171 11851 6177
rect 11793 6137 11805 6171
rect 11839 6168 11851 6171
rect 12728 6168 12756 6208
rect 15654 6196 15660 6208
rect 15712 6196 15718 6248
rect 15746 6196 15752 6248
rect 15804 6236 15810 6248
rect 16022 6236 16028 6248
rect 15804 6208 16028 6236
rect 15804 6196 15810 6208
rect 16022 6196 16028 6208
rect 16080 6196 16086 6248
rect 16298 6196 16304 6248
rect 16356 6236 16362 6248
rect 16669 6239 16727 6245
rect 16669 6236 16681 6239
rect 16356 6208 16681 6236
rect 16356 6196 16362 6208
rect 16669 6205 16681 6208
rect 16715 6205 16727 6239
rect 16669 6199 16727 6205
rect 11839 6140 12756 6168
rect 12805 6171 12863 6177
rect 11839 6137 11851 6140
rect 11793 6131 11851 6137
rect 12805 6137 12817 6171
rect 12851 6168 12863 6171
rect 12851 6140 13492 6168
rect 12851 6137 12863 6140
rect 12805 6131 12863 6137
rect 12342 6100 12348 6112
rect 11440 6072 12348 6100
rect 11333 6063 11391 6069
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12894 6100 12900 6112
rect 12492 6072 12537 6100
rect 12855 6072 12900 6100
rect 12492 6060 12498 6072
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13464 6109 13492 6140
rect 13538 6128 13544 6180
rect 13596 6168 13602 6180
rect 13909 6171 13967 6177
rect 13909 6168 13921 6171
rect 13596 6140 13921 6168
rect 13596 6128 13602 6140
rect 13909 6137 13921 6140
rect 13955 6168 13967 6171
rect 15286 6168 15292 6180
rect 13955 6140 15292 6168
rect 13955 6137 13967 6140
rect 13909 6131 13967 6137
rect 15286 6128 15292 6140
rect 15344 6128 15350 6180
rect 16390 6168 16396 6180
rect 15672 6140 16396 6168
rect 13449 6103 13507 6109
rect 13449 6069 13461 6103
rect 13495 6069 13507 6103
rect 13449 6063 13507 6069
rect 13817 6103 13875 6109
rect 13817 6069 13829 6103
rect 13863 6100 13875 6103
rect 13998 6100 14004 6112
rect 13863 6072 14004 6100
rect 13863 6069 13875 6072
rect 13817 6063 13875 6069
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 15672 6109 15700 6140
rect 16390 6128 16396 6140
rect 16448 6128 16454 6180
rect 16951 6168 16979 6344
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 18598 6304 18604 6316
rect 18559 6276 18604 6304
rect 18598 6264 18604 6276
rect 18656 6264 18662 6316
rect 19702 6304 19708 6316
rect 19663 6276 19708 6304
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 19889 6307 19947 6313
rect 19889 6273 19901 6307
rect 19935 6304 19947 6307
rect 20162 6304 20168 6316
rect 19935 6276 20168 6304
rect 19935 6273 19947 6276
rect 19889 6267 19947 6273
rect 20162 6264 20168 6276
rect 20220 6264 20226 6316
rect 20346 6264 20352 6316
rect 20404 6304 20410 6316
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 20404 6276 20821 6304
rect 20404 6264 20410 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 18414 6236 18420 6248
rect 18375 6208 18420 6236
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 19058 6196 19064 6248
rect 19116 6236 19122 6248
rect 20625 6239 20683 6245
rect 20625 6236 20637 6239
rect 19116 6208 20637 6236
rect 19116 6196 19122 6208
rect 20625 6205 20637 6208
rect 20671 6205 20683 6239
rect 20625 6199 20683 6205
rect 18509 6171 18567 6177
rect 18509 6168 18521 6171
rect 16951 6140 18521 6168
rect 18509 6137 18521 6140
rect 18555 6137 18567 6171
rect 18509 6131 18567 6137
rect 18966 6128 18972 6180
rect 19024 6168 19030 6180
rect 20717 6171 20775 6177
rect 20717 6168 20729 6171
rect 19024 6140 20729 6168
rect 19024 6128 19030 6140
rect 20717 6137 20729 6140
rect 20763 6137 20775 6171
rect 20717 6131 20775 6137
rect 15657 6103 15715 6109
rect 15657 6069 15669 6103
rect 15703 6069 15715 6103
rect 15657 6063 15715 6069
rect 15746 6060 15752 6112
rect 15804 6100 15810 6112
rect 16298 6100 16304 6112
rect 15804 6072 15849 6100
rect 16259 6072 16304 6100
rect 15804 6060 15810 6072
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 16666 6060 16672 6112
rect 16724 6100 16730 6112
rect 16761 6103 16819 6109
rect 16761 6100 16773 6103
rect 16724 6072 16773 6100
rect 16724 6060 16730 6072
rect 16761 6069 16773 6072
rect 16807 6069 16819 6103
rect 16761 6063 16819 6069
rect 18598 6060 18604 6112
rect 18656 6100 18662 6112
rect 19245 6103 19303 6109
rect 19245 6100 19257 6103
rect 18656 6072 19257 6100
rect 18656 6060 18662 6072
rect 19245 6069 19257 6072
rect 19291 6069 19303 6103
rect 19610 6100 19616 6112
rect 19571 6072 19616 6100
rect 19245 6063 19303 6069
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 20254 6100 20260 6112
rect 20215 6072 20260 6100
rect 20254 6060 20260 6072
rect 20312 6060 20318 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 7800 5868 7849 5896
rect 7800 5856 7806 5868
rect 7837 5865 7849 5868
rect 7883 5865 7895 5899
rect 9122 5896 9128 5908
rect 9083 5868 9128 5896
rect 7837 5859 7895 5865
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 6702 5831 6760 5837
rect 6702 5828 6714 5831
rect 4120 5800 6714 5828
rect 4120 5788 4126 5800
rect 6702 5797 6714 5800
rect 6748 5797 6760 5831
rect 7852 5828 7880 5859
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 9677 5899 9735 5905
rect 9677 5865 9689 5899
rect 9723 5896 9735 5899
rect 9766 5896 9772 5908
rect 9723 5868 9772 5896
rect 9723 5865 9735 5868
rect 9677 5859 9735 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 12989 5899 13047 5905
rect 12989 5896 13001 5899
rect 12492 5868 13001 5896
rect 12492 5856 12498 5868
rect 12989 5865 13001 5868
rect 13035 5865 13047 5899
rect 12989 5859 13047 5865
rect 13170 5856 13176 5908
rect 13228 5896 13234 5908
rect 15746 5896 15752 5908
rect 13228 5868 15752 5896
rect 13228 5856 13234 5868
rect 15746 5856 15752 5868
rect 15804 5896 15810 5908
rect 16022 5896 16028 5908
rect 15804 5868 16028 5896
rect 15804 5856 15810 5868
rect 16022 5856 16028 5868
rect 16080 5856 16086 5908
rect 16482 5856 16488 5908
rect 16540 5896 16546 5908
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 16540 5868 16681 5896
rect 16540 5856 16546 5868
rect 16669 5865 16681 5868
rect 16715 5865 16727 5899
rect 18046 5896 18052 5908
rect 16669 5859 16727 5865
rect 16776 5868 18052 5896
rect 11140 5831 11198 5837
rect 7852 5800 10364 5828
rect 6702 5791 6760 5797
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5760 6515 5763
rect 7650 5760 7656 5772
rect 6503 5732 7656 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 10042 5760 10048 5772
rect 10003 5732 10048 5760
rect 10042 5720 10048 5732
rect 10100 5760 10106 5772
rect 10226 5760 10232 5772
rect 10100 5732 10232 5760
rect 10100 5720 10106 5732
rect 10226 5720 10232 5732
rect 10284 5720 10290 5772
rect 10336 5760 10364 5800
rect 11140 5797 11152 5831
rect 11186 5828 11198 5831
rect 14090 5828 14096 5840
rect 11186 5800 14096 5828
rect 11186 5797 11198 5800
rect 11140 5791 11198 5797
rect 14090 5788 14096 5800
rect 14148 5788 14154 5840
rect 15470 5788 15476 5840
rect 15528 5837 15534 5840
rect 15528 5831 15592 5837
rect 15528 5797 15546 5831
rect 15580 5797 15592 5831
rect 15528 5791 15592 5797
rect 15528 5788 15534 5791
rect 15930 5788 15936 5840
rect 15988 5828 15994 5840
rect 16776 5828 16804 5868
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 18509 5899 18567 5905
rect 18509 5865 18521 5899
rect 18555 5865 18567 5899
rect 18509 5859 18567 5865
rect 15988 5800 16804 5828
rect 15988 5788 15994 5800
rect 17310 5788 17316 5840
rect 17368 5837 17374 5840
rect 17368 5831 17432 5837
rect 17368 5797 17386 5831
rect 17420 5797 17432 5831
rect 18524 5828 18552 5859
rect 19610 5856 19616 5908
rect 19668 5896 19674 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 19668 5868 20913 5896
rect 19668 5856 19674 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 19052 5831 19110 5837
rect 19052 5828 19064 5831
rect 18524 5800 19064 5828
rect 17368 5791 17432 5797
rect 19052 5797 19064 5800
rect 19098 5828 19110 5831
rect 20346 5828 20352 5840
rect 19098 5800 20352 5828
rect 19098 5797 19110 5800
rect 19052 5791 19110 5797
rect 17368 5788 17374 5791
rect 20346 5788 20352 5800
rect 20404 5788 20410 5840
rect 10962 5760 10968 5772
rect 10336 5732 10968 5760
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10336 5701 10364 5732
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12897 5763 12955 5769
rect 12897 5760 12909 5763
rect 12492 5732 12909 5760
rect 12492 5720 12498 5732
rect 12897 5729 12909 5732
rect 12943 5729 12955 5763
rect 13906 5760 13912 5772
rect 13867 5732 13912 5760
rect 12897 5723 12955 5729
rect 13906 5720 13912 5732
rect 13964 5720 13970 5772
rect 14001 5763 14059 5769
rect 14001 5729 14013 5763
rect 14047 5760 14059 5763
rect 14550 5760 14556 5772
rect 14047 5732 14556 5760
rect 14047 5729 14059 5732
rect 14001 5723 14059 5729
rect 14550 5720 14556 5732
rect 14608 5720 14614 5772
rect 15194 5720 15200 5772
rect 15252 5760 15258 5772
rect 15289 5763 15347 5769
rect 15289 5760 15301 5763
rect 15252 5732 15301 5760
rect 15252 5720 15258 5732
rect 15289 5729 15301 5732
rect 15335 5760 15347 5763
rect 17129 5763 17187 5769
rect 17129 5760 17141 5763
rect 15335 5732 17141 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 17129 5729 17141 5732
rect 17175 5760 17187 5763
rect 18785 5763 18843 5769
rect 18785 5760 18797 5763
rect 17175 5732 18797 5760
rect 17175 5729 17187 5732
rect 17129 5723 17187 5729
rect 18785 5729 18797 5732
rect 18831 5729 18843 5763
rect 18785 5723 18843 5729
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5661 10379 5695
rect 10870 5692 10876 5704
rect 10831 5664 10876 5692
rect 10321 5655 10379 5661
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 13173 5695 13231 5701
rect 13173 5661 13185 5695
rect 13219 5692 13231 5695
rect 13814 5692 13820 5704
rect 13219 5664 13820 5692
rect 13219 5661 13231 5664
rect 13173 5655 13231 5661
rect 13814 5652 13820 5664
rect 13872 5652 13878 5704
rect 14090 5652 14096 5704
rect 14148 5692 14154 5704
rect 14148 5664 14193 5692
rect 14148 5652 14154 5664
rect 12253 5627 12311 5633
rect 12253 5593 12265 5627
rect 12299 5624 12311 5627
rect 12986 5624 12992 5636
rect 12299 5596 12992 5624
rect 12299 5593 12311 5596
rect 12253 5587 12311 5593
rect 12986 5584 12992 5596
rect 13044 5584 13050 5636
rect 12529 5559 12587 5565
rect 12529 5525 12541 5559
rect 12575 5556 12587 5559
rect 13354 5556 13360 5568
rect 12575 5528 13360 5556
rect 12575 5525 12587 5528
rect 12529 5519 12587 5525
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 13538 5556 13544 5568
rect 13499 5528 13544 5556
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 18800 5556 18828 5723
rect 19058 5556 19064 5568
rect 18800 5528 19064 5556
rect 19058 5516 19064 5528
rect 19116 5516 19122 5568
rect 20162 5556 20168 5568
rect 20123 5528 20168 5556
rect 20162 5516 20168 5528
rect 20220 5516 20226 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 10321 5355 10379 5361
rect 10321 5321 10333 5355
rect 10367 5352 10379 5355
rect 10778 5352 10784 5364
rect 10367 5324 10784 5352
rect 10367 5321 10379 5324
rect 10321 5315 10379 5321
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 12618 5352 12624 5364
rect 12452 5324 12624 5352
rect 10870 5244 10876 5296
rect 10928 5284 10934 5296
rect 12452 5284 12480 5324
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 13814 5352 13820 5364
rect 13775 5324 13820 5352
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 14001 5355 14059 5361
rect 14001 5321 14013 5355
rect 14047 5352 14059 5355
rect 15194 5352 15200 5364
rect 14047 5324 15200 5352
rect 14047 5321 14059 5324
rect 14001 5315 14059 5321
rect 15194 5312 15200 5324
rect 15252 5312 15258 5364
rect 19426 5352 19432 5364
rect 19260 5324 19432 5352
rect 10928 5256 12480 5284
rect 10928 5244 10934 5256
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 10781 5219 10839 5225
rect 10781 5216 10793 5219
rect 10652 5188 10793 5216
rect 10652 5176 10658 5188
rect 10781 5185 10793 5188
rect 10827 5185 10839 5219
rect 10962 5216 10968 5228
rect 10923 5188 10968 5216
rect 10781 5179 10839 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 12452 5225 12480 5256
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5185 12495 5219
rect 13832 5216 13860 5312
rect 15212 5216 15240 5312
rect 15562 5216 15568 5228
rect 13832 5188 14228 5216
rect 15212 5188 15568 5216
rect 12437 5179 12495 5185
rect 12704 5151 12762 5157
rect 12704 5117 12716 5151
rect 12750 5148 12762 5151
rect 12986 5148 12992 5160
rect 12750 5120 12992 5148
rect 12750 5117 12762 5120
rect 12704 5111 12762 5117
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5148 14059 5151
rect 14093 5151 14151 5157
rect 14093 5148 14105 5151
rect 14047 5120 14105 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 14093 5117 14105 5120
rect 14139 5117 14151 5151
rect 14200 5148 14228 5188
rect 15562 5176 15568 5188
rect 15620 5216 15626 5228
rect 15933 5219 15991 5225
rect 15933 5216 15945 5219
rect 15620 5188 15945 5216
rect 15620 5176 15626 5188
rect 15933 5185 15945 5188
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 18877 5219 18935 5225
rect 18877 5185 18889 5219
rect 18923 5216 18935 5219
rect 19260 5216 19288 5324
rect 19426 5312 19432 5324
rect 19484 5352 19490 5364
rect 20625 5355 20683 5361
rect 20625 5352 20637 5355
rect 19484 5324 20637 5352
rect 19484 5312 19490 5324
rect 20625 5321 20637 5324
rect 20671 5321 20683 5355
rect 20625 5315 20683 5321
rect 18923 5188 19288 5216
rect 18923 5185 18935 5188
rect 18877 5179 18935 5185
rect 14349 5151 14407 5157
rect 14349 5148 14361 5151
rect 14200 5120 14361 5148
rect 14093 5111 14151 5117
rect 14349 5117 14361 5120
rect 14395 5117 14407 5151
rect 14349 5111 14407 5117
rect 14918 5108 14924 5160
rect 14976 5148 14982 5160
rect 16200 5151 16258 5157
rect 14976 5120 15884 5148
rect 14976 5108 14982 5120
rect 10689 5083 10747 5089
rect 10689 5049 10701 5083
rect 10735 5080 10747 5083
rect 15746 5080 15752 5092
rect 10735 5052 15752 5080
rect 10735 5049 10747 5052
rect 10689 5043 10747 5049
rect 15746 5040 15752 5052
rect 15804 5040 15810 5092
rect 15856 5080 15884 5120
rect 16200 5117 16212 5151
rect 16246 5148 16258 5151
rect 16482 5148 16488 5160
rect 16246 5120 16488 5148
rect 16246 5117 16258 5120
rect 16200 5111 16258 5117
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 18598 5148 18604 5160
rect 18559 5120 18604 5148
rect 18598 5108 18604 5120
rect 18656 5108 18662 5160
rect 19058 5108 19064 5160
rect 19116 5148 19122 5160
rect 19245 5151 19303 5157
rect 19245 5148 19257 5151
rect 19116 5120 19257 5148
rect 19116 5108 19122 5120
rect 19245 5117 19257 5120
rect 19291 5117 19303 5151
rect 19245 5111 19303 5117
rect 18046 5080 18052 5092
rect 15856 5052 18052 5080
rect 18046 5040 18052 5052
rect 18104 5040 18110 5092
rect 19512 5083 19570 5089
rect 19512 5049 19524 5083
rect 19558 5080 19570 5083
rect 20162 5080 20168 5092
rect 19558 5052 20168 5080
rect 19558 5049 19570 5052
rect 19512 5043 19570 5049
rect 20162 5040 20168 5052
rect 20220 5040 20226 5092
rect 11885 5015 11943 5021
rect 11885 4981 11897 5015
rect 11931 5012 11943 5015
rect 12342 5012 12348 5024
rect 11931 4984 12348 5012
rect 11931 4981 11943 4984
rect 11885 4975 11943 4981
rect 12342 4972 12348 4984
rect 12400 4972 12406 5024
rect 15470 5012 15476 5024
rect 15431 4984 15476 5012
rect 15470 4972 15476 4984
rect 15528 4972 15534 5024
rect 17310 5012 17316 5024
rect 17271 4984 17316 5012
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 18233 5015 18291 5021
rect 18233 4981 18245 5015
rect 18279 5012 18291 5015
rect 18598 5012 18604 5024
rect 18279 4984 18604 5012
rect 18279 4981 18291 4984
rect 18233 4975 18291 4981
rect 18598 4972 18604 4984
rect 18656 4972 18662 5024
rect 18693 5015 18751 5021
rect 18693 4981 18705 5015
rect 18739 5012 18751 5015
rect 19610 5012 19616 5024
rect 18739 4984 19616 5012
rect 18739 4981 18751 4984
rect 18693 4975 18751 4981
rect 19610 4972 19616 4984
rect 19668 4972 19674 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 12897 4811 12955 4817
rect 12492 4780 12537 4808
rect 12492 4768 12498 4780
rect 12897 4777 12909 4811
rect 12943 4808 12955 4811
rect 13538 4808 13544 4820
rect 12943 4780 13544 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 16025 4811 16083 4817
rect 16025 4777 16037 4811
rect 16071 4808 16083 4811
rect 16298 4808 16304 4820
rect 16071 4780 16304 4808
rect 16071 4777 16083 4780
rect 16025 4771 16083 4777
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 18049 4811 18107 4817
rect 18049 4777 18061 4811
rect 18095 4808 18107 4811
rect 18782 4808 18788 4820
rect 18095 4780 18788 4808
rect 18095 4777 18107 4780
rect 18049 4771 18107 4777
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 19610 4808 19616 4820
rect 19571 4780 19616 4808
rect 19610 4768 19616 4780
rect 19668 4768 19674 4820
rect 19981 4811 20039 4817
rect 19981 4777 19993 4811
rect 20027 4808 20039 4811
rect 20254 4808 20260 4820
rect 20027 4780 20260 4808
rect 20027 4777 20039 4780
rect 19981 4771 20039 4777
rect 20254 4768 20260 4780
rect 20312 4768 20318 4820
rect 9950 4700 9956 4752
rect 10008 4740 10014 4752
rect 16114 4740 16120 4752
rect 10008 4712 13952 4740
rect 16075 4712 16120 4740
rect 10008 4700 10014 4712
rect 12342 4632 12348 4684
rect 12400 4672 12406 4684
rect 13924 4681 13952 4712
rect 16114 4700 16120 4712
rect 16172 4700 16178 4752
rect 12805 4675 12863 4681
rect 12805 4672 12817 4675
rect 12400 4644 12817 4672
rect 12400 4632 12406 4644
rect 12805 4641 12817 4644
rect 12851 4641 12863 4675
rect 12805 4635 12863 4641
rect 13817 4675 13875 4681
rect 13817 4641 13829 4675
rect 13863 4641 13875 4675
rect 13817 4635 13875 4641
rect 13909 4675 13967 4681
rect 13909 4641 13921 4675
rect 13955 4672 13967 4675
rect 14366 4672 14372 4684
rect 13955 4644 14372 4672
rect 13955 4641 13967 4644
rect 13909 4635 13967 4641
rect 12986 4604 12992 4616
rect 12947 4576 12992 4604
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 12894 4496 12900 4548
rect 12952 4536 12958 4548
rect 13449 4539 13507 4545
rect 13449 4536 13461 4539
rect 12952 4508 13461 4536
rect 12952 4496 12958 4508
rect 13449 4505 13461 4508
rect 13495 4505 13507 4539
rect 13832 4536 13860 4635
rect 14366 4632 14372 4644
rect 14424 4632 14430 4684
rect 14461 4675 14519 4681
rect 14461 4641 14473 4675
rect 14507 4672 14519 4675
rect 15102 4672 15108 4684
rect 14507 4644 15108 4672
rect 14507 4641 14519 4644
rect 14461 4635 14519 4641
rect 15102 4632 15108 4644
rect 15160 4632 15166 4684
rect 18417 4675 18475 4681
rect 18417 4641 18429 4675
rect 18463 4672 18475 4675
rect 19061 4675 19119 4681
rect 19061 4672 19073 4675
rect 18463 4644 19073 4672
rect 18463 4641 18475 4644
rect 18417 4635 18475 4641
rect 19061 4641 19073 4644
rect 19107 4641 19119 4675
rect 19061 4635 19119 4641
rect 14090 4604 14096 4616
rect 14051 4576 14096 4604
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 16301 4607 16359 4613
rect 16301 4573 16313 4607
rect 16347 4604 16359 4607
rect 17310 4604 17316 4616
rect 16347 4576 17316 4604
rect 16347 4573 16359 4576
rect 16301 4567 16359 4573
rect 17310 4564 17316 4576
rect 17368 4564 17374 4616
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 18690 4604 18696 4616
rect 18651 4576 18696 4604
rect 18690 4564 18696 4576
rect 18748 4564 18754 4616
rect 20070 4604 20076 4616
rect 20031 4576 20076 4604
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20162 4564 20168 4616
rect 20220 4604 20226 4616
rect 20220 4576 20265 4604
rect 20220 4564 20226 4576
rect 16850 4536 16856 4548
rect 13832 4508 16856 4536
rect 13449 4499 13507 4505
rect 16850 4496 16856 4508
rect 16908 4536 16914 4548
rect 19978 4536 19984 4548
rect 16908 4508 19984 4536
rect 16908 4496 16914 4508
rect 19978 4496 19984 4508
rect 20036 4496 20042 4548
rect 11882 4428 11888 4480
rect 11940 4468 11946 4480
rect 14182 4468 14188 4480
rect 11940 4440 14188 4468
rect 11940 4428 11946 4440
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 14458 4428 14464 4480
rect 14516 4468 14522 4480
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 14516 4440 14657 4468
rect 14516 4428 14522 4440
rect 14645 4437 14657 4440
rect 14691 4437 14703 4471
rect 14645 4431 14703 4437
rect 15657 4471 15715 4477
rect 15657 4437 15669 4471
rect 15703 4468 15715 4471
rect 16298 4468 16304 4480
rect 15703 4440 16304 4468
rect 15703 4437 15715 4440
rect 15657 4431 15715 4437
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 11146 4264 11152 4276
rect 8956 4236 11152 4264
rect 3050 4088 3056 4140
rect 3108 4128 3114 4140
rect 8956 4128 8984 4236
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 12268 4236 13032 4264
rect 3108 4100 8984 4128
rect 3108 4088 3114 4100
rect 9950 4088 9956 4140
rect 10008 4128 10014 4140
rect 12268 4128 12296 4236
rect 12342 4156 12348 4208
rect 12400 4196 12406 4208
rect 12802 4196 12808 4208
rect 12400 4168 12808 4196
rect 12400 4156 12406 4168
rect 12802 4156 12808 4168
rect 12860 4156 12866 4208
rect 10008 4100 12296 4128
rect 13004 4128 13032 4236
rect 18690 4224 18696 4276
rect 18748 4264 18754 4276
rect 19429 4267 19487 4273
rect 19429 4264 19441 4267
rect 18748 4236 19441 4264
rect 18748 4224 18754 4236
rect 19429 4233 19441 4236
rect 19475 4233 19487 4267
rect 19429 4227 19487 4233
rect 19705 4267 19763 4273
rect 19705 4233 19717 4267
rect 19751 4264 19763 4267
rect 20070 4264 20076 4276
rect 19751 4236 20076 4264
rect 19751 4233 19763 4236
rect 19705 4227 19763 4233
rect 20070 4224 20076 4236
rect 20128 4224 20134 4276
rect 15470 4156 15476 4208
rect 15528 4196 15534 4208
rect 17954 4196 17960 4208
rect 15528 4168 15884 4196
rect 15528 4156 15534 4168
rect 13906 4128 13912 4140
rect 13004 4100 13912 4128
rect 10008 4088 10014 4100
rect 13906 4088 13912 4100
rect 13964 4088 13970 4140
rect 14550 4128 14556 4140
rect 14511 4100 14556 4128
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 15856 4137 15884 4168
rect 16132 4168 17960 4196
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4097 15899 4131
rect 15841 4091 15899 4097
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 8754 4060 8760 4072
rect 5868 4032 8760 4060
rect 5868 4020 5874 4032
rect 8754 4020 8760 4032
rect 8812 4020 8818 4072
rect 8938 4060 8944 4072
rect 8899 4032 8944 4060
rect 8938 4020 8944 4032
rect 8996 4020 9002 4072
rect 9214 4069 9220 4072
rect 9208 4023 9220 4069
rect 9272 4060 9278 4072
rect 9272 4032 9308 4060
rect 9214 4020 9220 4023
rect 9272 4020 9278 4032
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 10502 4060 10508 4072
rect 9732 4032 10508 4060
rect 9732 4020 9738 4032
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 11790 4069 11796 4072
rect 11781 4063 11796 4069
rect 11781 4029 11793 4063
rect 11781 4023 11796 4029
rect 11790 4020 11796 4023
rect 11848 4020 11854 4072
rect 12710 4060 12716 4072
rect 12671 4032 12716 4060
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 12986 4060 12992 4072
rect 12947 4032 12992 4060
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 15746 4060 15752 4072
rect 15659 4032 15752 4060
rect 15746 4020 15752 4032
rect 15804 4060 15810 4072
rect 16132 4060 16160 4168
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 20346 4196 20352 4208
rect 20272 4168 20352 4196
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 17862 4128 17868 4140
rect 17276 4100 17868 4128
rect 17276 4088 17282 4100
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 20272 4137 20300 4168
rect 20346 4156 20352 4168
rect 20404 4156 20410 4208
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 16298 4060 16304 4072
rect 15804 4032 16160 4060
rect 16259 4032 16304 4060
rect 15804 4020 15810 4032
rect 16298 4020 16304 4032
rect 16356 4020 16362 4072
rect 17402 4060 17408 4072
rect 17363 4032 17408 4060
rect 17402 4020 17408 4032
rect 17460 4020 17466 4072
rect 18046 4060 18052 4072
rect 18007 4032 18052 4060
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 20165 4063 20223 4069
rect 20165 4060 20177 4063
rect 18156 4032 20177 4060
rect 7466 3952 7472 4004
rect 7524 3992 7530 4004
rect 10042 3992 10048 4004
rect 7524 3964 10048 3992
rect 7524 3952 7530 3964
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 13449 3995 13507 4001
rect 13449 3961 13461 3995
rect 13495 3992 13507 3995
rect 14277 3995 14335 4001
rect 14277 3992 14289 3995
rect 13495 3964 14289 3992
rect 13495 3961 13507 3964
rect 13449 3955 13507 3961
rect 14277 3961 14289 3964
rect 14323 3961 14335 3995
rect 15654 3992 15660 4004
rect 15615 3964 15660 3992
rect 14277 3955 14335 3961
rect 15654 3952 15660 3964
rect 15712 3952 15718 4004
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 16577 3995 16635 4001
rect 16577 3992 16589 3995
rect 15988 3964 16589 3992
rect 15988 3952 15994 3964
rect 16577 3961 16589 3964
rect 16623 3961 16635 3995
rect 16577 3955 16635 3961
rect 17494 3952 17500 4004
rect 17552 3992 17558 4004
rect 18156 3992 18184 4032
rect 20165 4029 20177 4032
rect 20211 4029 20223 4063
rect 20714 4060 20720 4072
rect 20675 4032 20720 4060
rect 20165 4023 20223 4029
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 17552 3964 18184 3992
rect 18316 3995 18374 4001
rect 17552 3952 17558 3964
rect 18316 3961 18328 3995
rect 18362 3992 18374 3995
rect 18598 3992 18604 4004
rect 18362 3964 18604 3992
rect 18362 3961 18374 3964
rect 18316 3955 18374 3961
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 10134 3924 10140 3936
rect 2004 3896 10140 3924
rect 2004 3884 2010 3896
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10318 3924 10324 3936
rect 10279 3896 10324 3924
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 10965 3927 11023 3933
rect 10965 3893 10977 3927
rect 11011 3924 11023 3927
rect 11054 3924 11060 3936
rect 11011 3896 11060 3924
rect 11011 3893 11023 3896
rect 10965 3887 11023 3893
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11977 3927 12035 3933
rect 11977 3893 11989 3927
rect 12023 3924 12035 3927
rect 12526 3924 12532 3936
rect 12023 3896 12532 3924
rect 12023 3893 12035 3896
rect 11977 3887 12035 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 13906 3924 13912 3936
rect 13867 3896 13912 3924
rect 13906 3884 13912 3896
rect 13964 3884 13970 3936
rect 13998 3884 14004 3936
rect 14056 3924 14062 3936
rect 14369 3927 14427 3933
rect 14369 3924 14381 3927
rect 14056 3896 14381 3924
rect 14056 3884 14062 3896
rect 14369 3893 14381 3896
rect 14415 3893 14427 3927
rect 14369 3887 14427 3893
rect 15289 3927 15347 3933
rect 15289 3893 15301 3927
rect 15335 3924 15347 3927
rect 15378 3924 15384 3936
rect 15335 3896 15384 3924
rect 15335 3893 15347 3896
rect 15289 3887 15347 3893
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 17589 3927 17647 3933
rect 17589 3893 17601 3927
rect 17635 3924 17647 3927
rect 17954 3924 17960 3936
rect 17635 3896 17960 3924
rect 17635 3893 17647 3896
rect 17589 3887 17647 3893
rect 17954 3884 17960 3896
rect 18012 3884 18018 3936
rect 20070 3924 20076 3936
rect 20031 3896 20076 3924
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20901 3927 20959 3933
rect 20901 3893 20913 3927
rect 20947 3924 20959 3927
rect 21910 3924 21916 3936
rect 20947 3896 21916 3924
rect 20947 3893 20959 3896
rect 20901 3887 20959 3893
rect 21910 3884 21916 3896
rect 21968 3884 21974 3936
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 12342 3720 12348 3732
rect 4212 3692 12348 3720
rect 4212 3680 4218 3692
rect 12342 3680 12348 3692
rect 12400 3680 12406 3732
rect 12989 3723 13047 3729
rect 12989 3689 13001 3723
rect 13035 3689 13047 3723
rect 12989 3683 13047 3689
rect 290 3612 296 3664
rect 348 3652 354 3664
rect 9950 3652 9956 3664
rect 348 3624 9956 3652
rect 348 3612 354 3624
rect 9950 3612 9956 3624
rect 10008 3612 10014 3664
rect 10220 3655 10278 3661
rect 10220 3621 10232 3655
rect 10266 3652 10278 3655
rect 10318 3652 10324 3664
rect 10266 3624 10324 3652
rect 10266 3621 10278 3624
rect 10220 3615 10278 3621
rect 10318 3612 10324 3624
rect 10376 3652 10382 3664
rect 10870 3652 10876 3664
rect 10376 3624 10876 3652
rect 10376 3612 10382 3624
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 11425 3655 11483 3661
rect 11425 3621 11437 3655
rect 11471 3652 11483 3655
rect 11854 3655 11912 3661
rect 11854 3652 11866 3655
rect 11471 3624 11866 3652
rect 11471 3621 11483 3624
rect 11425 3615 11483 3621
rect 11854 3621 11866 3624
rect 11900 3621 11912 3655
rect 13004 3652 13032 3683
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 14608 3692 14657 3720
rect 14608 3680 14614 3692
rect 14645 3689 14657 3692
rect 14691 3689 14703 3723
rect 15746 3720 15752 3732
rect 14645 3683 14703 3689
rect 15304 3692 15752 3720
rect 13510 3655 13568 3661
rect 13510 3652 13522 3655
rect 13004 3624 13522 3652
rect 11854 3615 11912 3621
rect 13510 3621 13522 3624
rect 13556 3652 13568 3655
rect 13814 3652 13820 3664
rect 13556 3624 13820 3652
rect 13556 3621 13568 3624
rect 13510 3615 13568 3621
rect 13814 3612 13820 3624
rect 13872 3612 13878 3664
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 9674 3584 9680 3596
rect 5316 3556 9680 3584
rect 5316 3544 5322 3556
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 11609 3587 11667 3593
rect 11609 3584 11621 3587
rect 9968 3556 11621 3584
rect 8938 3476 8944 3528
rect 8996 3516 9002 3528
rect 9968 3525 9996 3556
rect 11609 3553 11621 3556
rect 11655 3584 11667 3587
rect 12618 3584 12624 3596
rect 11655 3556 12624 3584
rect 11655 3553 11667 3556
rect 11609 3547 11667 3553
rect 12618 3544 12624 3556
rect 12676 3584 12682 3596
rect 13265 3587 13323 3593
rect 13265 3584 13277 3587
rect 12676 3556 13277 3584
rect 12676 3544 12682 3556
rect 13265 3553 13277 3556
rect 13311 3553 13323 3587
rect 15304 3584 15332 3692
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 16945 3723 17003 3729
rect 16945 3689 16957 3723
rect 16991 3689 17003 3723
rect 18598 3720 18604 3732
rect 18559 3692 18604 3720
rect 16945 3683 17003 3689
rect 15832 3655 15890 3661
rect 15832 3621 15844 3655
rect 15878 3652 15890 3655
rect 16022 3652 16028 3664
rect 15878 3624 16028 3652
rect 15878 3621 15890 3624
rect 15832 3615 15890 3621
rect 16022 3612 16028 3624
rect 16080 3612 16086 3664
rect 16960 3652 16988 3683
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 17126 3652 17132 3664
rect 16960 3624 17132 3652
rect 17126 3612 17132 3624
rect 17184 3652 17190 3664
rect 17466 3655 17524 3661
rect 17466 3652 17478 3655
rect 17184 3624 17478 3652
rect 17184 3612 17190 3624
rect 17466 3621 17478 3624
rect 17512 3621 17524 3655
rect 17466 3615 17524 3621
rect 15562 3584 15568 3596
rect 13265 3547 13323 3553
rect 13372 3556 15332 3584
rect 15523 3556 15568 3584
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 8996 3488 9965 3516
rect 8996 3476 9002 3488
rect 9953 3485 9965 3488
rect 9999 3485 10011 3519
rect 13372 3516 13400 3556
rect 15562 3544 15568 3556
rect 15620 3584 15626 3596
rect 17221 3587 17279 3593
rect 17221 3584 17233 3587
rect 15620 3556 17233 3584
rect 15620 3544 15626 3556
rect 17221 3553 17233 3556
rect 17267 3584 17279 3587
rect 18046 3584 18052 3596
rect 17267 3556 18052 3584
rect 17267 3553 17279 3556
rect 17221 3547 17279 3553
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 18690 3544 18696 3596
rect 18748 3584 18754 3596
rect 19061 3587 19119 3593
rect 19061 3584 19073 3587
rect 18748 3556 19073 3584
rect 18748 3544 18754 3556
rect 19061 3553 19073 3556
rect 19107 3553 19119 3587
rect 19794 3584 19800 3596
rect 19755 3556 19800 3584
rect 19061 3547 19119 3553
rect 19794 3544 19800 3556
rect 19852 3544 19858 3596
rect 9953 3479 10011 3485
rect 12636 3488 13400 3516
rect 19337 3519 19395 3525
rect 12636 3460 12664 3488
rect 19337 3485 19349 3519
rect 19383 3516 19395 3519
rect 19518 3516 19524 3528
rect 19383 3488 19524 3516
rect 19383 3485 19395 3488
rect 19337 3479 19395 3485
rect 19518 3476 19524 3488
rect 19576 3476 19582 3528
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3516 20131 3519
rect 20346 3516 20352 3528
rect 20119 3488 20352 3516
rect 20119 3485 20131 3488
rect 20073 3479 20131 3485
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 11333 3451 11391 3457
rect 11333 3448 11345 3451
rect 11204 3420 11345 3448
rect 11204 3408 11210 3420
rect 11333 3417 11345 3420
rect 11379 3448 11391 3451
rect 11425 3451 11483 3457
rect 11425 3448 11437 3451
rect 11379 3420 11437 3448
rect 11379 3417 11391 3420
rect 11333 3411 11391 3417
rect 11425 3417 11437 3420
rect 11471 3417 11483 3451
rect 11425 3411 11483 3417
rect 12618 3408 12624 3460
rect 12676 3408 12682 3460
rect 3602 3340 3608 3392
rect 3660 3380 3666 3392
rect 13446 3380 13452 3392
rect 3660 3352 13452 3380
rect 3660 3340 3666 3352
rect 13446 3340 13452 3352
rect 13504 3340 13510 3392
rect 13906 3340 13912 3392
rect 13964 3380 13970 3392
rect 19702 3380 19708 3392
rect 13964 3352 19708 3380
rect 13964 3340 13970 3352
rect 19702 3340 19708 3352
rect 19760 3340 19766 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 10321 3179 10379 3185
rect 10321 3145 10333 3179
rect 10367 3176 10379 3179
rect 10505 3179 10563 3185
rect 10505 3176 10517 3179
rect 10367 3148 10517 3176
rect 10367 3145 10379 3148
rect 10321 3139 10379 3145
rect 10505 3145 10517 3148
rect 10551 3145 10563 3179
rect 10686 3176 10692 3188
rect 10647 3148 10692 3176
rect 10505 3139 10563 3145
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 10778 3136 10784 3188
rect 10836 3176 10842 3188
rect 12434 3176 12440 3188
rect 10836 3148 12440 3176
rect 10836 3136 10842 3148
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 13265 3179 13323 3185
rect 13265 3145 13277 3179
rect 13311 3176 13323 3179
rect 13998 3176 14004 3188
rect 13311 3148 14004 3176
rect 13311 3145 13323 3148
rect 13265 3139 13323 3145
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 16485 3179 16543 3185
rect 14240 3148 16160 3176
rect 14240 3136 14246 3148
rect 6549 3111 6607 3117
rect 6549 3077 6561 3111
rect 6595 3108 6607 3111
rect 8294 3108 8300 3120
rect 6595 3080 8300 3108
rect 6595 3077 6607 3080
rect 6549 3071 6607 3077
rect 8294 3068 8300 3080
rect 8352 3068 8358 3120
rect 10042 3068 10048 3120
rect 10100 3108 10106 3120
rect 15657 3111 15715 3117
rect 10100 3080 13676 3108
rect 10100 3068 10106 3080
rect 8570 3000 8576 3052
rect 8628 3040 8634 3052
rect 10505 3043 10563 3049
rect 8628 3012 10272 3040
rect 8628 3000 8634 3012
rect 10137 2975 10195 2981
rect 10137 2941 10149 2975
rect 10183 2941 10195 2975
rect 10244 2972 10272 3012
rect 10505 3009 10517 3043
rect 10551 3040 10563 3043
rect 10551 3012 11284 3040
rect 10551 3009 10563 3012
rect 10505 3003 10563 3009
rect 10778 2972 10784 2984
rect 10244 2944 10784 2972
rect 10137 2935 10195 2941
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 10042 2904 10048 2916
rect 8352 2876 10048 2904
rect 8352 2864 8358 2876
rect 10042 2864 10048 2876
rect 10100 2864 10106 2916
rect 10152 2904 10180 2935
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 11054 2972 11060 2984
rect 11015 2944 11060 2972
rect 11054 2932 11060 2944
rect 11112 2932 11118 2984
rect 11256 2972 11284 3012
rect 11330 3000 11336 3052
rect 11388 3040 11394 3052
rect 11388 3012 11433 3040
rect 11388 3000 11394 3012
rect 11514 2972 11520 2984
rect 11256 2944 11520 2972
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 11793 2975 11851 2981
rect 11793 2941 11805 2975
rect 11839 2972 11851 2975
rect 12342 2972 12348 2984
rect 11839 2944 12348 2972
rect 11839 2941 11851 2944
rect 11793 2935 11851 2941
rect 12342 2932 12348 2944
rect 12400 2932 12406 2984
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 13262 2972 13268 2984
rect 12483 2944 13268 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 13648 2981 13676 3080
rect 15657 3077 15669 3111
rect 15703 3108 15715 3111
rect 16022 3108 16028 3120
rect 15703 3080 16028 3108
rect 15703 3077 15715 3080
rect 15657 3071 15715 3077
rect 16022 3068 16028 3080
rect 16080 3068 16086 3120
rect 16132 3108 16160 3148
rect 16485 3145 16497 3179
rect 16531 3176 16543 3179
rect 17034 3176 17040 3188
rect 16531 3148 17040 3176
rect 16531 3145 16543 3148
rect 16485 3139 16543 3145
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 18049 3179 18107 3185
rect 18049 3145 18061 3179
rect 18095 3176 18107 3179
rect 18506 3176 18512 3188
rect 18095 3148 18512 3176
rect 18095 3145 18107 3148
rect 18049 3139 18107 3145
rect 18506 3136 18512 3148
rect 18564 3136 18570 3188
rect 19521 3111 19579 3117
rect 16132 3080 19472 3108
rect 13906 3040 13912 3052
rect 13867 3012 13912 3040
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 18598 3040 18604 3052
rect 18559 3012 18604 3040
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 19444 3040 19472 3080
rect 19521 3077 19533 3111
rect 19567 3108 19579 3111
rect 20254 3108 20260 3120
rect 19567 3080 20260 3108
rect 19567 3077 19579 3080
rect 19521 3071 19579 3077
rect 20254 3068 20260 3080
rect 20312 3068 20318 3120
rect 20070 3040 20076 3052
rect 19444 3012 20076 3040
rect 20070 3000 20076 3012
rect 20128 3040 20134 3052
rect 20128 3012 20576 3040
rect 20128 3000 20134 3012
rect 14550 2981 14556 2984
rect 13633 2975 13691 2981
rect 13633 2941 13645 2975
rect 13679 2941 13691 2975
rect 13633 2935 13691 2941
rect 14277 2975 14335 2981
rect 14277 2941 14289 2975
rect 14323 2941 14335 2975
rect 14544 2972 14556 2981
rect 14511 2944 14556 2972
rect 14277 2935 14335 2941
rect 14544 2935 14556 2944
rect 12713 2907 12771 2913
rect 12713 2904 12725 2907
rect 10152 2876 12725 2904
rect 12713 2873 12725 2876
rect 12759 2873 12771 2907
rect 14182 2904 14188 2916
rect 12713 2867 12771 2873
rect 13188 2876 14188 2904
rect 2498 2796 2504 2848
rect 2556 2836 2562 2848
rect 6549 2839 6607 2845
rect 6549 2836 6561 2839
rect 2556 2808 6561 2836
rect 2556 2796 2562 2808
rect 6549 2805 6561 2808
rect 6595 2805 6607 2839
rect 6549 2799 6607 2805
rect 9674 2796 9680 2848
rect 9732 2836 9738 2848
rect 10962 2836 10968 2848
rect 9732 2808 10968 2836
rect 9732 2796 9738 2808
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 11146 2796 11152 2848
rect 11204 2836 11210 2848
rect 11204 2808 11249 2836
rect 11204 2796 11210 2808
rect 11514 2796 11520 2848
rect 11572 2836 11578 2848
rect 11790 2836 11796 2848
rect 11572 2808 11796 2836
rect 11572 2796 11578 2808
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 11977 2839 12035 2845
rect 11977 2805 11989 2839
rect 12023 2836 12035 2839
rect 13188 2836 13216 2876
rect 14182 2864 14188 2876
rect 14240 2864 14246 2916
rect 14292 2904 14320 2935
rect 14550 2932 14556 2935
rect 14608 2932 14614 2984
rect 15930 2972 15936 2984
rect 15891 2944 15936 2972
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 17862 2972 17868 2984
rect 16132 2944 17868 2972
rect 15562 2904 15568 2916
rect 14292 2876 15568 2904
rect 15562 2864 15568 2876
rect 15620 2864 15626 2916
rect 16132 2904 16160 2944
rect 17862 2932 17868 2944
rect 17920 2932 17926 2984
rect 18509 2975 18567 2981
rect 18509 2941 18521 2975
rect 18555 2972 18567 2975
rect 18782 2972 18788 2984
rect 18555 2944 18788 2972
rect 18555 2941 18567 2944
rect 18509 2935 18567 2941
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2972 19395 2975
rect 19886 2972 19892 2984
rect 19383 2944 19892 2972
rect 19383 2941 19395 2944
rect 19337 2935 19395 2941
rect 19886 2932 19892 2944
rect 19944 2932 19950 2984
rect 19978 2932 19984 2984
rect 20036 2972 20042 2984
rect 20548 2981 20576 3012
rect 20533 2975 20591 2981
rect 20036 2944 20081 2972
rect 20036 2932 20042 2944
rect 20533 2941 20545 2975
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 15672 2876 16160 2904
rect 16853 2907 16911 2913
rect 12023 2808 13216 2836
rect 13725 2839 13783 2845
rect 12023 2805 12035 2808
rect 11977 2799 12035 2805
rect 13725 2805 13737 2839
rect 13771 2836 13783 2839
rect 15672 2836 15700 2876
rect 16853 2873 16865 2907
rect 16899 2904 16911 2907
rect 17497 2907 17555 2913
rect 17497 2904 17509 2907
rect 16899 2876 17509 2904
rect 16899 2873 16911 2876
rect 16853 2867 16911 2873
rect 17497 2873 17509 2876
rect 17543 2873 17555 2907
rect 18414 2904 18420 2916
rect 18375 2876 18420 2904
rect 17497 2867 17555 2873
rect 18414 2864 18420 2876
rect 18472 2904 18478 2916
rect 18877 2907 18935 2913
rect 18877 2904 18889 2907
rect 18472 2876 18889 2904
rect 18472 2864 18478 2876
rect 18877 2873 18889 2876
rect 18923 2873 18935 2907
rect 21358 2904 21364 2916
rect 18877 2867 18935 2873
rect 20180 2876 21364 2904
rect 13771 2808 15700 2836
rect 16117 2839 16175 2845
rect 13771 2805 13783 2808
rect 13725 2799 13783 2805
rect 16117 2805 16129 2839
rect 16163 2836 16175 2839
rect 16390 2836 16396 2848
rect 16163 2808 16396 2836
rect 16163 2805 16175 2808
rect 16117 2799 16175 2805
rect 16390 2796 16396 2808
rect 16448 2796 16454 2848
rect 16942 2796 16948 2848
rect 17000 2836 17006 2848
rect 20180 2845 20208 2876
rect 21358 2864 21364 2876
rect 21416 2864 21422 2916
rect 20165 2839 20223 2845
rect 17000 2808 17045 2836
rect 17000 2796 17006 2808
rect 20165 2805 20177 2839
rect 20211 2805 20223 2839
rect 20165 2799 20223 2805
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 22462 2836 22468 2848
rect 20763 2808 22468 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 22462 2796 22468 2808
rect 22520 2796 22526 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 10321 2635 10379 2641
rect 10321 2601 10333 2635
rect 10367 2632 10379 2635
rect 11146 2632 11152 2644
rect 10367 2604 11152 2632
rect 10367 2601 10379 2604
rect 10321 2595 10379 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 15841 2635 15899 2641
rect 15841 2632 15853 2635
rect 11348 2604 15853 2632
rect 4706 2456 4712 2508
rect 4764 2496 4770 2508
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 4764 2468 10701 2496
rect 4764 2456 4770 2468
rect 10689 2465 10701 2468
rect 10735 2465 10747 2499
rect 10689 2459 10747 2465
rect 10781 2499 10839 2505
rect 10781 2465 10793 2499
rect 10827 2496 10839 2499
rect 10962 2496 10968 2508
rect 10827 2468 10968 2496
rect 10827 2465 10839 2468
rect 10781 2459 10839 2465
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 10870 2428 10876 2440
rect 10831 2400 10876 2428
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 1394 2320 1400 2372
rect 1452 2360 1458 2372
rect 11348 2360 11376 2604
rect 15841 2601 15853 2604
rect 15887 2601 15899 2635
rect 15841 2595 15899 2601
rect 15933 2635 15991 2641
rect 15933 2601 15945 2635
rect 15979 2632 15991 2635
rect 16206 2632 16212 2644
rect 15979 2604 16212 2632
rect 15979 2601 15991 2604
rect 15933 2595 15991 2601
rect 16206 2592 16212 2604
rect 16264 2592 16270 2644
rect 17678 2592 17684 2644
rect 17736 2632 17742 2644
rect 17736 2604 19012 2632
rect 17736 2592 17742 2604
rect 12434 2524 12440 2576
rect 12492 2564 12498 2576
rect 13633 2567 13691 2573
rect 13633 2564 13645 2567
rect 12492 2536 13645 2564
rect 12492 2524 12498 2536
rect 13633 2533 13645 2536
rect 13679 2533 13691 2567
rect 13633 2527 13691 2533
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2465 11483 2499
rect 11425 2459 11483 2465
rect 11977 2499 12035 2505
rect 11977 2465 11989 2499
rect 12023 2496 12035 2499
rect 12066 2496 12072 2508
rect 12023 2468 12072 2496
rect 12023 2465 12035 2468
rect 11977 2459 12035 2465
rect 11440 2428 11468 2459
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 12250 2456 12256 2508
rect 12308 2496 12314 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12308 2468 12633 2496
rect 12308 2456 12314 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 13354 2496 13360 2508
rect 13315 2468 13360 2496
rect 12621 2459 12679 2465
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 14274 2496 14280 2508
rect 14235 2468 14280 2496
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14424 2468 14841 2496
rect 14424 2456 14430 2468
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 14829 2459 14887 2465
rect 16114 2456 16120 2508
rect 16172 2496 16178 2508
rect 16485 2499 16543 2505
rect 16485 2496 16497 2499
rect 16172 2468 16497 2496
rect 16172 2456 16178 2468
rect 16485 2465 16497 2468
rect 16531 2465 16543 2499
rect 16485 2459 16543 2465
rect 17313 2499 17371 2505
rect 17313 2465 17325 2499
rect 17359 2496 17371 2499
rect 17494 2496 17500 2508
rect 17359 2468 17500 2496
rect 17359 2465 17371 2468
rect 17313 2459 17371 2465
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 17770 2456 17776 2508
rect 17828 2496 17834 2508
rect 18984 2505 19012 2604
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 17828 2468 18337 2496
rect 17828 2456 17834 2468
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 18969 2499 19027 2505
rect 18969 2465 18981 2499
rect 19015 2465 19027 2499
rect 19518 2496 19524 2508
rect 19479 2468 19524 2496
rect 18969 2459 19027 2465
rect 19518 2456 19524 2468
rect 19576 2456 19582 2508
rect 20346 2496 20352 2508
rect 20307 2468 20352 2496
rect 20346 2456 20352 2468
rect 20404 2456 20410 2508
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 11440 2400 12817 2428
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 16022 2428 16028 2440
rect 15983 2400 16028 2428
rect 12805 2391 12863 2397
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 16942 2388 16948 2440
rect 17000 2388 17006 2440
rect 1452 2332 11376 2360
rect 11609 2363 11667 2369
rect 1452 2320 1458 2332
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 13078 2360 13084 2372
rect 11655 2332 13084 2360
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 13078 2320 13084 2332
rect 13136 2320 13142 2372
rect 14461 2363 14519 2369
rect 14461 2329 14473 2363
rect 14507 2360 14519 2363
rect 15286 2360 15292 2372
rect 14507 2332 15292 2360
rect 14507 2329 14519 2332
rect 14461 2323 14519 2329
rect 15286 2320 15292 2332
rect 15344 2320 15350 2372
rect 15838 2360 15844 2372
rect 15396 2332 15844 2360
rect 12161 2295 12219 2301
rect 12161 2261 12173 2295
rect 12207 2292 12219 2295
rect 13630 2292 13636 2304
rect 12207 2264 13636 2292
rect 12207 2261 12219 2264
rect 12161 2255 12219 2261
rect 13630 2252 13636 2264
rect 13688 2252 13694 2304
rect 15013 2295 15071 2301
rect 15013 2261 15025 2295
rect 15059 2292 15071 2295
rect 15396 2292 15424 2332
rect 15838 2320 15844 2332
rect 15896 2320 15902 2372
rect 16960 2360 16988 2388
rect 16224 2332 16988 2360
rect 15059 2264 15424 2292
rect 15473 2295 15531 2301
rect 15059 2261 15071 2264
rect 15013 2255 15071 2261
rect 15473 2261 15485 2295
rect 15519 2292 15531 2295
rect 16224 2292 16252 2332
rect 18598 2320 18604 2372
rect 18656 2360 18662 2372
rect 19705 2363 19763 2369
rect 19705 2360 19717 2363
rect 18656 2332 19717 2360
rect 18656 2320 18662 2332
rect 19705 2329 19717 2332
rect 19751 2329 19763 2363
rect 19705 2323 19763 2329
rect 15519 2264 16252 2292
rect 16669 2295 16727 2301
rect 15519 2261 15531 2264
rect 15473 2255 15531 2261
rect 16669 2261 16681 2295
rect 16715 2292 16727 2295
rect 16942 2292 16948 2304
rect 16715 2264 16948 2292
rect 16715 2261 16727 2264
rect 16669 2255 16727 2261
rect 16942 2252 16948 2264
rect 17000 2252 17006 2304
rect 17494 2292 17500 2304
rect 17455 2264 17500 2292
rect 17494 2252 17500 2264
rect 17552 2252 17558 2304
rect 18509 2295 18567 2301
rect 18509 2261 18521 2295
rect 18555 2292 18567 2295
rect 19058 2292 19064 2304
rect 18555 2264 19064 2292
rect 18555 2261 18567 2264
rect 18509 2255 18567 2261
rect 19058 2252 19064 2264
rect 19116 2252 19122 2304
rect 19153 2295 19211 2301
rect 19153 2261 19165 2295
rect 19199 2292 19211 2295
rect 19610 2292 19616 2304
rect 19199 2264 19616 2292
rect 19199 2261 19211 2264
rect 19153 2255 19211 2261
rect 19610 2252 19616 2264
rect 19668 2252 19674 2304
rect 20533 2295 20591 2301
rect 20533 2261 20545 2295
rect 20579 2292 20591 2295
rect 20806 2292 20812 2304
rect 20579 2264 20812 2292
rect 20579 2261 20591 2264
rect 20533 2255 20591 2261
rect 20806 2252 20812 2264
rect 20864 2252 20870 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
<< via1 >>
rect 13268 20680 13320 20732
rect 17960 20680 18012 20732
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 9128 20000 9180 20052
rect 11336 20000 11388 20052
rect 12532 20000 12584 20052
rect 13084 20000 13136 20052
rect 15292 20000 15344 20052
rect 7472 19932 7524 19984
rect 11612 19932 11664 19984
rect 16948 20000 17000 20052
rect 17500 20000 17552 20052
rect 18512 20043 18564 20052
rect 18512 20009 18521 20043
rect 18521 20009 18555 20043
rect 18555 20009 18564 20043
rect 18512 20000 18564 20009
rect 19064 20043 19116 20052
rect 19064 20009 19073 20043
rect 19073 20009 19107 20043
rect 19107 20009 19116 20043
rect 19064 20000 19116 20009
rect 19156 20000 19208 20052
rect 19248 20000 19300 20052
rect 6368 19864 6420 19916
rect 9404 19864 9456 19916
rect 10140 19907 10192 19916
rect 10140 19873 10149 19907
rect 10149 19873 10183 19907
rect 10183 19873 10192 19907
rect 10140 19864 10192 19873
rect 12256 19864 12308 19916
rect 12992 19864 13044 19916
rect 9220 19839 9272 19848
rect 9220 19805 9229 19839
rect 9229 19805 9263 19839
rect 9263 19805 9272 19839
rect 10232 19839 10284 19848
rect 9220 19796 9272 19805
rect 10232 19805 10241 19839
rect 10241 19805 10275 19839
rect 10275 19805 10284 19839
rect 10232 19796 10284 19805
rect 10324 19839 10376 19848
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 10324 19796 10376 19805
rect 12348 19796 12400 19848
rect 14280 19864 14332 19916
rect 15200 19864 15252 19916
rect 16028 19864 16080 19916
rect 16672 19907 16724 19916
rect 16672 19873 16681 19907
rect 16681 19873 16715 19907
rect 16715 19873 16724 19907
rect 16672 19864 16724 19873
rect 16856 19864 16908 19916
rect 18788 19864 18840 19916
rect 19156 19864 19208 19916
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 20536 19907 20588 19916
rect 16488 19796 16540 19848
rect 20536 19873 20545 19907
rect 20545 19873 20579 19907
rect 20579 19873 20588 19907
rect 20536 19864 20588 19873
rect 20904 19796 20956 19848
rect 18604 19728 18656 19780
rect 8668 19703 8720 19712
rect 8668 19669 8677 19703
rect 8677 19669 8711 19703
rect 8711 19669 8720 19703
rect 8668 19660 8720 19669
rect 9772 19703 9824 19712
rect 9772 19669 9781 19703
rect 9781 19669 9815 19703
rect 9815 19669 9824 19703
rect 9772 19660 9824 19669
rect 11888 19660 11940 19712
rect 18512 19660 18564 19712
rect 20260 19660 20312 19712
rect 20628 19660 20680 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 10232 19456 10284 19508
rect 17776 19456 17828 19508
rect 18972 19456 19024 19508
rect 8392 19295 8444 19304
rect 8392 19261 8401 19295
rect 8401 19261 8435 19295
rect 8435 19261 8444 19295
rect 8392 19252 8444 19261
rect 8484 19252 8536 19304
rect 9220 19184 9272 19236
rect 9956 19184 10008 19236
rect 10232 19184 10284 19236
rect 11704 19295 11756 19304
rect 11704 19261 11713 19295
rect 11713 19261 11747 19295
rect 11747 19261 11756 19295
rect 11704 19252 11756 19261
rect 14096 19295 14148 19304
rect 14096 19261 14105 19295
rect 14105 19261 14139 19295
rect 14139 19261 14148 19295
rect 14096 19252 14148 19261
rect 14188 19252 14240 19304
rect 12624 19184 12676 19236
rect 13636 19184 13688 19236
rect 2504 19116 2556 19168
rect 9588 19116 9640 19168
rect 9680 19116 9732 19168
rect 11428 19159 11480 19168
rect 11428 19125 11437 19159
rect 11437 19125 11471 19159
rect 11471 19125 11480 19159
rect 11428 19116 11480 19125
rect 11980 19116 12032 19168
rect 12440 19116 12492 19168
rect 12532 19116 12584 19168
rect 12900 19116 12952 19168
rect 13544 19116 13596 19168
rect 14556 19252 14608 19304
rect 15476 19252 15528 19304
rect 15568 19252 15620 19304
rect 16764 19252 16816 19304
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 15292 19184 15344 19236
rect 19340 19252 19392 19304
rect 19984 19295 20036 19304
rect 19984 19261 19993 19295
rect 19993 19261 20027 19295
rect 20027 19261 20036 19295
rect 19984 19252 20036 19261
rect 20352 19252 20404 19304
rect 18512 19184 18564 19236
rect 21364 19184 21416 19236
rect 15016 19116 15068 19168
rect 15844 19116 15896 19168
rect 16396 19116 16448 19168
rect 18696 19116 18748 19168
rect 19248 19116 19300 19168
rect 20168 19159 20220 19168
rect 20168 19125 20177 19159
rect 20177 19125 20211 19159
rect 20211 19125 20220 19159
rect 20168 19116 20220 19125
rect 20812 19116 20864 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 296 18912 348 18964
rect 7380 18776 7432 18828
rect 8392 18844 8444 18896
rect 8760 18776 8812 18828
rect 1400 18708 1452 18760
rect 4712 18572 4764 18624
rect 6184 18572 6236 18624
rect 9220 18912 9272 18964
rect 10140 18955 10192 18964
rect 10140 18921 10149 18955
rect 10149 18921 10183 18955
rect 10183 18921 10192 18955
rect 10140 18912 10192 18921
rect 12348 18912 12400 18964
rect 13636 18912 13688 18964
rect 15568 18912 15620 18964
rect 20076 18912 20128 18964
rect 9680 18844 9732 18896
rect 10232 18844 10284 18896
rect 10508 18844 10560 18896
rect 11428 18844 11480 18896
rect 12900 18887 12952 18896
rect 12900 18853 12934 18887
rect 12934 18853 12952 18887
rect 12900 18844 12952 18853
rect 19156 18887 19208 18896
rect 19156 18853 19165 18887
rect 19165 18853 19199 18887
rect 19199 18853 19208 18887
rect 19156 18844 19208 18853
rect 19432 18844 19484 18896
rect 9772 18776 9824 18828
rect 10140 18776 10192 18828
rect 10232 18708 10284 18760
rect 12440 18776 12492 18828
rect 14464 18776 14516 18828
rect 15752 18776 15804 18828
rect 16120 18776 16172 18828
rect 18604 18776 18656 18828
rect 18880 18819 18932 18828
rect 18880 18785 18889 18819
rect 18889 18785 18923 18819
rect 18923 18785 18932 18819
rect 18880 18776 18932 18785
rect 19524 18776 19576 18828
rect 9956 18640 10008 18692
rect 15384 18708 15436 18760
rect 17960 18708 18012 18760
rect 18512 18708 18564 18760
rect 11796 18572 11848 18624
rect 14004 18615 14056 18624
rect 14004 18581 14013 18615
rect 14013 18581 14047 18615
rect 14047 18581 14056 18615
rect 14004 18572 14056 18581
rect 19708 18640 19760 18692
rect 17224 18572 17276 18624
rect 19248 18572 19300 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 8208 18368 8260 18420
rect 12900 18368 12952 18420
rect 3056 18300 3108 18352
rect 8668 18232 8720 18284
rect 9680 18232 9732 18284
rect 11980 18300 12032 18352
rect 10324 18232 10376 18284
rect 10508 18275 10560 18284
rect 10508 18241 10517 18275
rect 10517 18241 10551 18275
rect 10551 18241 10560 18275
rect 10508 18232 10560 18241
rect 15292 18368 15344 18420
rect 15752 18368 15804 18420
rect 17868 18368 17920 18420
rect 17960 18368 18012 18420
rect 18144 18300 18196 18352
rect 4160 18164 4212 18216
rect 3608 18096 3660 18148
rect 8576 18096 8628 18148
rect 9588 18028 9640 18080
rect 9772 18028 9824 18080
rect 10140 18164 10192 18216
rect 10692 18164 10744 18216
rect 13728 18207 13780 18216
rect 13728 18173 13737 18207
rect 13737 18173 13771 18207
rect 13771 18173 13780 18207
rect 13728 18164 13780 18173
rect 17224 18232 17276 18284
rect 18972 18232 19024 18284
rect 19156 18232 19208 18284
rect 14004 18207 14056 18216
rect 14004 18173 14038 18207
rect 14038 18173 14056 18207
rect 14004 18164 14056 18173
rect 15384 18207 15436 18216
rect 9956 18028 10008 18080
rect 10048 18028 10100 18080
rect 10784 18028 10836 18080
rect 12072 18028 12124 18080
rect 13912 18096 13964 18148
rect 13084 18071 13136 18080
rect 13084 18037 13093 18071
rect 13093 18037 13127 18071
rect 13127 18037 13136 18071
rect 13084 18028 13136 18037
rect 13176 18071 13228 18080
rect 13176 18037 13185 18071
rect 13185 18037 13219 18071
rect 13219 18037 13228 18071
rect 13176 18028 13228 18037
rect 13728 18028 13780 18080
rect 15384 18173 15393 18207
rect 15393 18173 15427 18207
rect 15427 18173 15436 18207
rect 15384 18164 15436 18173
rect 17408 18207 17460 18216
rect 17408 18173 17417 18207
rect 17417 18173 17451 18207
rect 17451 18173 17460 18207
rect 17408 18164 17460 18173
rect 17776 18164 17828 18216
rect 18052 18164 18104 18216
rect 19800 18207 19852 18216
rect 19800 18173 19809 18207
rect 19809 18173 19843 18207
rect 19843 18173 19852 18207
rect 19800 18164 19852 18173
rect 19892 18164 19944 18216
rect 15936 18096 15988 18148
rect 16304 18096 16356 18148
rect 16120 18028 16172 18080
rect 17960 18096 18012 18148
rect 18696 18028 18748 18080
rect 19064 18028 19116 18080
rect 20720 18071 20772 18080
rect 20720 18037 20729 18071
rect 20729 18037 20763 18071
rect 20763 18037 20772 18071
rect 20720 18028 20772 18037
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 8760 17867 8812 17876
rect 8760 17833 8769 17867
rect 8769 17833 8803 17867
rect 8803 17833 8812 17867
rect 8760 17824 8812 17833
rect 9680 17824 9732 17876
rect 13084 17824 13136 17876
rect 848 17756 900 17808
rect 7380 17731 7432 17740
rect 7380 17697 7389 17731
rect 7389 17697 7423 17731
rect 7423 17697 7432 17731
rect 7380 17688 7432 17697
rect 8392 17688 8444 17740
rect 9956 17688 10008 17740
rect 11060 17688 11112 17740
rect 10876 17663 10928 17672
rect 10876 17629 10885 17663
rect 10885 17629 10919 17663
rect 10919 17629 10928 17663
rect 10876 17620 10928 17629
rect 11152 17484 11204 17536
rect 11520 17731 11572 17740
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 11980 17731 12032 17740
rect 11980 17697 11989 17731
rect 11989 17697 12023 17731
rect 12023 17697 12032 17731
rect 11980 17688 12032 17697
rect 13360 17620 13412 17672
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13912 17688 13964 17740
rect 18052 17824 18104 17876
rect 18420 17824 18472 17876
rect 18604 17867 18656 17876
rect 18604 17833 18613 17867
rect 18613 17833 18647 17867
rect 18647 17833 18656 17867
rect 18604 17824 18656 17833
rect 20536 17756 20588 17808
rect 15384 17688 15436 17740
rect 17224 17731 17276 17740
rect 17224 17697 17258 17731
rect 17258 17697 17276 17731
rect 17224 17688 17276 17697
rect 13544 17620 13596 17629
rect 15568 17620 15620 17672
rect 15660 17620 15712 17672
rect 16120 17663 16172 17672
rect 16120 17629 16129 17663
rect 16129 17629 16163 17663
rect 16163 17629 16172 17663
rect 16120 17620 16172 17629
rect 16948 17663 17000 17672
rect 16948 17629 16957 17663
rect 16957 17629 16991 17663
rect 16991 17629 17000 17663
rect 16948 17620 17000 17629
rect 18144 17620 18196 17672
rect 19248 17688 19300 17740
rect 11612 17552 11664 17604
rect 12256 17552 12308 17604
rect 12440 17552 12492 17604
rect 16856 17552 16908 17604
rect 18604 17552 18656 17604
rect 22468 17552 22520 17604
rect 14372 17484 14424 17536
rect 19800 17484 19852 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 7380 17280 7432 17332
rect 8392 17323 8444 17332
rect 8392 17289 8401 17323
rect 8401 17289 8435 17323
rect 8435 17289 8444 17323
rect 8392 17280 8444 17289
rect 9312 17280 9364 17332
rect 12440 17280 12492 17332
rect 13176 17280 13228 17332
rect 13360 17280 13412 17332
rect 15200 17280 15252 17332
rect 15384 17323 15436 17332
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 15568 17280 15620 17332
rect 20352 17280 20404 17332
rect 8760 17212 8812 17264
rect 8668 17144 8720 17196
rect 11612 17212 11664 17264
rect 12900 17212 12952 17264
rect 16120 17212 16172 17264
rect 11244 17187 11296 17196
rect 11244 17153 11253 17187
rect 11253 17153 11287 17187
rect 11287 17153 11296 17187
rect 11244 17144 11296 17153
rect 11888 17144 11940 17196
rect 13544 17144 13596 17196
rect 13912 17144 13964 17196
rect 15384 17144 15436 17196
rect 15752 17144 15804 17196
rect 15936 17187 15988 17196
rect 15936 17153 15945 17187
rect 15945 17153 15979 17187
rect 15979 17153 15988 17187
rect 15936 17144 15988 17153
rect 16948 17144 17000 17196
rect 19984 17187 20036 17196
rect 19984 17153 19993 17187
rect 19993 17153 20027 17187
rect 20027 17153 20036 17187
rect 19984 17144 20036 17153
rect 20904 17144 20956 17196
rect 11152 17119 11204 17128
rect 11152 17085 11161 17119
rect 11161 17085 11195 17119
rect 11195 17085 11204 17119
rect 11152 17076 11204 17085
rect 14004 17076 14056 17128
rect 14464 17076 14516 17128
rect 17316 17076 17368 17128
rect 17960 17076 18012 17128
rect 18052 17119 18104 17128
rect 18052 17085 18061 17119
rect 18061 17085 18095 17119
rect 18095 17085 18104 17119
rect 18052 17076 18104 17085
rect 7656 17008 7708 17060
rect 13452 17008 13504 17060
rect 15292 17008 15344 17060
rect 18604 17076 18656 17128
rect 18696 17076 18748 17128
rect 20536 17119 20588 17128
rect 20536 17085 20545 17119
rect 20545 17085 20579 17119
rect 20579 17085 20588 17119
rect 20536 17076 20588 17085
rect 18512 17008 18564 17060
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 9312 16940 9364 16992
rect 9680 16983 9732 16992
rect 9680 16949 9689 16983
rect 9689 16949 9723 16983
rect 9723 16949 9732 16983
rect 9680 16940 9732 16949
rect 10140 16983 10192 16992
rect 10140 16949 10149 16983
rect 10149 16949 10183 16983
rect 10183 16949 10192 16983
rect 10140 16940 10192 16949
rect 11060 16983 11112 16992
rect 11060 16949 11069 16983
rect 11069 16949 11103 16983
rect 11103 16949 11112 16983
rect 11060 16940 11112 16949
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 13544 16983 13596 16992
rect 13544 16949 13553 16983
rect 13553 16949 13587 16983
rect 13587 16949 13596 16983
rect 13544 16940 13596 16949
rect 16304 16940 16356 16992
rect 16580 16940 16632 16992
rect 17224 16940 17276 16992
rect 17960 16940 18012 16992
rect 18144 16940 18196 16992
rect 20996 17008 21048 17060
rect 19800 16940 19852 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 9036 16736 9088 16788
rect 13452 16779 13504 16788
rect 13452 16745 13461 16779
rect 13461 16745 13495 16779
rect 13495 16745 13504 16779
rect 13452 16736 13504 16745
rect 14188 16779 14240 16788
rect 14188 16745 14197 16779
rect 14197 16745 14231 16779
rect 14231 16745 14240 16779
rect 14188 16736 14240 16745
rect 6920 16668 6972 16720
rect 5816 16600 5868 16652
rect 7564 16600 7616 16652
rect 7656 16575 7708 16584
rect 7656 16541 7665 16575
rect 7665 16541 7699 16575
rect 7699 16541 7708 16575
rect 7656 16532 7708 16541
rect 10140 16668 10192 16720
rect 10876 16668 10928 16720
rect 13544 16668 13596 16720
rect 14372 16668 14424 16720
rect 18144 16736 18196 16788
rect 18512 16736 18564 16788
rect 14740 16668 14792 16720
rect 16120 16668 16172 16720
rect 20996 16736 21048 16788
rect 9128 16600 9180 16652
rect 10508 16600 10560 16652
rect 11796 16600 11848 16652
rect 8668 16575 8720 16584
rect 8668 16541 8677 16575
rect 8677 16541 8711 16575
rect 8711 16541 8720 16575
rect 8668 16532 8720 16541
rect 10416 16575 10468 16584
rect 10416 16541 10425 16575
rect 10425 16541 10459 16575
rect 10459 16541 10468 16575
rect 10416 16532 10468 16541
rect 7380 16396 7432 16448
rect 9496 16396 9548 16448
rect 10416 16396 10468 16448
rect 11152 16396 11204 16448
rect 12716 16532 12768 16584
rect 13636 16532 13688 16584
rect 13912 16532 13964 16584
rect 15200 16532 15252 16584
rect 15936 16575 15988 16584
rect 15936 16541 15945 16575
rect 15945 16541 15979 16575
rect 15979 16541 15988 16575
rect 16580 16600 16632 16652
rect 16948 16643 17000 16652
rect 16948 16609 16957 16643
rect 16957 16609 16991 16643
rect 16991 16609 17000 16643
rect 16948 16600 17000 16609
rect 17040 16600 17092 16652
rect 18512 16600 18564 16652
rect 19156 16600 19208 16652
rect 15936 16532 15988 16541
rect 19432 16532 19484 16584
rect 15660 16464 15712 16516
rect 17592 16464 17644 16516
rect 19708 16575 19760 16584
rect 19708 16541 19717 16575
rect 19717 16541 19751 16575
rect 19751 16541 19760 16575
rect 19708 16532 19760 16541
rect 19800 16575 19852 16584
rect 19800 16541 19809 16575
rect 19809 16541 19843 16575
rect 19843 16541 19852 16575
rect 19800 16532 19852 16541
rect 21916 16600 21968 16652
rect 12072 16439 12124 16448
rect 12072 16405 12081 16439
rect 12081 16405 12115 16439
rect 12115 16405 12124 16439
rect 12072 16396 12124 16405
rect 12164 16396 12216 16448
rect 16488 16396 16540 16448
rect 20444 16439 20496 16448
rect 20444 16405 20453 16439
rect 20453 16405 20487 16439
rect 20487 16405 20496 16439
rect 20444 16396 20496 16405
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 6920 15988 6972 16040
rect 7380 15988 7432 16040
rect 9680 16192 9732 16244
rect 10416 16192 10468 16244
rect 9496 16031 9548 16040
rect 9496 15997 9505 16031
rect 9505 15997 9539 16031
rect 9539 15997 9548 16031
rect 9496 15988 9548 15997
rect 12164 16124 12216 16176
rect 11612 16099 11664 16108
rect 11612 16065 11621 16099
rect 11621 16065 11655 16099
rect 11655 16065 11664 16099
rect 11612 16056 11664 16065
rect 8208 15895 8260 15904
rect 8208 15861 8217 15895
rect 8217 15861 8251 15895
rect 8251 15861 8260 15895
rect 8208 15852 8260 15861
rect 11152 15988 11204 16040
rect 11520 16031 11572 16040
rect 11520 15997 11529 16031
rect 11529 15997 11563 16031
rect 11563 15997 11572 16031
rect 11520 15988 11572 15997
rect 15292 16124 15344 16176
rect 15936 16124 15988 16176
rect 16488 16192 16540 16244
rect 19432 16235 19484 16244
rect 16856 16167 16908 16176
rect 16856 16133 16865 16167
rect 16865 16133 16899 16167
rect 16899 16133 16908 16167
rect 16856 16124 16908 16133
rect 16120 16056 16172 16108
rect 17500 16099 17552 16108
rect 17500 16065 17509 16099
rect 17509 16065 17543 16099
rect 17543 16065 17552 16099
rect 17500 16056 17552 16065
rect 19432 16201 19441 16235
rect 19441 16201 19475 16235
rect 19475 16201 19484 16235
rect 19432 16192 19484 16201
rect 19156 16124 19208 16176
rect 19892 16056 19944 16108
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 11244 15852 11296 15904
rect 13544 15988 13596 16040
rect 13728 15988 13780 16040
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 15200 15988 15252 16040
rect 16304 16031 16356 16040
rect 16304 15997 16313 16031
rect 16313 15997 16347 16031
rect 16347 15997 16356 16031
rect 16304 15988 16356 15997
rect 16580 15988 16632 16040
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 19800 15988 19852 16040
rect 20904 15988 20956 16040
rect 13084 15920 13136 15972
rect 12348 15852 12400 15904
rect 17408 15920 17460 15972
rect 17684 15920 17736 15972
rect 13912 15852 13964 15904
rect 14464 15852 14516 15904
rect 15568 15895 15620 15904
rect 15568 15861 15577 15895
rect 15577 15861 15611 15895
rect 15611 15861 15620 15895
rect 15568 15852 15620 15861
rect 15844 15895 15896 15904
rect 15844 15861 15853 15895
rect 15853 15861 15887 15895
rect 15887 15861 15896 15895
rect 15844 15852 15896 15861
rect 15936 15852 15988 15904
rect 16488 15852 16540 15904
rect 19156 15852 19208 15904
rect 20628 15852 20680 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 7656 15648 7708 15700
rect 11060 15648 11112 15700
rect 6920 15580 6972 15632
rect 9128 15580 9180 15632
rect 11244 15580 11296 15632
rect 11796 15580 11848 15632
rect 13912 15648 13964 15700
rect 14188 15648 14240 15700
rect 16856 15648 16908 15700
rect 17500 15648 17552 15700
rect 15568 15580 15620 15632
rect 15752 15623 15804 15632
rect 15752 15589 15761 15623
rect 15761 15589 15795 15623
rect 15795 15589 15804 15623
rect 15752 15580 15804 15589
rect 8116 15512 8168 15564
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 10048 15512 10100 15564
rect 12440 15512 12492 15564
rect 12808 15555 12860 15564
rect 12808 15521 12817 15555
rect 12817 15521 12851 15555
rect 12851 15521 12860 15555
rect 12808 15512 12860 15521
rect 16488 15555 16540 15564
rect 16488 15521 16497 15555
rect 16497 15521 16531 15555
rect 16531 15521 16540 15555
rect 16488 15512 16540 15521
rect 17684 15512 17736 15564
rect 18052 15512 18104 15564
rect 19432 15580 19484 15632
rect 20076 15555 20128 15564
rect 11888 15444 11940 15496
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 13544 15487 13596 15496
rect 12348 15444 12400 15453
rect 12900 15376 12952 15428
rect 11704 15351 11756 15360
rect 11704 15317 11713 15351
rect 11713 15317 11747 15351
rect 11747 15317 11756 15351
rect 11704 15308 11756 15317
rect 13544 15453 13553 15487
rect 13553 15453 13587 15487
rect 13587 15453 13596 15487
rect 13544 15444 13596 15453
rect 15568 15444 15620 15496
rect 16580 15487 16632 15496
rect 16580 15453 16589 15487
rect 16589 15453 16623 15487
rect 16623 15453 16632 15487
rect 16580 15444 16632 15453
rect 20076 15521 20085 15555
rect 20085 15521 20119 15555
rect 20119 15521 20128 15555
rect 20076 15512 20128 15521
rect 20260 15487 20312 15496
rect 20260 15453 20269 15487
rect 20269 15453 20303 15487
rect 20303 15453 20312 15487
rect 20260 15444 20312 15453
rect 13728 15308 13780 15360
rect 14924 15351 14976 15360
rect 14924 15317 14933 15351
rect 14933 15317 14967 15351
rect 14967 15317 14976 15351
rect 14924 15308 14976 15317
rect 20720 15376 20772 15428
rect 16856 15308 16908 15360
rect 19800 15351 19852 15360
rect 19800 15317 19809 15351
rect 19809 15317 19843 15351
rect 19843 15317 19852 15351
rect 19800 15308 19852 15317
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 8116 15104 8168 15156
rect 6184 15011 6236 15020
rect 6184 14977 6193 15011
rect 6193 14977 6227 15011
rect 6227 14977 6236 15011
rect 6184 14968 6236 14977
rect 6920 14968 6972 15020
rect 7380 14968 7432 15020
rect 9680 15104 9732 15156
rect 12808 15104 12860 15156
rect 20076 15104 20128 15156
rect 14924 15036 14976 15088
rect 11704 14968 11756 15020
rect 12440 14968 12492 15020
rect 13084 15011 13136 15020
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13084 14968 13136 14977
rect 13544 14968 13596 15020
rect 5540 14900 5592 14952
rect 6092 14943 6144 14952
rect 6092 14909 6101 14943
rect 6101 14909 6135 14943
rect 6135 14909 6144 14943
rect 6092 14900 6144 14909
rect 11152 14900 11204 14952
rect 15476 14968 15528 15020
rect 15936 14968 15988 15020
rect 16120 14968 16172 15020
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 20536 15036 20588 15088
rect 16856 14968 16908 14977
rect 17776 14968 17828 15020
rect 19800 14968 19852 15020
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 20996 14968 21048 15020
rect 15292 14900 15344 14952
rect 8300 14832 8352 14884
rect 8576 14832 8628 14884
rect 9036 14764 9088 14816
rect 9680 14764 9732 14816
rect 11704 14807 11756 14816
rect 11704 14773 11713 14807
rect 11713 14773 11747 14807
rect 11747 14773 11756 14807
rect 11704 14764 11756 14773
rect 12716 14764 12768 14816
rect 15016 14807 15068 14816
rect 15016 14773 15025 14807
rect 15025 14773 15059 14807
rect 15059 14773 15068 14807
rect 15016 14764 15068 14773
rect 15660 14764 15712 14816
rect 20168 14900 20220 14952
rect 20904 14832 20956 14884
rect 19248 14764 19300 14816
rect 19708 14764 19760 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 8576 14603 8628 14612
rect 8576 14569 8585 14603
rect 8585 14569 8619 14603
rect 8619 14569 8628 14603
rect 8576 14560 8628 14569
rect 9036 14603 9088 14612
rect 9036 14569 9045 14603
rect 9045 14569 9079 14603
rect 9079 14569 9088 14603
rect 9036 14560 9088 14569
rect 9680 14603 9732 14612
rect 9680 14569 9689 14603
rect 9689 14569 9723 14603
rect 9723 14569 9732 14603
rect 9680 14560 9732 14569
rect 12440 14603 12492 14612
rect 12440 14569 12449 14603
rect 12449 14569 12483 14603
rect 12483 14569 12492 14603
rect 12440 14560 12492 14569
rect 13084 14560 13136 14612
rect 15292 14603 15344 14612
rect 15292 14569 15301 14603
rect 15301 14569 15335 14603
rect 15335 14569 15344 14603
rect 15292 14560 15344 14569
rect 15660 14603 15712 14612
rect 15660 14569 15669 14603
rect 15669 14569 15703 14603
rect 15703 14569 15712 14603
rect 15660 14560 15712 14569
rect 15844 14560 15896 14612
rect 17684 14603 17736 14612
rect 17684 14569 17693 14603
rect 17693 14569 17727 14603
rect 17727 14569 17736 14603
rect 17684 14560 17736 14569
rect 6920 14492 6972 14544
rect 8208 14492 8260 14544
rect 11060 14492 11112 14544
rect 12348 14492 12400 14544
rect 13636 14492 13688 14544
rect 14556 14492 14608 14544
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 12072 14424 12124 14476
rect 13544 14424 13596 14476
rect 14372 14467 14424 14476
rect 14372 14433 14381 14467
rect 14381 14433 14415 14467
rect 14415 14433 14424 14467
rect 14372 14424 14424 14433
rect 10140 14399 10192 14408
rect 8300 14331 8352 14340
rect 8300 14297 8309 14331
rect 8309 14297 8343 14331
rect 8343 14297 8352 14331
rect 10140 14365 10149 14399
rect 10149 14365 10183 14399
rect 10183 14365 10192 14399
rect 10140 14356 10192 14365
rect 8300 14288 8352 14297
rect 9220 14220 9272 14272
rect 15568 14356 15620 14408
rect 16212 14356 16264 14408
rect 17592 14424 17644 14476
rect 19800 14492 19852 14544
rect 20260 14467 20312 14476
rect 20260 14433 20269 14467
rect 20269 14433 20303 14467
rect 20303 14433 20312 14467
rect 20260 14424 20312 14433
rect 17960 14399 18012 14408
rect 17960 14365 17969 14399
rect 17969 14365 18003 14399
rect 18003 14365 18012 14399
rect 17960 14356 18012 14365
rect 20076 14356 20128 14408
rect 10508 14220 10560 14272
rect 13636 14220 13688 14272
rect 19984 14263 20036 14272
rect 19984 14229 19993 14263
rect 19993 14229 20027 14263
rect 20027 14229 20036 14263
rect 19984 14220 20036 14229
rect 20444 14263 20496 14272
rect 20444 14229 20453 14263
rect 20453 14229 20487 14263
rect 20487 14229 20496 14263
rect 20444 14220 20496 14229
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 11704 14016 11756 14068
rect 12716 14059 12768 14068
rect 12716 14025 12725 14059
rect 12725 14025 12759 14059
rect 12759 14025 12768 14059
rect 12716 14016 12768 14025
rect 16488 14016 16540 14068
rect 16948 14016 17000 14068
rect 17592 14059 17644 14068
rect 15752 13948 15804 14000
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 19708 14059 19760 14068
rect 19708 14025 19717 14059
rect 19717 14025 19751 14059
rect 19751 14025 19760 14059
rect 19708 14016 19760 14025
rect 20904 14059 20956 14068
rect 20904 14025 20913 14059
rect 20913 14025 20947 14059
rect 20947 14025 20956 14059
rect 20904 14016 20956 14025
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 11796 13923 11848 13932
rect 11796 13889 11805 13923
rect 11805 13889 11839 13923
rect 11839 13889 11848 13923
rect 11796 13880 11848 13889
rect 12348 13880 12400 13932
rect 13176 13923 13228 13932
rect 13176 13889 13185 13923
rect 13185 13889 13219 13923
rect 13219 13889 13228 13923
rect 13176 13880 13228 13889
rect 13544 13880 13596 13932
rect 14188 13923 14240 13932
rect 14188 13889 14197 13923
rect 14197 13889 14231 13923
rect 14231 13889 14240 13923
rect 14188 13880 14240 13889
rect 13636 13812 13688 13864
rect 13728 13812 13780 13864
rect 15016 13880 15068 13932
rect 15568 13923 15620 13932
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 15844 13812 15896 13864
rect 16304 13812 16356 13864
rect 16856 13812 16908 13864
rect 19064 13812 19116 13864
rect 19800 13880 19852 13932
rect 20720 13855 20772 13864
rect 20720 13821 20729 13855
rect 20729 13821 20763 13855
rect 20763 13821 20772 13855
rect 20720 13812 20772 13821
rect 10048 13744 10100 13796
rect 9588 13676 9640 13728
rect 10600 13719 10652 13728
rect 10600 13685 10609 13719
rect 10609 13685 10643 13719
rect 10643 13685 10652 13719
rect 10600 13676 10652 13685
rect 14096 13719 14148 13728
rect 14096 13685 14105 13719
rect 14105 13685 14139 13719
rect 14139 13685 14148 13719
rect 14096 13676 14148 13685
rect 14556 13676 14608 13728
rect 15292 13719 15344 13728
rect 15292 13685 15301 13719
rect 15301 13685 15335 13719
rect 15335 13685 15344 13719
rect 15292 13676 15344 13685
rect 15476 13744 15528 13796
rect 15660 13744 15712 13796
rect 16672 13744 16724 13796
rect 18788 13744 18840 13796
rect 20076 13787 20128 13796
rect 20076 13753 20085 13787
rect 20085 13753 20119 13787
rect 20119 13753 20128 13787
rect 20076 13744 20128 13753
rect 18052 13719 18104 13728
rect 18052 13685 18061 13719
rect 18061 13685 18095 13719
rect 18095 13685 18104 13719
rect 18052 13676 18104 13685
rect 18420 13719 18472 13728
rect 18420 13685 18429 13719
rect 18429 13685 18463 13719
rect 18463 13685 18472 13719
rect 18420 13676 18472 13685
rect 18696 13676 18748 13728
rect 18972 13676 19024 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 10968 13472 11020 13524
rect 11612 13472 11664 13524
rect 11980 13472 12032 13524
rect 13176 13515 13228 13524
rect 13176 13481 13185 13515
rect 13185 13481 13219 13515
rect 13219 13481 13228 13515
rect 13176 13472 13228 13481
rect 14556 13515 14608 13524
rect 14556 13481 14565 13515
rect 14565 13481 14599 13515
rect 14599 13481 14608 13515
rect 14556 13472 14608 13481
rect 17040 13472 17092 13524
rect 18052 13472 18104 13524
rect 20168 13472 20220 13524
rect 11060 13404 11112 13456
rect 11796 13404 11848 13456
rect 13636 13404 13688 13456
rect 13820 13404 13872 13456
rect 14004 13404 14056 13456
rect 14096 13404 14148 13456
rect 15752 13404 15804 13456
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 12348 13379 12400 13388
rect 12348 13345 12357 13379
rect 12357 13345 12391 13379
rect 12391 13345 12400 13379
rect 12348 13336 12400 13345
rect 12532 13336 12584 13388
rect 13176 13336 13228 13388
rect 13728 13336 13780 13388
rect 16396 13336 16448 13388
rect 16580 13336 16632 13388
rect 17592 13336 17644 13388
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 10600 13268 10652 13320
rect 11060 13200 11112 13252
rect 12624 13311 12676 13320
rect 12624 13277 12633 13311
rect 12633 13277 12667 13311
rect 12667 13277 12676 13311
rect 12624 13268 12676 13277
rect 13544 13200 13596 13252
rect 14004 13268 14056 13320
rect 14740 13311 14792 13320
rect 14740 13277 14749 13311
rect 14749 13277 14783 13311
rect 14783 13277 14792 13311
rect 14740 13268 14792 13277
rect 16856 13268 16908 13320
rect 17684 13268 17736 13320
rect 18972 13336 19024 13388
rect 19432 13336 19484 13388
rect 19248 13311 19300 13320
rect 19248 13277 19257 13311
rect 19257 13277 19291 13311
rect 19291 13277 19300 13311
rect 19248 13268 19300 13277
rect 20260 13311 20312 13320
rect 16672 13200 16724 13252
rect 17224 13200 17276 13252
rect 18420 13200 18472 13252
rect 19064 13200 19116 13252
rect 20260 13277 20269 13311
rect 20269 13277 20303 13311
rect 20303 13277 20312 13311
rect 20260 13268 20312 13277
rect 19984 13200 20036 13252
rect 10784 13175 10836 13184
rect 10784 13141 10793 13175
rect 10793 13141 10827 13175
rect 10827 13141 10836 13175
rect 10784 13132 10836 13141
rect 12440 13132 12492 13184
rect 13820 13132 13872 13184
rect 15752 13175 15804 13184
rect 15752 13141 15761 13175
rect 15761 13141 15795 13175
rect 15795 13141 15804 13175
rect 15752 13132 15804 13141
rect 16304 13132 16356 13184
rect 17776 13132 17828 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 9220 12928 9272 12980
rect 11060 12971 11112 12980
rect 8484 12792 8536 12844
rect 11060 12937 11069 12971
rect 11069 12937 11103 12971
rect 11103 12937 11112 12971
rect 11060 12928 11112 12937
rect 14280 12928 14332 12980
rect 10876 12860 10928 12912
rect 12072 12903 12124 12912
rect 10784 12792 10836 12844
rect 12072 12869 12081 12903
rect 12081 12869 12115 12903
rect 12115 12869 12124 12903
rect 15844 12928 15896 12980
rect 16580 12971 16632 12980
rect 16580 12937 16589 12971
rect 16589 12937 16623 12971
rect 16623 12937 16632 12971
rect 16580 12928 16632 12937
rect 18604 12928 18656 12980
rect 19064 12928 19116 12980
rect 12072 12860 12124 12869
rect 16212 12860 16264 12912
rect 12992 12792 13044 12844
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 10600 12724 10652 12776
rect 11888 12724 11940 12776
rect 12164 12724 12216 12776
rect 10508 12656 10560 12708
rect 11428 12699 11480 12708
rect 11428 12665 11437 12699
rect 11437 12665 11471 12699
rect 11471 12665 11480 12699
rect 11428 12656 11480 12665
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 14188 12724 14240 12776
rect 13360 12656 13412 12708
rect 14372 12588 14424 12640
rect 15752 12792 15804 12844
rect 17592 12792 17644 12844
rect 18604 12792 18656 12844
rect 19800 12792 19852 12844
rect 16488 12724 16540 12776
rect 17960 12724 18012 12776
rect 18144 12767 18196 12776
rect 18144 12733 18153 12767
rect 18153 12733 18187 12767
rect 18187 12733 18196 12767
rect 18144 12724 18196 12733
rect 19984 12724 20036 12776
rect 14556 12656 14608 12708
rect 14740 12656 14792 12708
rect 17592 12656 17644 12708
rect 15752 12631 15804 12640
rect 15752 12597 15761 12631
rect 15761 12597 15795 12631
rect 15795 12597 15804 12631
rect 15752 12588 15804 12597
rect 15844 12588 15896 12640
rect 16212 12631 16264 12640
rect 16212 12597 16221 12631
rect 16221 12597 16255 12631
rect 16255 12597 16264 12631
rect 16212 12588 16264 12597
rect 20628 12656 20680 12708
rect 20536 12588 20588 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 10324 12316 10376 12368
rect 12624 12384 12676 12436
rect 16948 12384 17000 12436
rect 17868 12427 17920 12436
rect 17868 12393 17877 12427
rect 17877 12393 17911 12427
rect 17911 12393 17920 12427
rect 17868 12384 17920 12393
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 20444 12427 20496 12436
rect 20444 12393 20453 12427
rect 20453 12393 20487 12427
rect 20487 12393 20496 12427
rect 20444 12384 20496 12393
rect 13820 12316 13872 12368
rect 15752 12316 15804 12368
rect 17960 12316 18012 12368
rect 18420 12316 18472 12368
rect 8484 12248 8536 12300
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 9496 12180 9548 12232
rect 9404 12112 9456 12164
rect 10876 12248 10928 12300
rect 12256 12248 12308 12300
rect 12532 12248 12584 12300
rect 18144 12248 18196 12300
rect 19248 12248 19300 12300
rect 9036 12044 9088 12096
rect 13360 12180 13412 12232
rect 11796 12044 11848 12096
rect 15108 12180 15160 12232
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 18604 12223 18656 12232
rect 14556 12044 14608 12096
rect 17132 12087 17184 12096
rect 17132 12053 17141 12087
rect 17141 12053 17175 12087
rect 17175 12053 17184 12087
rect 17132 12044 17184 12053
rect 17224 12044 17276 12096
rect 17868 12044 17920 12096
rect 18604 12189 18613 12223
rect 18613 12189 18647 12223
rect 18647 12189 18656 12223
rect 18604 12180 18656 12189
rect 19616 12180 19668 12232
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 10140 11840 10192 11892
rect 12348 11840 12400 11892
rect 13544 11840 13596 11892
rect 15844 11840 15896 11892
rect 19432 11840 19484 11892
rect 8852 11747 8904 11756
rect 8852 11713 8861 11747
rect 8861 11713 8895 11747
rect 8895 11713 8904 11747
rect 8852 11704 8904 11713
rect 14096 11772 14148 11824
rect 10876 11747 10928 11756
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 12256 11704 12308 11756
rect 9496 11636 9548 11688
rect 11796 11636 11848 11688
rect 12532 11568 12584 11620
rect 12624 11568 12676 11620
rect 13360 11568 13412 11620
rect 15568 11704 15620 11756
rect 17684 11704 17736 11756
rect 17224 11679 17276 11688
rect 17224 11645 17233 11679
rect 17233 11645 17267 11679
rect 17267 11645 17276 11679
rect 17224 11636 17276 11645
rect 18236 11772 18288 11824
rect 18604 11772 18656 11824
rect 18696 11704 18748 11756
rect 19248 11747 19300 11756
rect 19248 11713 19257 11747
rect 19257 11713 19291 11747
rect 19291 11713 19300 11747
rect 19248 11704 19300 11713
rect 19616 11636 19668 11688
rect 15292 11568 15344 11620
rect 15476 11568 15528 11620
rect 18512 11568 18564 11620
rect 18696 11568 18748 11620
rect 18880 11568 18932 11620
rect 19984 11611 20036 11620
rect 19984 11577 20018 11611
rect 20018 11577 20036 11611
rect 19984 11568 20036 11577
rect 8668 11543 8720 11552
rect 8668 11509 8677 11543
rect 8677 11509 8711 11543
rect 8711 11509 8720 11543
rect 8668 11500 8720 11509
rect 8760 11543 8812 11552
rect 8760 11509 8769 11543
rect 8769 11509 8803 11543
rect 8803 11509 8812 11543
rect 8760 11500 8812 11509
rect 11428 11500 11480 11552
rect 11704 11543 11756 11552
rect 11704 11509 11713 11543
rect 11713 11509 11747 11543
rect 11747 11509 11756 11543
rect 11704 11500 11756 11509
rect 12440 11500 12492 11552
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 14280 11543 14332 11552
rect 14280 11509 14289 11543
rect 14289 11509 14323 11543
rect 14323 11509 14332 11543
rect 14280 11500 14332 11509
rect 15016 11500 15068 11552
rect 15752 11543 15804 11552
rect 15752 11509 15761 11543
rect 15761 11509 15795 11543
rect 15795 11509 15804 11543
rect 15752 11500 15804 11509
rect 16212 11500 16264 11552
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 17316 11543 17368 11552
rect 16856 11500 16908 11509
rect 17316 11509 17325 11543
rect 17325 11509 17359 11543
rect 17359 11509 17368 11543
rect 17316 11500 17368 11509
rect 18604 11500 18656 11552
rect 19248 11500 19300 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 8668 11296 8720 11348
rect 10140 11271 10192 11280
rect 10140 11237 10149 11271
rect 10149 11237 10183 11271
rect 10183 11237 10192 11271
rect 10140 11228 10192 11237
rect 10232 11271 10284 11280
rect 10232 11237 10241 11271
rect 10241 11237 10275 11271
rect 10275 11237 10284 11271
rect 10232 11228 10284 11237
rect 10600 11228 10652 11280
rect 11704 11296 11756 11348
rect 14004 11296 14056 11348
rect 14188 11296 14240 11348
rect 15660 11296 15712 11348
rect 16580 11296 16632 11348
rect 17868 11296 17920 11348
rect 20260 11296 20312 11348
rect 7472 11160 7524 11212
rect 9036 11160 9088 11212
rect 9404 11160 9456 11212
rect 11060 11203 11112 11212
rect 11060 11169 11094 11203
rect 11094 11169 11112 11203
rect 13268 11228 13320 11280
rect 18604 11228 18656 11280
rect 19248 11228 19300 11280
rect 19340 11228 19392 11280
rect 11060 11160 11112 11169
rect 13820 11160 13872 11212
rect 15568 11160 15620 11212
rect 13728 11092 13780 11144
rect 14004 11092 14056 11144
rect 17224 11160 17276 11212
rect 17408 11160 17460 11212
rect 8668 11024 8720 11076
rect 8852 11024 8904 11076
rect 13820 11024 13872 11076
rect 15844 11024 15896 11076
rect 12256 10956 12308 11008
rect 15568 10999 15620 11008
rect 15568 10965 15577 10999
rect 15577 10965 15611 10999
rect 15611 10965 15620 10999
rect 15568 10956 15620 10965
rect 18604 11092 18656 11144
rect 18972 11092 19024 11144
rect 19708 11160 19760 11212
rect 20260 11135 20312 11144
rect 19064 11024 19116 11076
rect 20260 11101 20269 11135
rect 20269 11101 20303 11135
rect 20303 11101 20312 11135
rect 20260 11092 20312 11101
rect 16948 10956 17000 11008
rect 18788 10999 18840 11008
rect 18788 10965 18797 10999
rect 18797 10965 18831 10999
rect 18831 10965 18840 10999
rect 18788 10956 18840 10965
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 8760 10752 8812 10804
rect 11980 10752 12032 10804
rect 12348 10752 12400 10804
rect 12440 10795 12492 10804
rect 12440 10761 12449 10795
rect 12449 10761 12483 10795
rect 12483 10761 12492 10795
rect 12440 10752 12492 10761
rect 14280 10752 14332 10804
rect 17316 10752 17368 10804
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 9128 10548 9180 10600
rect 12624 10684 12676 10736
rect 15200 10684 15252 10736
rect 11152 10659 11204 10668
rect 11152 10625 11161 10659
rect 11161 10625 11195 10659
rect 11195 10625 11204 10659
rect 11152 10616 11204 10625
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 12256 10616 12308 10668
rect 15292 10616 15344 10668
rect 8576 10480 8628 10532
rect 14280 10548 14332 10600
rect 14096 10480 14148 10532
rect 15200 10480 15252 10532
rect 15568 10548 15620 10600
rect 17960 10616 18012 10668
rect 16580 10591 16632 10600
rect 16580 10557 16614 10591
rect 16614 10557 16632 10591
rect 16212 10480 16264 10532
rect 16580 10548 16632 10557
rect 16672 10480 16724 10532
rect 16948 10480 17000 10532
rect 8944 10412 8996 10464
rect 10968 10455 11020 10464
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 11060 10455 11112 10464
rect 11060 10421 11069 10455
rect 11069 10421 11103 10455
rect 11103 10421 11112 10455
rect 11060 10412 11112 10421
rect 12624 10412 12676 10464
rect 13268 10412 13320 10464
rect 13544 10412 13596 10464
rect 13728 10412 13780 10464
rect 13820 10412 13872 10464
rect 17868 10548 17920 10600
rect 18788 10548 18840 10600
rect 19340 10548 19392 10600
rect 17132 10480 17184 10532
rect 20536 10480 20588 10532
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 18972 10412 19024 10464
rect 20628 10412 20680 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 10600 10208 10652 10260
rect 11244 10208 11296 10260
rect 8668 10140 8720 10192
rect 11152 10140 11204 10192
rect 13360 10208 13412 10260
rect 13820 10251 13872 10260
rect 13820 10217 13829 10251
rect 13829 10217 13863 10251
rect 13863 10217 13872 10251
rect 13820 10208 13872 10217
rect 14372 10251 14424 10260
rect 14372 10217 14381 10251
rect 14381 10217 14415 10251
rect 14415 10217 14424 10251
rect 14372 10208 14424 10217
rect 15016 10208 15068 10260
rect 15476 10208 15528 10260
rect 17132 10251 17184 10260
rect 17132 10217 17141 10251
rect 17141 10217 17175 10251
rect 17175 10217 17184 10251
rect 17132 10208 17184 10217
rect 17592 10251 17644 10260
rect 17592 10217 17601 10251
rect 17601 10217 17635 10251
rect 17635 10217 17644 10251
rect 17592 10208 17644 10217
rect 20260 10208 20312 10260
rect 20536 10251 20588 10260
rect 20536 10217 20545 10251
rect 20545 10217 20579 10251
rect 20579 10217 20588 10251
rect 20536 10208 20588 10217
rect 12256 10140 12308 10192
rect 15108 10140 15160 10192
rect 16764 10140 16816 10192
rect 18788 10140 18840 10192
rect 19984 10140 20036 10192
rect 20628 10140 20680 10192
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 8760 9936 8812 9988
rect 9220 9936 9272 9988
rect 13636 10004 13688 10056
rect 14556 10004 14608 10056
rect 9128 9868 9180 9920
rect 12716 9868 12768 9920
rect 14372 9936 14424 9988
rect 16856 10072 16908 10124
rect 18512 10115 18564 10124
rect 15384 9936 15436 9988
rect 18512 10081 18521 10115
rect 18521 10081 18555 10115
rect 18555 10081 18564 10115
rect 18512 10072 18564 10081
rect 18420 10004 18472 10056
rect 18788 10047 18840 10056
rect 18788 10013 18797 10047
rect 18797 10013 18831 10047
rect 18831 10013 18840 10047
rect 18788 10004 18840 10013
rect 19064 9936 19116 9988
rect 19340 9868 19392 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 15292 9664 15344 9716
rect 17132 9664 17184 9716
rect 17776 9664 17828 9716
rect 18512 9664 18564 9716
rect 18788 9664 18840 9716
rect 11152 9639 11204 9648
rect 11152 9605 11161 9639
rect 11161 9605 11195 9639
rect 11195 9605 11204 9639
rect 11152 9596 11204 9605
rect 16212 9639 16264 9648
rect 16212 9605 16221 9639
rect 16221 9605 16255 9639
rect 16255 9605 16264 9639
rect 16212 9596 16264 9605
rect 17960 9596 18012 9648
rect 18328 9596 18380 9648
rect 19340 9664 19392 9716
rect 7656 9528 7708 9580
rect 10416 9460 10468 9512
rect 12348 9460 12400 9512
rect 12532 9460 12584 9512
rect 14188 9460 14240 9512
rect 14648 9460 14700 9512
rect 9128 9392 9180 9444
rect 11244 9392 11296 9444
rect 15292 9460 15344 9512
rect 17224 9528 17276 9580
rect 16028 9460 16080 9512
rect 20444 9571 20496 9580
rect 20444 9537 20453 9571
rect 20453 9537 20487 9571
rect 20487 9537 20496 9571
rect 20444 9528 20496 9537
rect 20628 9571 20680 9580
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 18972 9460 19024 9512
rect 15844 9392 15896 9444
rect 16488 9392 16540 9444
rect 18420 9435 18472 9444
rect 18420 9401 18429 9435
rect 18429 9401 18463 9435
rect 18463 9401 18472 9435
rect 18420 9392 18472 9401
rect 9220 9324 9272 9376
rect 11428 9367 11480 9376
rect 11428 9333 11437 9367
rect 11437 9333 11471 9367
rect 11471 9333 11480 9367
rect 11428 9324 11480 9333
rect 12072 9324 12124 9376
rect 13544 9324 13596 9376
rect 13636 9324 13688 9376
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 15568 9324 15620 9376
rect 17408 9324 17460 9376
rect 17592 9324 17644 9376
rect 18512 9367 18564 9376
rect 18512 9333 18521 9367
rect 18521 9333 18555 9367
rect 18555 9333 18564 9367
rect 18512 9324 18564 9333
rect 19892 9324 19944 9376
rect 20352 9367 20404 9376
rect 20352 9333 20361 9367
rect 20361 9333 20395 9367
rect 20395 9333 20404 9367
rect 20352 9324 20404 9333
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 8576 9163 8628 9172
rect 8576 9129 8585 9163
rect 8585 9129 8619 9163
rect 8619 9129 8628 9163
rect 8576 9120 8628 9129
rect 9680 9120 9732 9172
rect 10416 9163 10468 9172
rect 10416 9129 10425 9163
rect 10425 9129 10459 9163
rect 10459 9129 10468 9163
rect 10416 9120 10468 9129
rect 10968 9120 11020 9172
rect 11428 9120 11480 9172
rect 3424 9052 3476 9104
rect 12532 9052 12584 9104
rect 13636 9052 13688 9104
rect 15200 9120 15252 9172
rect 15476 9120 15528 9172
rect 17960 9120 18012 9172
rect 10968 8984 11020 9036
rect 11152 9027 11204 9036
rect 8576 8916 8628 8968
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 12348 8984 12400 9036
rect 13544 8984 13596 9036
rect 15936 8984 15988 9036
rect 16948 9027 17000 9036
rect 16948 8993 16957 9027
rect 16957 8993 16991 9027
rect 16991 8993 17000 9027
rect 16948 8984 17000 8993
rect 17684 9052 17736 9104
rect 19248 9120 19300 9172
rect 19800 9052 19852 9104
rect 20076 8984 20128 9036
rect 8208 8848 8260 8900
rect 11244 8959 11296 8968
rect 11244 8925 11253 8959
rect 11253 8925 11287 8959
rect 11287 8925 11296 8959
rect 11244 8916 11296 8925
rect 10784 8848 10836 8900
rect 15660 8916 15712 8968
rect 15844 8959 15896 8968
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 15568 8848 15620 8900
rect 16672 8848 16724 8900
rect 18328 8916 18380 8968
rect 11704 8823 11756 8832
rect 11704 8789 11713 8823
rect 11713 8789 11747 8823
rect 11747 8789 11756 8823
rect 11704 8780 11756 8789
rect 14188 8823 14240 8832
rect 14188 8789 14197 8823
rect 14197 8789 14231 8823
rect 14231 8789 14240 8823
rect 14188 8780 14240 8789
rect 14740 8780 14792 8832
rect 15108 8780 15160 8832
rect 16488 8780 16540 8832
rect 17776 8780 17828 8832
rect 19064 8780 19116 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 8576 8619 8628 8628
rect 8576 8585 8585 8619
rect 8585 8585 8619 8619
rect 8619 8585 8628 8619
rect 8576 8576 8628 8585
rect 11060 8576 11112 8628
rect 10968 8508 11020 8560
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 9588 8372 9640 8424
rect 10416 8372 10468 8424
rect 10876 8372 10928 8424
rect 11152 8372 11204 8424
rect 11704 8415 11756 8424
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 14096 8508 14148 8560
rect 13636 8440 13688 8492
rect 14740 8483 14792 8492
rect 14740 8449 14749 8483
rect 14749 8449 14783 8483
rect 14783 8449 14792 8483
rect 14740 8440 14792 8449
rect 14280 8372 14332 8424
rect 15292 8372 15344 8424
rect 15844 8576 15896 8628
rect 15568 8483 15620 8492
rect 15568 8449 15577 8483
rect 15577 8449 15611 8483
rect 15611 8449 15620 8483
rect 15568 8440 15620 8449
rect 16580 8440 16632 8492
rect 6920 8304 6972 8356
rect 10784 8304 10836 8356
rect 11244 8304 11296 8356
rect 12072 8304 12124 8356
rect 13728 8304 13780 8356
rect 14372 8304 14424 8356
rect 15016 8304 15068 8356
rect 16948 8372 17000 8424
rect 11152 8236 11204 8288
rect 13176 8279 13228 8288
rect 13176 8245 13185 8279
rect 13185 8245 13219 8279
rect 13219 8245 13228 8279
rect 13176 8236 13228 8245
rect 13268 8236 13320 8288
rect 14280 8236 14332 8288
rect 16304 8304 16356 8356
rect 15292 8236 15344 8288
rect 18144 8304 18196 8356
rect 18604 8576 18656 8628
rect 19800 8508 19852 8560
rect 18604 8483 18656 8492
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 18604 8440 18656 8449
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20076 8440 20128 8449
rect 19892 8415 19944 8424
rect 19892 8381 19901 8415
rect 19901 8381 19935 8415
rect 19935 8381 19944 8415
rect 19892 8372 19944 8381
rect 17224 8279 17276 8288
rect 17224 8245 17233 8279
rect 17233 8245 17267 8279
rect 17267 8245 17276 8279
rect 17224 8236 17276 8245
rect 17960 8236 18012 8288
rect 19984 8279 20036 8288
rect 19984 8245 19993 8279
rect 19993 8245 20027 8279
rect 20027 8245 20036 8279
rect 19984 8236 20036 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 11152 8032 11204 8084
rect 9680 7896 9732 7948
rect 11060 7896 11112 7948
rect 13636 7964 13688 8016
rect 14188 7964 14240 8016
rect 14096 7896 14148 7948
rect 18052 8032 18104 8084
rect 20076 8032 20128 8084
rect 20352 8032 20404 8084
rect 18604 7964 18656 8016
rect 16764 7896 16816 7948
rect 17776 7896 17828 7948
rect 20628 7896 20680 7948
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 10876 7828 10928 7880
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 16304 7871 16356 7880
rect 11796 7692 11848 7744
rect 12072 7692 12124 7744
rect 13268 7692 13320 7744
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 16672 7871 16724 7880
rect 16672 7837 16681 7871
rect 16681 7837 16715 7871
rect 16715 7837 16724 7871
rect 16672 7828 16724 7837
rect 17776 7692 17828 7744
rect 17868 7692 17920 7744
rect 18788 7692 18840 7744
rect 19064 7692 19116 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 9312 7488 9364 7540
rect 10784 7488 10836 7540
rect 12072 7352 12124 7404
rect 13544 7420 13596 7472
rect 15200 7420 15252 7472
rect 16304 7488 16356 7540
rect 16764 7488 16816 7540
rect 17776 7488 17828 7540
rect 19984 7488 20036 7540
rect 13636 7352 13688 7404
rect 14188 7352 14240 7404
rect 17408 7420 17460 7472
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 13176 7284 13228 7336
rect 13820 7284 13872 7336
rect 17868 7352 17920 7404
rect 18696 7352 18748 7404
rect 17224 7284 17276 7336
rect 17960 7284 18012 7336
rect 18512 7284 18564 7336
rect 19432 7327 19484 7336
rect 9404 7259 9456 7268
rect 9404 7225 9438 7259
rect 9438 7225 9456 7259
rect 9404 7216 9456 7225
rect 12256 7148 12308 7200
rect 13912 7216 13964 7268
rect 16580 7216 16632 7268
rect 18512 7191 18564 7200
rect 18512 7157 18521 7191
rect 18521 7157 18555 7191
rect 18555 7157 18564 7191
rect 18512 7148 18564 7157
rect 19432 7293 19441 7327
rect 19441 7293 19475 7327
rect 19475 7293 19484 7327
rect 19432 7284 19484 7293
rect 20628 7395 20680 7404
rect 20628 7361 20637 7395
rect 20637 7361 20671 7395
rect 20671 7361 20680 7395
rect 20628 7352 20680 7361
rect 19248 7148 19300 7200
rect 20444 7191 20496 7200
rect 20444 7157 20453 7191
rect 20453 7157 20487 7191
rect 20487 7157 20496 7191
rect 20444 7148 20496 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 9680 6987 9732 6996
rect 9680 6953 9689 6987
rect 9689 6953 9723 6987
rect 9723 6953 9732 6987
rect 9680 6944 9732 6953
rect 14372 6944 14424 6996
rect 9128 6876 9180 6928
rect 7656 6740 7708 6792
rect 9036 6808 9088 6860
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 10324 6808 10376 6860
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 12072 6876 12124 6928
rect 15384 6876 15436 6928
rect 18604 6944 18656 6996
rect 20628 6944 20680 6996
rect 19892 6876 19944 6928
rect 13452 6808 13504 6860
rect 14004 6808 14056 6860
rect 14464 6808 14516 6860
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 18696 6808 18748 6860
rect 19432 6851 19484 6860
rect 19432 6817 19466 6851
rect 19466 6817 19484 6851
rect 19432 6808 19484 6817
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 9404 6672 9456 6724
rect 9128 6604 9180 6656
rect 10876 6604 10928 6656
rect 10968 6604 11020 6656
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 15292 6740 15344 6792
rect 15936 6783 15988 6792
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 15936 6740 15988 6749
rect 16304 6783 16356 6792
rect 16304 6749 16313 6783
rect 16313 6749 16347 6783
rect 16347 6749 16356 6783
rect 16304 6740 16356 6749
rect 13728 6715 13780 6724
rect 13728 6681 13737 6715
rect 13737 6681 13771 6715
rect 13771 6681 13780 6715
rect 13728 6672 13780 6681
rect 15200 6672 15252 6724
rect 14096 6604 14148 6656
rect 16120 6604 16172 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 9036 6443 9088 6452
rect 9036 6409 9045 6443
rect 9045 6409 9079 6443
rect 9079 6409 9088 6443
rect 9036 6400 9088 6409
rect 10048 6400 10100 6452
rect 10140 6400 10192 6452
rect 10968 6400 11020 6452
rect 11060 6400 11112 6452
rect 13544 6400 13596 6452
rect 15292 6443 15344 6452
rect 15292 6409 15301 6443
rect 15301 6409 15335 6443
rect 15335 6409 15344 6443
rect 15292 6400 15344 6409
rect 16396 6400 16448 6452
rect 6092 6264 6144 6316
rect 10232 6332 10284 6384
rect 12072 6332 12124 6384
rect 12440 6332 12492 6384
rect 18512 6400 18564 6452
rect 7656 6239 7708 6248
rect 7656 6205 7665 6239
rect 7665 6205 7699 6239
rect 7699 6205 7708 6239
rect 7656 6196 7708 6205
rect 10968 6264 11020 6316
rect 12992 6307 13044 6316
rect 12992 6273 13001 6307
rect 13001 6273 13035 6307
rect 13035 6273 13044 6307
rect 12992 6264 13044 6273
rect 14096 6307 14148 6316
rect 14096 6273 14105 6307
rect 14105 6273 14139 6307
rect 14139 6273 14148 6307
rect 14096 6264 14148 6273
rect 15476 6264 15528 6316
rect 15936 6264 15988 6316
rect 16488 6264 16540 6316
rect 7748 6128 7800 6180
rect 9128 6128 9180 6180
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 10784 6103 10836 6112
rect 10784 6069 10793 6103
rect 10793 6069 10827 6103
rect 10827 6069 10836 6103
rect 10784 6060 10836 6069
rect 12164 6196 12216 6248
rect 15660 6196 15712 6248
rect 15752 6196 15804 6248
rect 16028 6196 16080 6248
rect 16304 6196 16356 6248
rect 12348 6060 12400 6112
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12900 6103 12952 6112
rect 12440 6060 12492 6069
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 13544 6128 13596 6180
rect 15292 6128 15344 6180
rect 14004 6060 14056 6112
rect 16396 6128 16448 6180
rect 20720 6332 20772 6384
rect 18604 6307 18656 6316
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 18604 6264 18656 6273
rect 19708 6307 19760 6316
rect 19708 6273 19717 6307
rect 19717 6273 19751 6307
rect 19751 6273 19760 6307
rect 19708 6264 19760 6273
rect 20168 6264 20220 6316
rect 20352 6264 20404 6316
rect 18420 6239 18472 6248
rect 18420 6205 18429 6239
rect 18429 6205 18463 6239
rect 18463 6205 18472 6239
rect 18420 6196 18472 6205
rect 19064 6196 19116 6248
rect 18972 6128 19024 6180
rect 15752 6103 15804 6112
rect 15752 6069 15761 6103
rect 15761 6069 15795 6103
rect 15795 6069 15804 6103
rect 16304 6103 16356 6112
rect 15752 6060 15804 6069
rect 16304 6069 16313 6103
rect 16313 6069 16347 6103
rect 16347 6069 16356 6103
rect 16304 6060 16356 6069
rect 16672 6060 16724 6112
rect 18604 6060 18656 6112
rect 19616 6103 19668 6112
rect 19616 6069 19625 6103
rect 19625 6069 19659 6103
rect 19659 6069 19668 6103
rect 19616 6060 19668 6069
rect 20260 6103 20312 6112
rect 20260 6069 20269 6103
rect 20269 6069 20303 6103
rect 20303 6069 20312 6103
rect 20260 6060 20312 6069
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 7748 5856 7800 5908
rect 9128 5899 9180 5908
rect 4068 5788 4120 5840
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 9772 5856 9824 5908
rect 12440 5856 12492 5908
rect 13176 5856 13228 5908
rect 15752 5856 15804 5908
rect 16028 5856 16080 5908
rect 16488 5856 16540 5908
rect 7656 5720 7708 5772
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 10232 5720 10284 5772
rect 14096 5788 14148 5840
rect 15476 5788 15528 5840
rect 15936 5788 15988 5840
rect 18052 5856 18104 5908
rect 17316 5788 17368 5840
rect 19616 5856 19668 5908
rect 20352 5788 20404 5840
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 10968 5720 11020 5772
rect 12440 5720 12492 5772
rect 13912 5763 13964 5772
rect 13912 5729 13921 5763
rect 13921 5729 13955 5763
rect 13955 5729 13964 5763
rect 13912 5720 13964 5729
rect 14556 5720 14608 5772
rect 15200 5720 15252 5772
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 13820 5652 13872 5704
rect 14096 5695 14148 5704
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 12992 5584 13044 5636
rect 13360 5516 13412 5568
rect 13544 5559 13596 5568
rect 13544 5525 13553 5559
rect 13553 5525 13587 5559
rect 13587 5525 13596 5559
rect 13544 5516 13596 5525
rect 19064 5516 19116 5568
rect 20168 5559 20220 5568
rect 20168 5525 20177 5559
rect 20177 5525 20211 5559
rect 20211 5525 20220 5559
rect 20168 5516 20220 5525
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 10784 5312 10836 5364
rect 10876 5244 10928 5296
rect 12624 5312 12676 5364
rect 13820 5355 13872 5364
rect 13820 5321 13829 5355
rect 13829 5321 13863 5355
rect 13863 5321 13872 5355
rect 13820 5312 13872 5321
rect 15200 5312 15252 5364
rect 10600 5176 10652 5228
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 12992 5108 13044 5160
rect 15568 5176 15620 5228
rect 19432 5312 19484 5364
rect 14924 5108 14976 5160
rect 15752 5040 15804 5092
rect 16488 5108 16540 5160
rect 18604 5151 18656 5160
rect 18604 5117 18613 5151
rect 18613 5117 18647 5151
rect 18647 5117 18656 5151
rect 18604 5108 18656 5117
rect 19064 5108 19116 5160
rect 18052 5040 18104 5092
rect 20168 5040 20220 5092
rect 12348 4972 12400 5024
rect 15476 5015 15528 5024
rect 15476 4981 15485 5015
rect 15485 4981 15519 5015
rect 15519 4981 15528 5015
rect 15476 4972 15528 4981
rect 17316 5015 17368 5024
rect 17316 4981 17325 5015
rect 17325 4981 17359 5015
rect 17359 4981 17368 5015
rect 17316 4972 17368 4981
rect 18604 4972 18656 5024
rect 19616 4972 19668 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 13544 4768 13596 4820
rect 16304 4768 16356 4820
rect 18788 4768 18840 4820
rect 19616 4811 19668 4820
rect 19616 4777 19625 4811
rect 19625 4777 19659 4811
rect 19659 4777 19668 4811
rect 19616 4768 19668 4777
rect 20260 4768 20312 4820
rect 9956 4700 10008 4752
rect 16120 4743 16172 4752
rect 12348 4632 12400 4684
rect 16120 4709 16129 4743
rect 16129 4709 16163 4743
rect 16163 4709 16172 4743
rect 16120 4700 16172 4709
rect 12992 4607 13044 4616
rect 12992 4573 13001 4607
rect 13001 4573 13035 4607
rect 13035 4573 13044 4607
rect 12992 4564 13044 4573
rect 12900 4496 12952 4548
rect 14372 4632 14424 4684
rect 15108 4632 15160 4684
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 17316 4564 17368 4616
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 18696 4607 18748 4616
rect 18696 4573 18705 4607
rect 18705 4573 18739 4607
rect 18739 4573 18748 4607
rect 18696 4564 18748 4573
rect 20076 4607 20128 4616
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 20168 4607 20220 4616
rect 20168 4573 20177 4607
rect 20177 4573 20211 4607
rect 20211 4573 20220 4607
rect 20168 4564 20220 4573
rect 16856 4496 16908 4548
rect 19984 4496 20036 4548
rect 11888 4428 11940 4480
rect 14188 4428 14240 4480
rect 14464 4428 14516 4480
rect 16304 4428 16356 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 3056 4088 3108 4140
rect 11152 4224 11204 4276
rect 9956 4088 10008 4140
rect 12348 4156 12400 4208
rect 12808 4156 12860 4208
rect 18696 4224 18748 4276
rect 20076 4224 20128 4276
rect 15476 4156 15528 4208
rect 13912 4088 13964 4140
rect 14556 4131 14608 4140
rect 14556 4097 14565 4131
rect 14565 4097 14599 4131
rect 14599 4097 14608 4131
rect 14556 4088 14608 4097
rect 5816 4020 5868 4072
rect 8760 4020 8812 4072
rect 8944 4063 8996 4072
rect 8944 4029 8953 4063
rect 8953 4029 8987 4063
rect 8987 4029 8996 4063
rect 8944 4020 8996 4029
rect 9220 4063 9272 4072
rect 9220 4029 9254 4063
rect 9254 4029 9272 4063
rect 9220 4020 9272 4029
rect 9680 4020 9732 4072
rect 10508 4020 10560 4072
rect 11796 4063 11848 4072
rect 11796 4029 11827 4063
rect 11827 4029 11848 4063
rect 11796 4020 11848 4029
rect 12716 4063 12768 4072
rect 12716 4029 12725 4063
rect 12725 4029 12759 4063
rect 12759 4029 12768 4063
rect 12716 4020 12768 4029
rect 12992 4063 13044 4072
rect 12992 4029 13001 4063
rect 13001 4029 13035 4063
rect 13035 4029 13044 4063
rect 12992 4020 13044 4029
rect 15752 4063 15804 4072
rect 15752 4029 15761 4063
rect 15761 4029 15795 4063
rect 15795 4029 15804 4063
rect 17960 4156 18012 4208
rect 17224 4088 17276 4140
rect 17868 4088 17920 4140
rect 20352 4156 20404 4208
rect 16304 4063 16356 4072
rect 15752 4020 15804 4029
rect 16304 4029 16313 4063
rect 16313 4029 16347 4063
rect 16347 4029 16356 4063
rect 16304 4020 16356 4029
rect 17408 4063 17460 4072
rect 17408 4029 17417 4063
rect 17417 4029 17451 4063
rect 17451 4029 17460 4063
rect 17408 4020 17460 4029
rect 18052 4063 18104 4072
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 7472 3952 7524 4004
rect 10048 3952 10100 4004
rect 15660 3995 15712 4004
rect 15660 3961 15669 3995
rect 15669 3961 15703 3995
rect 15703 3961 15712 3995
rect 15660 3952 15712 3961
rect 15936 3952 15988 4004
rect 17500 3952 17552 4004
rect 20720 4063 20772 4072
rect 20720 4029 20729 4063
rect 20729 4029 20763 4063
rect 20763 4029 20772 4063
rect 20720 4020 20772 4029
rect 18604 3952 18656 4004
rect 1952 3884 2004 3936
rect 10140 3884 10192 3936
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 11060 3884 11112 3936
rect 12532 3884 12584 3936
rect 13912 3927 13964 3936
rect 13912 3893 13921 3927
rect 13921 3893 13955 3927
rect 13955 3893 13964 3927
rect 13912 3884 13964 3893
rect 14004 3884 14056 3936
rect 15384 3884 15436 3936
rect 17960 3884 18012 3936
rect 20076 3927 20128 3936
rect 20076 3893 20085 3927
rect 20085 3893 20119 3927
rect 20119 3893 20128 3927
rect 20076 3884 20128 3893
rect 21916 3884 21968 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 4160 3680 4212 3732
rect 12348 3680 12400 3732
rect 296 3612 348 3664
rect 9956 3612 10008 3664
rect 10324 3612 10376 3664
rect 10876 3612 10928 3664
rect 14556 3680 14608 3732
rect 13820 3612 13872 3664
rect 5264 3544 5316 3596
rect 9680 3544 9732 3596
rect 8944 3476 8996 3528
rect 12624 3544 12676 3596
rect 15752 3680 15804 3732
rect 18604 3723 18656 3732
rect 16028 3612 16080 3664
rect 18604 3689 18613 3723
rect 18613 3689 18647 3723
rect 18647 3689 18656 3723
rect 18604 3680 18656 3689
rect 17132 3612 17184 3664
rect 15568 3587 15620 3596
rect 15568 3553 15577 3587
rect 15577 3553 15611 3587
rect 15611 3553 15620 3587
rect 15568 3544 15620 3553
rect 18052 3544 18104 3596
rect 18696 3544 18748 3596
rect 19800 3587 19852 3596
rect 19800 3553 19809 3587
rect 19809 3553 19843 3587
rect 19843 3553 19852 3587
rect 19800 3544 19852 3553
rect 19524 3476 19576 3528
rect 20352 3476 20404 3528
rect 11152 3408 11204 3460
rect 12624 3408 12676 3460
rect 3608 3340 3660 3392
rect 13452 3340 13504 3392
rect 13912 3340 13964 3392
rect 19708 3340 19760 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 10692 3179 10744 3188
rect 10692 3145 10701 3179
rect 10701 3145 10735 3179
rect 10735 3145 10744 3179
rect 10692 3136 10744 3145
rect 10784 3136 10836 3188
rect 12440 3136 12492 3188
rect 14004 3136 14056 3188
rect 14188 3136 14240 3188
rect 8300 3068 8352 3120
rect 10048 3068 10100 3120
rect 8576 3000 8628 3052
rect 8300 2864 8352 2916
rect 10048 2864 10100 2916
rect 10784 2932 10836 2984
rect 11060 2975 11112 2984
rect 11060 2941 11069 2975
rect 11069 2941 11103 2975
rect 11103 2941 11112 2975
rect 11060 2932 11112 2941
rect 11336 3043 11388 3052
rect 11336 3009 11345 3043
rect 11345 3009 11379 3043
rect 11379 3009 11388 3043
rect 11336 3000 11388 3009
rect 11520 2932 11572 2984
rect 12348 2932 12400 2984
rect 13268 2932 13320 2984
rect 16028 3068 16080 3120
rect 17040 3136 17092 3188
rect 18512 3136 18564 3188
rect 13912 3043 13964 3052
rect 13912 3009 13921 3043
rect 13921 3009 13955 3043
rect 13955 3009 13964 3043
rect 13912 3000 13964 3009
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 20260 3068 20312 3120
rect 20076 3000 20128 3052
rect 14556 2975 14608 2984
rect 14556 2941 14590 2975
rect 14590 2941 14608 2975
rect 2504 2796 2556 2848
rect 9680 2796 9732 2848
rect 10968 2796 11020 2848
rect 11152 2839 11204 2848
rect 11152 2805 11161 2839
rect 11161 2805 11195 2839
rect 11195 2805 11204 2839
rect 11152 2796 11204 2805
rect 11520 2796 11572 2848
rect 11796 2796 11848 2848
rect 14188 2864 14240 2916
rect 14556 2932 14608 2941
rect 15936 2975 15988 2984
rect 15936 2941 15945 2975
rect 15945 2941 15979 2975
rect 15979 2941 15988 2975
rect 15936 2932 15988 2941
rect 15568 2864 15620 2916
rect 17868 2932 17920 2984
rect 18788 2932 18840 2984
rect 19892 2932 19944 2984
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 18420 2907 18472 2916
rect 18420 2873 18429 2907
rect 18429 2873 18463 2907
rect 18463 2873 18472 2907
rect 18420 2864 18472 2873
rect 16396 2796 16448 2848
rect 16948 2839 17000 2848
rect 16948 2805 16957 2839
rect 16957 2805 16991 2839
rect 16991 2805 17000 2839
rect 21364 2864 21416 2916
rect 16948 2796 17000 2805
rect 22468 2796 22520 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 11152 2592 11204 2644
rect 4712 2456 4764 2508
rect 10968 2456 11020 2508
rect 10876 2431 10928 2440
rect 10876 2397 10885 2431
rect 10885 2397 10919 2431
rect 10919 2397 10928 2431
rect 10876 2388 10928 2397
rect 1400 2320 1452 2372
rect 16212 2592 16264 2644
rect 17684 2592 17736 2644
rect 12440 2524 12492 2576
rect 12072 2456 12124 2508
rect 12256 2456 12308 2508
rect 13360 2499 13412 2508
rect 13360 2465 13369 2499
rect 13369 2465 13403 2499
rect 13403 2465 13412 2499
rect 13360 2456 13412 2465
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 14372 2456 14424 2508
rect 16120 2456 16172 2508
rect 17500 2456 17552 2508
rect 17776 2456 17828 2508
rect 19524 2499 19576 2508
rect 19524 2465 19533 2499
rect 19533 2465 19567 2499
rect 19567 2465 19576 2499
rect 19524 2456 19576 2465
rect 20352 2499 20404 2508
rect 20352 2465 20361 2499
rect 20361 2465 20395 2499
rect 20395 2465 20404 2499
rect 20352 2456 20404 2465
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 16948 2388 17000 2440
rect 13084 2320 13136 2372
rect 15292 2320 15344 2372
rect 13636 2252 13688 2304
rect 15844 2320 15896 2372
rect 18604 2320 18656 2372
rect 16948 2252 17000 2304
rect 17500 2295 17552 2304
rect 17500 2261 17509 2295
rect 17509 2261 17543 2295
rect 17543 2261 17552 2295
rect 17500 2252 17552 2261
rect 19064 2252 19116 2304
rect 19616 2252 19668 2304
rect 20812 2252 20864 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
<< metal2 >>
rect 294 22320 350 22800
rect 846 22320 902 22800
rect 1398 22320 1454 22800
rect 1950 22320 2006 22800
rect 2502 22320 2558 22800
rect 3054 22320 3110 22800
rect 3606 22320 3662 22800
rect 4158 22320 4214 22800
rect 4710 22320 4766 22800
rect 5262 22320 5318 22800
rect 5814 22320 5870 22800
rect 6366 22320 6422 22800
rect 6918 22320 6974 22800
rect 7470 22320 7526 22800
rect 8022 22320 8078 22800
rect 8574 22320 8630 22800
rect 9126 22320 9182 22800
rect 9678 22320 9734 22800
rect 10230 22320 10286 22800
rect 10782 22320 10838 22800
rect 11334 22320 11390 22800
rect 11978 22320 12034 22800
rect 12530 22320 12586 22800
rect 13082 22320 13138 22800
rect 13634 22320 13690 22800
rect 14186 22320 14242 22800
rect 14738 22320 14794 22800
rect 15290 22320 15346 22800
rect 15842 22320 15898 22800
rect 16394 22320 16450 22800
rect 16946 22320 17002 22800
rect 17498 22320 17554 22800
rect 17958 22536 18014 22545
rect 17958 22471 18014 22480
rect 308 18970 336 22320
rect 296 18964 348 18970
rect 296 18906 348 18912
rect 860 17814 888 22320
rect 1412 18766 1440 22320
rect 1964 22250 1992 22320
rect 1504 22222 1992 22250
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1504 18442 1532 22222
rect 2516 19174 2544 22320
rect 2504 19168 2556 19174
rect 2504 19110 2556 19116
rect 1412 18414 1532 18442
rect 848 17808 900 17814
rect 848 17750 900 17756
rect 1412 13297 1440 18414
rect 3068 18358 3096 22320
rect 3056 18352 3108 18358
rect 3056 18294 3108 18300
rect 3620 18154 3648 22320
rect 4172 18222 4200 22320
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4724 18630 4752 22320
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 3608 18148 3660 18154
rect 3608 18090 3660 18096
rect 5276 18034 5304 22320
rect 5276 18006 5580 18034
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 3422 17232 3478 17241
rect 3422 17167 3478 17176
rect 1398 13288 1454 13297
rect 1398 13223 1454 13232
rect 3436 9110 3464 17167
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 5552 14958 5580 18006
rect 5828 16658 5856 22320
rect 6380 19922 6408 22320
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 6196 15026 6224 18566
rect 6932 16726 6960 22320
rect 7484 19990 7512 22320
rect 8036 20346 8064 22320
rect 8036 20318 8248 20346
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7472 19984 7524 19990
rect 7472 19926 7524 19932
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7392 17746 7420 18770
rect 8220 18426 8248 20318
rect 8588 19394 8616 22320
rect 9140 20058 9168 22320
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 8496 19366 8616 19394
rect 8496 19310 8524 19366
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8404 18902 8432 19246
rect 8392 18896 8444 18902
rect 8392 18838 8444 18844
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8680 18290 8708 19654
rect 9232 19242 9260 19790
rect 9220 19236 9272 19242
rect 9220 19178 9272 19184
rect 9232 18970 9260 19178
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 7392 17338 7420 17682
rect 8404 17338 8432 17682
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 7392 16454 7420 17274
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7392 16046 7420 16390
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 6932 15638 6960 15982
rect 6920 15632 6972 15638
rect 6920 15574 6972 15580
rect 7392 15026 7420 15982
rect 7576 15586 7604 16594
rect 7668 16590 7696 17002
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7668 15706 7696 16526
rect 8208 15904 8260 15910
rect 8588 15881 8616 18090
rect 8772 17882 8800 18770
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 8772 17270 8800 17818
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8680 16590 8708 17138
rect 9324 16998 9352 17274
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9048 16794 9076 16934
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8208 15846 8260 15852
rect 8574 15872 8630 15881
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 7576 15558 7696 15586
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 6104 6322 6132 14894
rect 6932 14550 6960 14962
rect 6920 14544 6972 14550
rect 6920 14486 6972 14492
rect 7668 12322 7696 15558
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8128 15162 8156 15506
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8220 14550 8248 15846
rect 8574 15807 8630 15816
rect 9140 15638 9168 16594
rect 9128 15632 9180 15638
rect 9128 15574 9180 15580
rect 8300 14884 8352 14890
rect 8300 14826 8352 14832
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 8312 14346 8340 14826
rect 8588 14618 8616 14826
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 9048 14618 9076 14758
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7576 12294 7696 12322
rect 8496 12306 8524 12786
rect 8484 12300 8536 12306
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7484 11218 7512 12174
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 4068 5840 4120 5846
rect 4066 5808 4068 5817
rect 4120 5808 4122 5817
rect 4066 5743 4122 5752
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 296 3664 348 3670
rect 296 3606 348 3612
rect 308 480 336 3606
rect 846 2952 902 2961
rect 846 2887 902 2896
rect 860 480 888 2887
rect 1400 2372 1452 2378
rect 1400 2314 1452 2320
rect 1412 480 1440 2314
rect 1964 480 1992 3878
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2516 480 2544 2790
rect 3068 480 3096 4082
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3620 480 3648 3334
rect 4172 480 4200 3674
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4724 480 4752 2450
rect 5276 480 5304 3538
rect 5828 480 5856 4014
rect 6366 3496 6422 3505
rect 6366 3431 6422 3440
rect 6380 480 6408 3431
rect 6932 480 6960 8298
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7484 480 7512 3946
rect 7576 3641 7604 12294
rect 8484 12242 8536 12248
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8680 11354 8708 11494
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8576 10532 8628 10538
rect 8576 10474 8628 10480
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7668 9586 7696 9998
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8588 9178 8616 10474
rect 8680 10198 8708 11018
rect 8772 10810 8800 11494
rect 8864 11082 8892 11698
rect 9048 11218 9076 12038
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 9048 10674 9076 11154
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9140 10606 9168 15574
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9232 13938 9260 14214
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9232 12986 9260 13874
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9324 12866 9352 16934
rect 9232 12838 9352 12866
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 6254 7696 6734
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7668 5778 7696 6190
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7760 5914 7788 6122
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 7562 3632 7618 3641
rect 7562 3567 7618 3576
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8220 2530 8248 8842
rect 8588 8634 8616 8910
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8772 4078 8800 9930
rect 8956 5794 8984 10406
rect 9232 9994 9260 12838
rect 9416 12322 9444 19858
rect 9692 19802 9720 22320
rect 10244 19938 10272 22320
rect 10140 19916 10192 19922
rect 10244 19910 10456 19938
rect 10140 19858 10192 19864
rect 9692 19774 9904 19802
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9600 18170 9628 19110
rect 9692 18902 9720 19110
rect 9680 18896 9732 18902
rect 9680 18838 9732 18844
rect 9692 18290 9720 18838
rect 9784 18834 9812 19654
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9600 18142 9720 18170
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9508 16046 9536 16390
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9600 13734 9628 18022
rect 9692 17882 9720 18142
rect 9772 18080 9824 18086
rect 9770 18048 9772 18057
rect 9824 18048 9826 18057
rect 9770 17983 9826 17992
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9876 17105 9904 19774
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9968 18698 9996 19178
rect 10152 18970 10180 19858
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10244 19514 10272 19790
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 10336 19258 10364 19790
rect 10244 19242 10364 19258
rect 10232 19236 10364 19242
rect 10284 19230 10364 19236
rect 10232 19178 10284 19184
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10244 18902 10272 19178
rect 10232 18896 10284 18902
rect 10232 18838 10284 18844
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 10152 18222 10180 18770
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 9956 18080 10008 18086
rect 10048 18080 10100 18086
rect 9956 18022 10008 18028
rect 10046 18048 10048 18057
rect 10100 18048 10102 18057
rect 9968 17746 9996 18022
rect 10046 17983 10102 17992
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9862 17096 9918 17105
rect 9862 17031 9918 17040
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16250 9720 16934
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 15162 9720 15506
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14618 9720 14758
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9324 12294 9444 12322
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9140 9450 9168 9862
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9140 8498 9168 9386
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 8974 9260 9318
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 6934 9168 7278
rect 9128 6928 9180 6934
rect 9128 6870 9180 6876
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9048 6458 9076 6802
rect 9140 6662 9168 6870
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 9140 5914 9168 6122
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 8956 5766 9168 5794
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8956 3534 8984 4014
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8312 2922 8340 3062
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8036 2502 8248 2530
rect 8036 480 8064 2502
rect 8588 480 8616 2994
rect 9140 480 9168 5766
rect 9232 4078 9260 8910
rect 9324 7546 9352 12294
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9416 11218 9444 12106
rect 9508 11694 9536 12174
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9600 8430 9628 13670
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9178 9720 9998
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9416 6730 9444 7210
rect 9692 7002 9720 7890
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5914 9812 6054
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9968 4758 9996 17682
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10152 16726 10180 16934
rect 10140 16720 10192 16726
rect 10140 16662 10192 16668
rect 10046 15600 10102 15609
rect 10046 15535 10048 15544
rect 10100 15535 10102 15544
rect 10048 15506 10100 15512
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10060 13802 10088 14418
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10152 13977 10180 14350
rect 10138 13968 10194 13977
rect 10138 13903 10194 13912
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10152 11898 10180 13330
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10244 11286 10272 18702
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10336 16697 10364 18226
rect 10428 17241 10456 19910
rect 10508 18896 10560 18902
rect 10508 18838 10560 18844
rect 10520 18290 10548 18838
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10414 17232 10470 17241
rect 10414 17167 10470 17176
rect 10322 16688 10378 16697
rect 10322 16623 10378 16632
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10428 16454 10456 16526
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10428 16250 10456 16390
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10520 14278 10548 16594
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10414 13968 10470 13977
rect 10414 13903 10470 13912
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10336 12374 10364 13262
rect 10428 12594 10456 13903
rect 10520 12714 10548 14214
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10612 13326 10640 13670
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10612 12782 10640 13262
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10428 12566 10548 12594
rect 10324 12368 10376 12374
rect 10324 12310 10376 12316
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10152 10577 10180 11222
rect 10138 10568 10194 10577
rect 10138 10503 10194 10512
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10428 9518 10456 9998
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10428 9178 10456 9454
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10428 8430 10456 9114
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10060 6458 10088 6802
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10152 6458 10180 6734
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10232 6384 10284 6390
rect 10152 6332 10232 6338
rect 10152 6326 10284 6332
rect 10152 6310 10272 6326
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 9956 4752 10008 4758
rect 9956 4694 10008 4700
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9692 3602 9720 4014
rect 9968 3670 9996 4082
rect 10060 4010 10088 5714
rect 10152 5710 10180 6310
rect 10232 5772 10284 5778
rect 10336 5760 10364 6802
rect 10284 5732 10364 5760
rect 10232 5714 10284 5720
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10152 3942 10180 5646
rect 10230 4720 10286 4729
rect 10230 4655 10286 4664
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10060 2922 10088 3062
rect 10048 2916 10100 2922
rect 10048 2858 10100 2864
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9692 480 9720 2790
rect 10244 480 10272 4655
rect 10520 4078 10548 12566
rect 10600 11280 10652 11286
rect 10600 11222 10652 11228
rect 10612 10266 10640 11222
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10612 5234 10640 10202
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10336 3670 10364 3878
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10704 3194 10732 18158
rect 10796 18086 10824 22320
rect 11348 20058 11376 22320
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11612 19984 11664 19990
rect 11612 19926 11664 19932
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11440 18902 11468 19110
rect 11428 18896 11480 18902
rect 11428 18838 11480 18844
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 11518 17776 11574 17785
rect 11060 17740 11112 17746
rect 11518 17711 11520 17720
rect 11060 17682 11112 17688
rect 11572 17711 11574 17720
rect 11520 17682 11572 17688
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10888 16726 10916 17614
rect 11072 17082 11100 17682
rect 11624 17610 11652 19926
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11164 17134 11192 17478
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 10980 17054 11100 17082
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 10980 15586 11008 17054
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11072 15706 11100 16934
rect 11256 16538 11284 17138
rect 11164 16510 11284 16538
rect 11164 16454 11192 16510
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 11164 16046 11192 16390
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11518 16144 11574 16153
rect 11624 16114 11652 17206
rect 11518 16079 11574 16088
rect 11612 16108 11664 16114
rect 11532 16046 11560 16079
rect 11612 16050 11664 16056
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 10980 15558 11100 15586
rect 11072 14634 11100 15558
rect 11164 14958 11192 15846
rect 11256 15638 11284 15846
rect 11244 15632 11296 15638
rect 11244 15574 11296 15580
rect 11716 15450 11744 19246
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11808 17082 11836 18566
rect 11900 17202 11928 19654
rect 11992 19174 12020 22320
rect 12544 20058 12572 22320
rect 13096 20058 13124 22320
rect 13268 20732 13320 20738
rect 13268 20674 13320 20680
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11980 18352 12032 18358
rect 11980 18294 12032 18300
rect 11992 17746 12020 18294
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 12268 18034 12296 19858
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12360 19258 12388 19790
rect 12360 19242 12664 19258
rect 12360 19236 12676 19242
rect 12360 19230 12624 19236
rect 12360 18970 12388 19230
rect 12624 19178 12676 19184
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12452 18834 12480 19110
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12544 18193 12572 19110
rect 12912 18902 12940 19110
rect 12900 18896 12952 18902
rect 12900 18838 12952 18844
rect 12900 18420 12952 18426
rect 12900 18362 12952 18368
rect 12530 18184 12586 18193
rect 12530 18119 12586 18128
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11808 17054 11928 17082
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11808 15638 11836 16594
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11900 15502 11928 17054
rect 12084 16538 12112 18022
rect 12268 18006 12388 18034
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 11992 16510 12112 16538
rect 11624 15422 11744 15450
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 11624 14634 11652 15422
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11716 15026 11744 15302
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 10980 14606 11100 14634
rect 11164 14606 11652 14634
rect 10980 13530 11008 14606
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11072 13462 11100 14486
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10796 12850 10824 13126
rect 11072 12986 11100 13194
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10888 12306 10916 12854
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10888 11762 10916 12242
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11072 10792 11100 11154
rect 11164 11121 11192 14606
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11716 14074 11744 14758
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11426 12744 11482 12753
rect 11426 12679 11428 12688
rect 11480 12679 11482 12688
rect 11428 12650 11480 12656
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11150 11112 11206 11121
rect 11440 11098 11468 11494
rect 11624 11234 11652 13466
rect 11808 13462 11836 13874
rect 11992 13530 12020 16510
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12084 16153 12112 16390
rect 12176 16182 12204 16390
rect 12164 16176 12216 16182
rect 12070 16144 12126 16153
rect 12164 16118 12216 16124
rect 12070 16079 12126 16088
rect 12162 16008 12218 16017
rect 12162 15943 12218 15952
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11978 13288 12034 13297
rect 11978 13223 12034 13232
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11808 11694 11836 12038
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11354 11744 11494
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11624 11206 11836 11234
rect 11702 11112 11758 11121
rect 11440 11070 11652 11098
rect 11150 11047 11206 11056
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11072 10764 11284 10792
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10980 9178 11008 10406
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10796 8362 10824 8842
rect 10980 8566 11008 8978
rect 11072 8634 11100 10406
rect 11164 10198 11192 10610
rect 11256 10266 11284 10764
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11164 9654 11192 10134
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11244 9444 11296 9450
rect 11244 9386 11296 9392
rect 11150 9072 11206 9081
rect 11150 9007 11152 9016
rect 11204 9007 11206 9016
rect 11152 8978 11204 8984
rect 11256 8974 11284 9386
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11440 9178 11468 9318
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11244 8968 11296 8974
rect 11164 8916 11244 8922
rect 11164 8910 11296 8916
rect 11164 8894 11284 8910
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10796 7886 10824 8298
rect 10888 7886 10916 8366
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10796 7546 10824 7822
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10980 6866 11008 8502
rect 11164 8430 11192 8894
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11164 8090 11192 8230
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11256 7970 11284 8298
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11164 7942 11284 7970
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10796 5370 10824 6054
rect 10888 5710 10916 6598
rect 10980 6458 11008 6598
rect 11072 6458 11100 7890
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10980 5778 11008 6258
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10888 5302 10916 5646
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10980 5234 11008 5714
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 11164 4282 11192 7942
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11624 7154 11652 11070
rect 11702 11047 11758 11056
rect 11716 8922 11744 11047
rect 11808 10554 11836 11206
rect 11900 10674 11928 12718
rect 11992 10810 12020 13223
rect 12084 12918 12112 14418
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 12176 12782 12204 15943
rect 12164 12776 12216 12782
rect 12070 12744 12126 12753
rect 12164 12718 12216 12724
rect 12070 12679 12126 12688
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11808 10526 11928 10554
rect 11716 8894 11836 8922
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11716 8430 11744 8774
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11808 7750 11836 8894
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11624 7126 11744 7154
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10796 2990 10824 3130
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10782 2816 10838 2825
rect 10782 2751 10838 2760
rect 10796 480 10824 2751
rect 10888 2446 10916 3606
rect 10966 3088 11022 3097
rect 10966 3023 11022 3032
rect 10980 2854 11008 3023
rect 11072 2990 11100 3878
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 3176 11192 3402
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11164 3148 11376 3176
rect 11348 3058 11376 3148
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11532 2854 11560 2926
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11164 2650 11192 2790
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 10980 1601 11008 2450
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11716 1986 11744 7126
rect 11900 4486 11928 10526
rect 12084 9466 12112 12679
rect 12268 12628 12296 17546
rect 12360 16017 12388 18006
rect 12440 17604 12492 17610
rect 12440 17546 12492 17552
rect 12452 17338 12480 17546
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12346 16008 12402 16017
rect 12346 15943 12402 15952
rect 12348 15904 12400 15910
rect 12346 15872 12348 15881
rect 12400 15872 12402 15881
rect 12346 15807 12402 15816
rect 12360 15586 12388 15807
rect 12360 15570 12480 15586
rect 12360 15564 12492 15570
rect 12360 15558 12440 15564
rect 12440 15506 12492 15512
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12360 14550 12388 15438
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12452 14618 12480 14962
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12360 13938 12388 14486
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12544 13394 12572 18119
rect 12912 17270 12940 18362
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12728 15042 12756 16526
rect 12806 16008 12862 16017
rect 12912 15994 12940 16934
rect 12862 15966 12940 15994
rect 12806 15943 12862 15952
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12820 15162 12848 15506
rect 12912 15434 12940 15966
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12728 15014 12848 15042
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12728 14074 12756 14758
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 11992 9438 12112 9466
rect 12176 12600 12296 12628
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11796 4072 11848 4078
rect 11794 4040 11796 4049
rect 11848 4040 11850 4049
rect 11794 3975 11850 3984
rect 11796 2848 11848 2854
rect 11992 2825 12020 9438
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 9042 12112 9318
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12084 8362 12112 8978
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12084 7410 12112 7686
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 6934 12112 7346
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 12072 6384 12124 6390
rect 12176 6361 12204 12600
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12268 11762 12296 12242
rect 12360 11898 12388 13330
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12782 12480 13126
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12636 12442 12664 13262
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12268 11014 12296 11698
rect 12544 11626 12572 12242
rect 12636 11626 12664 12378
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12452 10810 12480 11494
rect 12820 11257 12848 15014
rect 12912 12730 12940 15370
rect 13004 12850 13032 19858
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 13096 17882 13124 18022
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 13188 17338 13216 18022
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13084 15972 13136 15978
rect 13084 15914 13136 15920
rect 13096 15026 13124 15914
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13096 14618 13124 14962
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13188 13530 13216 13874
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 12912 12702 13032 12730
rect 12806 11248 12862 11257
rect 12806 11183 12862 11192
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 10198 12296 10610
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12360 9602 12388 10746
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12636 10470 12664 10678
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12360 9574 12480 9602
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12360 9042 12388 9454
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12072 6326 12124 6332
rect 12162 6352 12218 6361
rect 11796 2790 11848 2796
rect 11978 2816 12034 2825
rect 11348 1958 11744 1986
rect 10966 1592 11022 1601
rect 10966 1527 11022 1536
rect 11348 480 11376 1958
rect 11808 1442 11836 2790
rect 11978 2751 12034 2760
rect 12084 2514 12112 6326
rect 12162 6287 12218 6296
rect 12164 6248 12216 6254
rect 12162 6216 12164 6225
rect 12216 6216 12218 6225
rect 12162 6151 12218 6160
rect 12268 2514 12296 7142
rect 12452 6390 12480 9574
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12544 9110 12572 9454
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12440 6384 12492 6390
rect 12440 6326 12492 6332
rect 12636 6202 12664 10406
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12544 6174 12664 6202
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12360 5953 12388 6054
rect 12346 5944 12402 5953
rect 12452 5914 12480 6054
rect 12346 5879 12402 5888
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12360 4690 12388 4966
rect 12452 4826 12480 5714
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12544 4706 12572 6174
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12452 4678 12572 4706
rect 12348 4208 12400 4214
rect 12348 4150 12400 4156
rect 12360 3738 12388 4150
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12452 3194 12480 4678
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12348 2984 12400 2990
rect 12400 2944 12480 2972
rect 12348 2926 12400 2932
rect 12452 2582 12480 2944
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 11808 1414 12020 1442
rect 11992 480 12020 1414
rect 12544 480 12572 3878
rect 12636 3602 12664 5306
rect 12728 4078 12756 9862
rect 12820 4214 12848 11183
rect 13004 9568 13032 12702
rect 13188 10044 13216 13330
rect 13280 11286 13308 20674
rect 13648 19242 13676 22320
rect 14200 19310 14228 22320
rect 14752 20346 14780 22320
rect 14752 20318 15056 20346
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13556 17678 13584 19110
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13372 17338 13400 17614
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13372 16674 13400 17274
rect 13556 17202 13584 17614
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13452 17060 13504 17066
rect 13452 17002 13504 17008
rect 13464 16794 13492 17002
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13556 16726 13584 16934
rect 13544 16720 13596 16726
rect 13372 16646 13492 16674
rect 13544 16662 13596 16668
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13372 12238 13400 12650
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13268 11280 13320 11286
rect 13268 11222 13320 11228
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13280 10146 13308 10406
rect 13372 10266 13400 11562
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13280 10118 13400 10146
rect 13188 10016 13308 10044
rect 13004 9540 13124 9568
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12912 4554 12940 6054
rect 13004 5642 13032 6258
rect 12992 5636 13044 5642
rect 12992 5578 13044 5584
rect 13004 5166 13032 5578
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 13004 4622 13032 5102
rect 12992 4616 13044 4622
rect 13096 4604 13124 9540
rect 13280 8294 13308 10016
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13188 7342 13216 8230
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13174 5944 13230 5953
rect 13174 5879 13176 5888
rect 13228 5879 13230 5888
rect 13176 5850 13228 5856
rect 13096 4576 13216 4604
rect 12992 4558 13044 4564
rect 12900 4548 12952 4554
rect 12900 4490 12952 4496
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12716 4072 12768 4078
rect 12992 4072 13044 4078
rect 12716 4014 12768 4020
rect 12990 4040 12992 4049
rect 13044 4040 13046 4049
rect 12990 3975 13046 3984
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12636 3097 12664 3402
rect 12622 3088 12678 3097
rect 12622 3023 12678 3032
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 13096 480 13124 2314
rect 13188 1601 13216 4576
rect 13280 2990 13308 7686
rect 13372 6746 13400 10118
rect 13464 6866 13492 16646
rect 13648 16590 13676 18906
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 14016 18222 14044 18566
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 13740 18086 13768 18158
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13740 16046 13768 18022
rect 13924 17746 13952 18090
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13924 16590 13952 17138
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 13912 16584 13964 16590
rect 13912 16526 13964 16532
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13556 15502 13584 15982
rect 13924 15910 13952 16526
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 15706 13952 15846
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 14016 15586 14044 17070
rect 13924 15558 14044 15586
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13556 15026 13584 15438
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13556 14482 13584 14962
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13648 14362 13676 14486
rect 13556 14334 13676 14362
rect 13556 13938 13584 14334
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13648 13870 13676 14214
rect 13740 13870 13768 15302
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13556 11898 13584 13194
rect 13648 12889 13676 13398
rect 13740 13394 13768 13806
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13832 13274 13860 13398
rect 13740 13246 13860 13274
rect 13634 12880 13690 12889
rect 13634 12815 13690 12824
rect 13634 11928 13690 11937
rect 13544 11892 13596 11898
rect 13634 11863 13690 11872
rect 13544 11834 13596 11840
rect 13648 10962 13676 11863
rect 13740 11150 13768 13246
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13832 12850 13860 13126
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13832 11558 13860 12310
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 11218 13860 11494
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13556 10934 13676 10962
rect 13556 10470 13584 10934
rect 13832 10554 13860 11018
rect 13740 10526 13860 10554
rect 13740 10470 13768 10526
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13740 10146 13768 10406
rect 13832 10266 13860 10406
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13740 10118 13860 10146
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13648 9382 13676 9998
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13556 9042 13584 9318
rect 13648 9110 13676 9318
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13648 8022 13676 8434
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13556 7478 13584 7822
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 13648 7410 13676 7958
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13372 6718 13492 6746
rect 13740 6730 13768 8298
rect 13832 7342 13860 10118
rect 13924 9081 13952 15558
rect 14108 13818 14136 19246
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14200 16153 14228 16730
rect 14186 16144 14242 16153
rect 14186 16079 14242 16088
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14200 15706 14228 15982
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14188 13932 14240 13938
rect 14292 13920 14320 19858
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 16726 14412 17478
rect 14476 17134 14504 18770
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14240 13892 14320 13920
rect 14188 13874 14240 13880
rect 14016 13790 14136 13818
rect 14016 13462 14044 13790
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14108 13462 14136 13670
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 14004 13320 14056 13326
rect 14200 13274 14228 13874
rect 14004 13262 14056 13268
rect 14016 11354 14044 13262
rect 14108 13246 14228 13274
rect 14108 11937 14136 13246
rect 14280 12980 14332 12986
rect 14384 12968 14412 14418
rect 14332 12940 14412 12968
rect 14280 12922 14332 12928
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14094 11928 14150 11937
rect 14094 11863 14150 11872
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 13910 9072 13966 9081
rect 13910 9007 13966 9016
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13372 2514 13400 5510
rect 13464 3398 13492 6718
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13556 6186 13584 6394
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 13924 5778 13952 7210
rect 14016 6866 14044 11086
rect 14108 10538 14136 11766
rect 14200 11354 14228 12718
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 14200 9518 14228 11290
rect 14292 10810 14320 11494
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 8566 14136 9318
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 14200 8022 14228 8774
rect 14292 8430 14320 10542
rect 14384 10266 14412 12582
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14384 8362 14412 9930
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14280 8288 14332 8294
rect 14332 8236 14412 8242
rect 14280 8230 14412 8236
rect 14292 8214 14412 8230
rect 14188 8016 14240 8022
rect 14188 7958 14240 7964
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14108 6746 14136 7890
rect 14200 7410 14228 7958
rect 14188 7404 14240 7410
rect 14240 7364 14320 7392
rect 14188 7346 14240 7352
rect 14292 6798 14320 7364
rect 14384 7002 14412 8214
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14476 6866 14504 15846
rect 14568 14550 14596 19246
rect 15028 19174 15056 20318
rect 15304 20058 15332 22320
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 15212 17338 15240 19858
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15304 18426 15332 19178
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15396 18222 15424 18702
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15396 17338 15424 17682
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14740 16720 14792 16726
rect 14738 16688 14740 16697
rect 14792 16688 14794 16697
rect 14738 16623 14794 16632
rect 14752 16289 14780 16623
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 14738 16280 14794 16289
rect 14738 16215 14794 16224
rect 15212 16046 15240 16526
rect 15304 16182 15332 17002
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15396 15892 15424 17138
rect 15212 15864 15424 15892
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14924 15360 14976 15366
rect 14924 15302 14976 15308
rect 14936 15094 14964 15302
rect 14924 15088 14976 15094
rect 14924 15030 14976 15036
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 15028 13938 15056 14758
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14568 13530 14596 13670
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14752 12714 14780 13262
rect 14556 12708 14608 12714
rect 14556 12650 14608 12656
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 14568 12102 14596 12650
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 10062 14596 12038
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 15028 10266 15056 11494
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15120 10198 15148 12174
rect 15212 10742 15240 15864
rect 15488 15026 15516 19246
rect 15580 18970 15608 19246
rect 15856 19174 15884 22320
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 15764 18426 15792 18770
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15580 17338 15608 17614
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15672 16522 15700 17614
rect 15764 17202 15792 18362
rect 15936 18148 15988 18154
rect 15936 18090 15988 18096
rect 15948 17202 15976 18090
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 15948 16590 15976 17138
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15658 16416 15714 16425
rect 15658 16351 15714 16360
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 15638 15608 15846
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15580 15502 15608 15574
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15304 14618 15332 14894
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15580 14414 15608 15438
rect 15672 14906 15700 16351
rect 15936 16176 15988 16182
rect 15750 16144 15806 16153
rect 15936 16118 15988 16124
rect 15750 16079 15806 16088
rect 15764 15638 15792 16079
rect 15948 15910 15976 16118
rect 15844 15904 15896 15910
rect 15936 15904 15988 15910
rect 15844 15846 15896 15852
rect 15934 15872 15936 15881
rect 15988 15872 15990 15881
rect 15752 15632 15804 15638
rect 15752 15574 15804 15580
rect 15672 14878 15792 14906
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15672 14618 15700 14758
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15764 14226 15792 14878
rect 15856 14618 15884 15846
rect 15934 15807 15990 15816
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15396 14198 15792 14226
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15304 11626 15332 13670
rect 15396 11937 15424 14198
rect 15752 14000 15804 14006
rect 15658 13968 15714 13977
rect 15568 13932 15620 13938
rect 15752 13942 15804 13948
rect 15658 13903 15714 13912
rect 15568 13874 15620 13880
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15382 11928 15438 11937
rect 15382 11863 15438 11872
rect 15488 11778 15516 13738
rect 15396 11750 15516 11778
rect 15580 11762 15608 13874
rect 15672 13802 15700 13903
rect 15660 13796 15712 13802
rect 15660 13738 15712 13744
rect 15568 11756 15620 11762
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 15108 10192 15160 10198
rect 14738 10160 14794 10169
rect 15108 10134 15160 10140
rect 14738 10095 14794 10104
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14648 9512 14700 9518
rect 14568 9472 14648 9500
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14016 6718 14136 6746
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14016 6118 14044 6718
rect 14096 6656 14148 6662
rect 14476 6610 14504 6802
rect 14096 6598 14148 6604
rect 14108 6322 14136 6598
rect 14292 6582 14504 6610
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14108 5846 14136 6258
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13556 4826 13584 5510
rect 13832 5370 13860 5646
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13924 4146 13952 5714
rect 14108 5710 14136 5782
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14108 4622 14136 5646
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13832 3210 13860 3606
rect 13924 3398 13952 3878
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13832 3182 13952 3210
rect 14016 3194 14044 3878
rect 14200 3194 14228 4422
rect 13924 3058 13952 3182
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13174 1592 13230 1601
rect 13174 1527 13230 1536
rect 13648 480 13676 2246
rect 14200 480 14228 2858
rect 14292 2514 14320 6582
rect 14568 5778 14596 9472
rect 14752 9500 14780 10095
rect 15106 10024 15162 10033
rect 15106 9959 15162 9968
rect 14700 9472 14780 9500
rect 14648 9454 14700 9460
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 15120 8838 15148 9959
rect 15212 9178 15240 10474
rect 15304 10010 15332 10610
rect 15396 10146 15424 11750
rect 15568 11698 15620 11704
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15488 10266 15516 11562
rect 15580 11218 15608 11698
rect 15672 11354 15700 13738
rect 15764 13462 15792 13942
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15752 13456 15804 13462
rect 15752 13398 15804 13404
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15764 12850 15792 13126
rect 15856 12986 15884 13806
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15764 12374 15792 12582
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15752 12232 15804 12238
rect 15856 12220 15884 12582
rect 15804 12192 15884 12220
rect 15752 12174 15804 12180
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15750 11792 15806 11801
rect 15750 11727 15806 11736
rect 15764 11558 15792 11727
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15580 10606 15608 10950
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15658 10568 15714 10577
rect 15658 10503 15714 10512
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15396 10118 15516 10146
rect 15304 9994 15424 10010
rect 15304 9988 15436 9994
rect 15304 9982 15384 9988
rect 15304 9722 15332 9982
rect 15384 9930 15436 9936
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15304 9518 15332 9658
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15488 9178 15516 10118
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15580 8906 15608 9318
rect 15672 8974 15700 10503
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 14752 8498 14780 8774
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14924 5160 14976 5166
rect 15028 5148 15056 8298
rect 14976 5120 15056 5148
rect 14924 5102 14976 5108
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 15120 4690 15148 8774
rect 15580 8498 15608 8842
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15672 8378 15700 8910
rect 15764 8514 15792 11494
rect 15856 11082 15884 11834
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 15856 8974 15884 9386
rect 15948 9042 15976 14962
rect 16040 9518 16068 19858
rect 16408 19174 16436 22320
rect 16960 20058 16988 22320
rect 17512 20058 17540 22320
rect 17972 20738 18000 22471
rect 18050 22320 18106 22800
rect 18602 22320 18658 22800
rect 19154 22320 19210 22800
rect 19706 22320 19762 22800
rect 20258 22320 20314 22800
rect 20810 22320 20866 22800
rect 21362 22320 21418 22800
rect 21914 22320 21970 22800
rect 22466 22320 22522 22800
rect 17960 20732 18012 20738
rect 17960 20674 18012 20680
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 16132 18086 16160 18770
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 16132 17678 16160 18022
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16120 17264 16172 17270
rect 16120 17206 16172 17212
rect 16132 16726 16160 17206
rect 16316 16998 16344 18090
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16120 16720 16172 16726
rect 16118 16688 16120 16697
rect 16172 16688 16174 16697
rect 16118 16623 16174 16632
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16132 15026 16160 16050
rect 16316 16046 16344 16934
rect 16500 16833 16528 19790
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16486 16824 16542 16833
rect 16486 16759 16542 16768
rect 16592 16658 16620 16934
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16500 16250 16528 16390
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16304 16040 16356 16046
rect 16224 16000 16304 16028
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 16224 14906 16252 16000
rect 16580 16040 16632 16046
rect 16304 15982 16356 15988
rect 16486 16008 16542 16017
rect 16580 15982 16632 15988
rect 16486 15943 16542 15952
rect 16500 15910 16528 15943
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16132 14878 16252 14906
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8634 15884 8910
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15764 8486 15884 8514
rect 15304 8294 15332 8366
rect 15672 8350 15792 8378
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15658 7440 15714 7449
rect 15212 6730 15240 7414
rect 15658 7375 15714 7384
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 15212 5778 15240 6666
rect 15304 6458 15332 6734
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15212 5370 15240 5714
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15304 4865 15332 6122
rect 15290 4856 15346 4865
rect 15290 4791 15346 4800
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 14384 2514 14412 4626
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14476 1442 14504 4422
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14568 3738 14596 4082
rect 15396 3942 15424 6870
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15488 5846 15516 6258
rect 15672 6254 15700 7375
rect 15764 6254 15792 8350
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15488 5030 15516 5782
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15488 4214 15516 4966
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14568 2990 14596 3674
rect 15580 3602 15608 5170
rect 15672 4010 15700 6190
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15764 5914 15792 6054
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15752 5092 15804 5098
rect 15752 5034 15804 5040
rect 15764 4078 15792 5034
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15856 3890 15884 8486
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16132 6746 16160 14878
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16224 13852 16252 14350
rect 16500 14074 16528 15506
rect 16592 15502 16620 15982
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16304 13864 16356 13870
rect 16224 13824 16304 13852
rect 16224 12918 16252 13824
rect 16304 13806 16356 13812
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16224 12646 16252 12854
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16316 11914 16344 13126
rect 16408 12889 16436 13330
rect 16394 12880 16450 12889
rect 16394 12815 16450 12824
rect 16500 12782 16528 14010
rect 16684 13802 16712 19858
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16672 13796 16724 13802
rect 16672 13738 16724 13744
rect 16776 13682 16804 19246
rect 16868 17610 16896 19858
rect 18064 19700 18092 22320
rect 18510 22128 18566 22137
rect 18510 22063 18566 22072
rect 18524 20058 18552 22063
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18616 19786 18644 22320
rect 19062 21584 19118 21593
rect 19062 21519 19118 21528
rect 18694 21176 18750 21185
rect 18694 21111 18750 21120
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 17972 19672 18092 19700
rect 18512 19712 18564 19718
rect 17776 19508 17828 19514
rect 17776 19450 17828 19456
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16960 17202 16988 17614
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 16856 16176 16908 16182
rect 16856 16118 16908 16124
rect 16868 15706 16896 16118
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16868 15026 16896 15302
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16960 14074 16988 16594
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16684 13654 16804 13682
rect 16684 13410 16712 13654
rect 16580 13388 16632 13394
rect 16684 13382 16804 13410
rect 16580 13330 16632 13336
rect 16592 12986 16620 13330
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16316 11886 16436 11914
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 11257 16252 11494
rect 16302 11384 16358 11393
rect 16302 11319 16358 11328
rect 16210 11248 16266 11257
rect 16210 11183 16266 11192
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 16224 9654 16252 10474
rect 16316 10169 16344 11319
rect 16302 10160 16358 10169
rect 16302 10095 16358 10104
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 16316 7886 16344 8298
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16316 7546 16344 7822
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16304 6792 16356 6798
rect 15948 6322 15976 6734
rect 16132 6718 16252 6746
rect 16304 6734 16356 6740
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 16028 6248 16080 6254
rect 15948 6196 16028 6202
rect 15948 6190 16080 6196
rect 15948 6174 16068 6190
rect 15948 5846 15976 6174
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 16040 4570 16068 5850
rect 16132 4758 16160 6598
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 16040 4542 16160 4570
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15764 3862 15884 3890
rect 15764 3738 15792 3862
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 15580 2922 15608 3538
rect 15948 2990 15976 3946
rect 16028 3664 16080 3670
rect 16028 3606 16080 3612
rect 16040 3126 16068 3606
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 15568 2916 15620 2922
rect 15568 2858 15620 2864
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 16040 2446 16068 3062
rect 16132 2514 16160 4542
rect 16224 2650 16252 6718
rect 16316 6254 16344 6734
rect 16408 6458 16436 11886
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16592 10606 16620 11290
rect 16684 10713 16712 13194
rect 16670 10704 16726 10713
rect 16670 10639 16726 10648
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16672 10532 16724 10538
rect 16672 10474 16724 10480
rect 16578 10432 16634 10441
rect 16578 10367 16634 10376
rect 16488 9444 16540 9450
rect 16488 9386 16540 9392
rect 16500 8838 16528 9386
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16592 8650 16620 10367
rect 16684 8906 16712 10474
rect 16776 10198 16804 13382
rect 16868 13326 16896 13806
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16960 12442 16988 14010
rect 17052 13530 17080 16594
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17144 12186 17172 19246
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17236 18290 17264 18566
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17236 17746 17264 18226
rect 17788 18222 17816 19450
rect 17972 18850 18000 19672
rect 18512 19654 18564 19660
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18524 19242 18552 19654
rect 18512 19236 18564 19242
rect 18512 19178 18564 19184
rect 18708 19174 18736 21111
rect 18970 20224 19026 20233
rect 18970 20159 19026 20168
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18800 19394 18828 19858
rect 18984 19514 19012 20159
rect 19076 20058 19104 21519
rect 19168 20058 19196 22320
rect 19246 20632 19302 20641
rect 19246 20567 19302 20576
rect 19260 20058 19288 20567
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19062 19816 19118 19825
rect 19062 19751 19118 19760
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18800 19366 19012 19394
rect 18786 19272 18842 19281
rect 18786 19207 18842 19216
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 17880 18822 18000 18850
rect 18604 18828 18656 18834
rect 17880 18426 17908 18822
rect 18604 18770 18656 18776
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 17972 18426 18000 18702
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17776 18216 17828 18222
rect 17776 18158 17828 18164
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 17420 18057 17448 18158
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17406 18048 17462 18057
rect 17406 17983 17462 17992
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17774 17232 17830 17241
rect 17774 17167 17830 17176
rect 17316 17128 17368 17134
rect 17316 17070 17368 17076
rect 17682 17096 17738 17105
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17236 13258 17264 16934
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17328 12753 17356 17070
rect 17682 17031 17738 17040
rect 17592 16516 17644 16522
rect 17592 16458 17644 16464
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17408 15972 17460 15978
rect 17408 15914 17460 15920
rect 17420 14770 17448 15914
rect 17512 15706 17540 16050
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17604 15609 17632 16458
rect 17696 15978 17724 17031
rect 17684 15972 17736 15978
rect 17684 15914 17736 15920
rect 17590 15600 17646 15609
rect 17590 15535 17646 15544
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17420 14742 17540 14770
rect 17314 12744 17370 12753
rect 17314 12679 17370 12688
rect 17052 12158 17172 12186
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16868 10130 16896 11494
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16960 10538 16988 10950
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16854 10024 16910 10033
rect 16854 9959 16910 9968
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16500 8622 16620 8650
rect 16500 7154 16528 8622
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16592 7274 16620 8434
rect 16684 7886 16712 8842
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16670 7712 16726 7721
rect 16670 7647 16726 7656
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16500 7126 16620 7154
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16408 6186 16436 6394
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16396 6180 16448 6186
rect 16396 6122 16448 6128
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 16316 4826 16344 6054
rect 16500 5914 16528 6258
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16500 5166 16528 5850
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16316 4078 16344 4422
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16592 3505 16620 7126
rect 16684 6225 16712 7647
rect 16776 7546 16804 7890
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16670 6216 16726 6225
rect 16670 6151 16726 6160
rect 16684 6118 16712 6151
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16868 4554 16896 9959
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16960 8430 16988 8978
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16960 6866 16988 8366
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16578 3496 16634 3505
rect 16578 3431 16634 3440
rect 17052 3194 17080 12158
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17144 11234 17172 12038
rect 17236 11694 17264 12038
rect 17328 11778 17356 12679
rect 17328 11750 17448 11778
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17144 11218 17264 11234
rect 17144 11212 17276 11218
rect 17144 11206 17224 11212
rect 17224 11154 17276 11160
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 17144 10266 17172 10474
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17144 4729 17172 9658
rect 17236 9586 17264 11154
rect 17328 10810 17356 11494
rect 17420 11218 17448 11750
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17406 11112 17462 11121
rect 17406 11047 17462 11056
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17314 10704 17370 10713
rect 17314 10639 17370 10648
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17236 7342 17264 8230
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17328 5930 17356 10639
rect 17420 9382 17448 11047
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17512 7562 17540 14742
rect 17696 14618 17724 15506
rect 17788 15026 17816 17167
rect 17972 17134 18000 18090
rect 18064 17882 18092 18158
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18156 17678 18184 18294
rect 18524 17898 18552 18702
rect 18432 17882 18552 17898
rect 18616 17882 18644 18770
rect 18694 18184 18750 18193
rect 18694 18119 18750 18128
rect 18708 18086 18736 18119
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18420 17876 18552 17882
rect 18472 17870 18552 17876
rect 18420 17818 18472 17824
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 17960 16992 18012 16998
rect 17958 16960 17960 16969
rect 18012 16960 18014 16969
rect 17958 16895 18014 16904
rect 18064 16436 18092 17070
rect 18524 17066 18552 17870
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18616 17134 18644 17546
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18512 17060 18564 17066
rect 18512 17002 18564 17008
rect 18144 16992 18196 16998
rect 18708 16980 18736 17070
rect 18616 16952 18736 16980
rect 18616 16946 18644 16952
rect 18144 16934 18196 16940
rect 18156 16794 18184 16934
rect 18524 16918 18644 16946
rect 18524 16794 18552 16918
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 17972 16408 18092 16436
rect 17972 16028 18000 16408
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18052 16040 18104 16046
rect 17972 16000 18052 16028
rect 18052 15982 18104 15988
rect 18064 15570 18092 15982
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17684 14612 17736 14618
rect 17684 14554 17736 14560
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17604 14074 17632 14418
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17604 13394 17632 14010
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17604 12850 17632 13330
rect 17696 13326 17724 14554
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17788 13190 17816 14962
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 17972 12782 18000 14350
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18064 13530 18092 13670
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 18432 13258 18460 13670
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18524 12968 18552 16594
rect 18800 13954 18828 19207
rect 18880 18828 18932 18834
rect 18880 18770 18932 18776
rect 18616 13926 18828 13954
rect 18616 12986 18644 13926
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18432 12940 18552 12968
rect 18604 12980 18656 12986
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 17592 12708 17644 12714
rect 17592 12650 17644 12656
rect 17604 10266 17632 12650
rect 17868 12436 17920 12442
rect 17788 12396 17868 12424
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17696 10470 17724 11698
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17604 8956 17632 9318
rect 17696 9110 17724 10406
rect 17788 9722 17816 12396
rect 17868 12378 17920 12384
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17880 11354 17908 12038
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17972 10674 18000 12310
rect 18156 12306 18184 12718
rect 18432 12374 18460 12940
rect 18604 12922 18656 12928
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18616 12238 18644 12786
rect 18604 12232 18656 12238
rect 18510 12200 18566 12209
rect 18604 12174 18656 12180
rect 18510 12135 18566 12144
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18236 11824 18288 11830
rect 18234 11792 18236 11801
rect 18288 11792 18290 11801
rect 18234 11727 18290 11736
rect 18524 11626 18552 12135
rect 18616 11830 18644 12174
rect 18604 11824 18656 11830
rect 18604 11766 18656 11772
rect 18708 11762 18736 13670
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18604 11552 18656 11558
rect 18524 11500 18604 11506
rect 18524 11494 18656 11500
rect 18524 11478 18644 11494
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17868 10600 17920 10606
rect 17920 10548 18000 10554
rect 17868 10542 18000 10548
rect 17880 10526 18000 10542
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17972 9654 18000 10526
rect 18524 10441 18552 11478
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 18616 11150 18644 11222
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18510 10432 18566 10441
rect 18510 10367 18566 10376
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18420 10056 18472 10062
rect 18418 10024 18420 10033
rect 18472 10024 18474 10033
rect 18418 9959 18474 9968
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18524 9722 18552 10066
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 17958 9208 18014 9217
rect 17958 9143 17960 9152
rect 18012 9143 18014 9152
rect 17960 9114 18012 9120
rect 17684 9104 17736 9110
rect 17684 9046 17736 9052
rect 18340 8974 18368 9590
rect 18418 9480 18474 9489
rect 18418 9415 18420 9424
rect 18472 9415 18474 9424
rect 18420 9386 18472 9392
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18328 8968 18380 8974
rect 17604 8928 17724 8956
rect 17512 7534 17632 7562
rect 17408 7472 17460 7478
rect 17408 7414 17460 7420
rect 17236 5902 17356 5930
rect 17130 4720 17186 4729
rect 17130 4655 17186 4664
rect 17236 4146 17264 5902
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 17328 5030 17356 5782
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 17328 4622 17356 4966
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17420 4078 17448 7414
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 17500 4004 17552 4010
rect 17500 3946 17552 3952
rect 17132 3664 17184 3670
rect 17512 3641 17540 3946
rect 17132 3606 17184 3612
rect 17498 3632 17554 3641
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 17144 3058 17172 3606
rect 17498 3567 17554 3576
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16224 2553 16252 2586
rect 16210 2544 16266 2553
rect 16120 2508 16172 2514
rect 16210 2479 16266 2488
rect 16120 2450 16172 2456
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 15292 2372 15344 2378
rect 15292 2314 15344 2320
rect 15844 2372 15896 2378
rect 15844 2314 15896 2320
rect 14476 1414 14780 1442
rect 14752 480 14780 1414
rect 15304 480 15332 2314
rect 15856 480 15884 2314
rect 16408 480 16436 2790
rect 16960 2446 16988 2790
rect 17512 2514 17540 3567
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 16960 480 16988 2246
rect 17512 480 17540 2246
rect 17604 649 17632 7534
rect 17696 2650 17724 8928
rect 17958 8936 18014 8945
rect 18328 8910 18380 8916
rect 17958 8871 18014 8880
rect 17776 8832 17828 8838
rect 17972 8820 18000 8871
rect 17776 8774 17828 8780
rect 17880 8792 18000 8820
rect 17788 7954 17816 8774
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17880 7857 17908 8792
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18142 8528 18198 8537
rect 18142 8463 18198 8472
rect 18156 8362 18184 8463
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17866 7848 17922 7857
rect 17866 7783 17922 7792
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17788 7546 17816 7686
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17880 7410 17908 7686
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17972 7342 18000 8230
rect 18050 8120 18106 8129
rect 18050 8055 18052 8064
rect 18104 8055 18106 8064
rect 18052 8026 18104 8032
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18524 7342 18552 9318
rect 18616 8634 18644 11086
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18616 8022 18644 8434
rect 18604 8016 18656 8022
rect 18604 7958 18656 7964
rect 18616 7392 18644 7958
rect 18708 7562 18736 11562
rect 18800 11370 18828 13738
rect 18892 11626 18920 18770
rect 18984 18290 19012 19366
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 19076 18170 19104 19751
rect 19168 18902 19196 19858
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19156 18896 19208 18902
rect 19260 18873 19288 19110
rect 19156 18838 19208 18844
rect 19246 18864 19302 18873
rect 19246 18799 19302 18808
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 18984 18142 19104 18170
rect 18984 13734 19012 18142
rect 19064 18080 19116 18086
rect 19064 18022 19116 18028
rect 19076 16561 19104 18022
rect 19168 16776 19196 18226
rect 19260 17746 19288 18566
rect 19352 17785 19380 19246
rect 19444 18902 19472 19858
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19338 17776 19394 17785
rect 19248 17740 19300 17746
rect 19338 17711 19394 17720
rect 19248 17682 19300 17688
rect 19168 16748 19288 16776
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 19062 16552 19118 16561
rect 19062 16487 19118 16496
rect 19168 16182 19196 16594
rect 19156 16176 19208 16182
rect 19156 16118 19208 16124
rect 19156 15904 19208 15910
rect 19260 15881 19288 16748
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19444 16250 19472 16526
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19156 15846 19208 15852
rect 19246 15872 19302 15881
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18984 12866 19012 13330
rect 19076 13258 19104 13806
rect 19064 13252 19116 13258
rect 19064 13194 19116 13200
rect 19076 12986 19104 13194
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19168 12889 19196 15846
rect 19246 15807 19302 15816
rect 19260 14822 19288 15807
rect 19444 15638 19472 16186
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19260 13410 19288 14758
rect 19260 13382 19380 13410
rect 19248 13320 19300 13326
rect 19246 13288 19248 13297
rect 19300 13288 19302 13297
rect 19246 13223 19302 13232
rect 19246 13152 19302 13161
rect 19352 13138 19380 13382
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19302 13110 19380 13138
rect 19246 13087 19302 13096
rect 19154 12880 19210 12889
rect 18984 12838 19104 12866
rect 19076 12764 19104 12838
rect 19154 12815 19210 12824
rect 18970 12744 19026 12753
rect 19076 12736 19196 12764
rect 18970 12679 19026 12688
rect 18880 11620 18932 11626
rect 18880 11562 18932 11568
rect 18800 11342 18920 11370
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18800 10606 18828 10950
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18788 10192 18840 10198
rect 18788 10134 18840 10140
rect 18800 10062 18828 10134
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18800 7750 18828 9658
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18708 7534 18828 7562
rect 18696 7404 18748 7410
rect 18616 7364 18696 7392
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18524 6458 18552 7142
rect 18616 7002 18644 7364
rect 18696 7346 18748 7352
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 17774 6352 17830 6361
rect 17774 6287 17830 6296
rect 18418 6352 18474 6361
rect 18616 6322 18644 6938
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18418 6287 18474 6296
rect 18604 6316 18656 6322
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17788 2514 17816 6287
rect 18432 6254 18460 6287
rect 18604 6258 18656 6264
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18064 5817 18092 5850
rect 18050 5808 18106 5817
rect 18050 5743 18106 5752
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 18050 5264 18106 5273
rect 18050 5199 18106 5208
rect 18064 5098 18092 5199
rect 18616 5166 18644 6054
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18052 5092 18104 5098
rect 18052 5034 18104 5040
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 17960 4208 18012 4214
rect 17958 4176 17960 4185
rect 18012 4176 18014 4185
rect 17868 4140 17920 4146
rect 17958 4111 18014 4120
rect 17868 4082 17920 4088
rect 17880 2990 17908 4082
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 17880 2009 17908 2926
rect 17866 2000 17922 2009
rect 17866 1935 17922 1944
rect 17972 1034 18000 3878
rect 18064 3602 18092 4014
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18524 3194 18552 4558
rect 18616 4162 18644 4966
rect 18708 4622 18736 6802
rect 18800 4826 18828 7534
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18708 4282 18736 4558
rect 18696 4276 18748 4282
rect 18696 4218 18748 4224
rect 18616 4134 18736 4162
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 18616 3738 18644 3946
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18616 3058 18644 3674
rect 18708 3602 18736 4134
rect 18786 4040 18842 4049
rect 18786 3975 18842 3984
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18800 2990 18828 3975
rect 18788 2984 18840 2990
rect 18418 2952 18474 2961
rect 18418 2887 18420 2896
rect 18472 2887 18474 2896
rect 18786 2952 18788 2961
rect 18840 2952 18842 2961
rect 18786 2887 18842 2896
rect 18420 2858 18472 2864
rect 18604 2372 18656 2378
rect 18604 2314 18656 2320
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1006 18092 1034
rect 17590 640 17646 649
rect 17590 575 17646 584
rect 18064 480 18092 1006
rect 18616 480 18644 2314
rect 18892 1057 18920 11342
rect 18984 11150 19012 12679
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18984 9518 19012 10406
rect 19076 9994 19104 11018
rect 19064 9988 19116 9994
rect 19064 9930 19116 9936
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18970 9072 19026 9081
rect 18970 9007 19026 9016
rect 18984 6186 19012 9007
rect 19076 8838 19104 9930
rect 19168 9738 19196 12736
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19260 11762 19288 12242
rect 19444 11898 19472 13330
rect 19536 12458 19564 18770
rect 19720 18698 19748 22320
rect 20272 20210 20300 22320
rect 20088 20182 20300 20210
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19812 17542 19840 18158
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19706 16824 19762 16833
rect 19706 16759 19762 16768
rect 19720 16590 19748 16759
rect 19812 16590 19840 16934
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19812 16046 19840 16526
rect 19904 16114 19932 18158
rect 19996 17202 20024 19246
rect 20088 18970 20116 20182
rect 20824 19938 20852 22320
rect 20536 19916 20588 19922
rect 20824 19910 21036 19938
rect 20536 19858 20588 19864
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 20180 17921 20208 19110
rect 20272 18329 20300 19654
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20258 18320 20314 18329
rect 20258 18255 20314 18264
rect 20166 17912 20222 17921
rect 20166 17847 20222 17856
rect 20364 17338 20392 19246
rect 20548 17814 20576 19858
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20536 17808 20588 17814
rect 20536 17750 20588 17756
rect 20640 17377 20668 19654
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20626 17368 20682 17377
rect 20352 17332 20404 17338
rect 20626 17303 20682 17312
rect 20352 17274 20404 17280
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19800 16040 19852 16046
rect 19800 15982 19852 15988
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19812 15026 19840 15302
rect 20088 15162 20116 15506
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19720 14074 19748 14758
rect 19812 14550 19840 14962
rect 19800 14544 19852 14550
rect 19800 14486 19852 14492
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19812 13938 19840 14486
rect 19996 14278 20024 14962
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 20088 13802 20116 14350
rect 20076 13796 20128 13802
rect 20076 13738 20128 13744
rect 20180 13530 20208 14894
rect 20272 14482 20300 15438
rect 20456 15065 20484 16390
rect 20548 15094 20576 17070
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20536 15088 20588 15094
rect 20442 15056 20498 15065
rect 20536 15030 20588 15036
rect 20442 14991 20498 15000
rect 20640 14657 20668 15846
rect 20732 15609 20760 18022
rect 20824 16017 20852 19110
rect 20916 17202 20944 19790
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 21008 17066 21036 19910
rect 21376 19242 21404 22320
rect 21364 19236 21416 19242
rect 21364 19178 21416 19184
rect 20996 17060 21048 17066
rect 20996 17002 21048 17008
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20904 16040 20956 16046
rect 20810 16008 20866 16017
rect 20904 15982 20956 15988
rect 20810 15943 20866 15952
rect 20718 15600 20774 15609
rect 20718 15535 20774 15544
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20626 14648 20682 14657
rect 20626 14583 20682 14592
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20456 13705 20484 14214
rect 20732 13870 20760 15370
rect 20916 14890 20944 15982
rect 21008 15026 21036 16730
rect 21928 16658 21956 22320
rect 22480 17610 22508 22320
rect 22468 17604 22520 17610
rect 22468 17546 22520 17552
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 20904 14884 20956 14890
rect 20904 14826 20956 14832
rect 20902 14104 20958 14113
rect 20902 14039 20904 14048
rect 20956 14039 20958 14048
rect 20904 14010 20956 14016
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20442 13696 20498 13705
rect 20442 13631 20498 13640
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20442 13288 20498 13297
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19536 12430 19748 12458
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19260 11558 19288 11698
rect 19628 11694 19656 12174
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 19248 11552 19300 11558
rect 19720 11506 19748 12430
rect 19248 11494 19300 11500
rect 19260 11370 19288 11494
rect 19628 11478 19748 11506
rect 19260 11342 19380 11370
rect 19352 11286 19380 11342
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 19159 9710 19196 9738
rect 19159 9353 19187 9710
rect 19154 9344 19210 9353
rect 19154 9279 19210 9288
rect 19260 9178 19288 11222
rect 19522 10840 19578 10849
rect 19522 10775 19578 10784
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19352 9926 19380 10542
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19352 9722 19380 9862
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19430 9480 19486 9489
rect 19430 9415 19486 9424
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19246 9072 19302 9081
rect 19246 9007 19302 9016
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 19076 7177 19104 7686
rect 19260 7290 19288 9007
rect 19444 7342 19472 9415
rect 19536 8945 19564 10775
rect 19522 8936 19578 8945
rect 19522 8871 19578 8880
rect 19432 7336 19484 7342
rect 19260 7262 19380 7290
rect 19432 7278 19484 7284
rect 19248 7200 19300 7206
rect 19062 7168 19118 7177
rect 19248 7142 19300 7148
rect 19062 7103 19118 7112
rect 19076 6254 19104 7103
rect 19064 6248 19116 6254
rect 19260 6225 19288 7142
rect 19064 6190 19116 6196
rect 19246 6216 19302 6225
rect 18972 6180 19024 6186
rect 19246 6151 19302 6160
rect 18972 6122 19024 6128
rect 18984 3913 19012 6122
rect 19352 6100 19380 7262
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19260 6072 19380 6100
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 19076 5166 19104 5510
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 18970 3904 19026 3913
rect 18970 3839 19026 3848
rect 19260 3505 19288 6072
rect 19444 5370 19472 6802
rect 19628 6202 19656 11478
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19720 10441 19748 11154
rect 19706 10432 19762 10441
rect 19706 10367 19762 10376
rect 19720 6322 19748 10367
rect 19812 9110 19840 12786
rect 19996 12782 20024 13194
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 19996 12442 20024 12718
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 19996 10198 20024 11562
rect 20272 11354 20300 13262
rect 20442 13223 20498 13232
rect 20456 12442 20484 13223
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20272 10266 20300 11086
rect 20548 10690 20576 12582
rect 20456 10662 20576 10690
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 19984 10192 20036 10198
rect 19984 10134 20036 10140
rect 20456 10033 20484 10662
rect 20640 10554 20668 12650
rect 20536 10532 20588 10538
rect 20640 10526 20760 10554
rect 20536 10474 20588 10480
rect 20548 10266 20576 10474
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20640 10198 20668 10406
rect 20628 10192 20680 10198
rect 20628 10134 20680 10140
rect 20442 10024 20498 10033
rect 20732 10010 20760 10526
rect 20442 9959 20498 9968
rect 20640 9982 20760 10010
rect 20456 9586 20484 9959
rect 20640 9738 20668 9982
rect 20548 9710 20668 9738
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 19800 9104 19852 9110
rect 19800 9046 19852 9052
rect 19800 8560 19852 8566
rect 19800 8502 19852 8508
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19628 6174 19748 6202
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19628 5914 19656 6054
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19616 5024 19668 5030
rect 19616 4966 19668 4972
rect 19628 4826 19656 4966
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19524 3528 19576 3534
rect 19246 3496 19302 3505
rect 19524 3470 19576 3476
rect 19246 3431 19302 3440
rect 19536 2514 19564 3470
rect 19720 3398 19748 6174
rect 19812 3602 19840 8502
rect 19904 8430 19932 9318
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 20088 8498 20116 8978
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19996 7546 20024 8230
rect 20088 8090 20116 8434
rect 20364 8090 20392 9318
rect 20076 8084 20128 8090
rect 20076 8026 20128 8032
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 20444 7200 20496 7206
rect 20548 7188 20576 9710
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20640 7954 20668 9522
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20640 7410 20668 7890
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20496 7160 20576 7188
rect 20444 7142 20496 7148
rect 19892 6928 19944 6934
rect 19892 6870 19944 6876
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19904 2990 19932 6870
rect 20456 6769 20484 7142
rect 20640 7002 20668 7346
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20442 6760 20498 6769
rect 20442 6695 20498 6704
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20168 6316 20220 6322
rect 20168 6258 20220 6264
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 20180 5574 20208 6258
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 20180 5098 20208 5510
rect 20168 5092 20220 5098
rect 20168 5034 20220 5040
rect 20180 4622 20208 5034
rect 20272 4826 20300 6054
rect 20364 5846 20392 6258
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19996 2990 20024 4490
rect 20088 4282 20116 4558
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 20364 4214 20392 5782
rect 20352 4208 20404 4214
rect 20352 4150 20404 4156
rect 20732 4078 20760 6326
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 20088 3058 20116 3878
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20260 3120 20312 3126
rect 20260 3062 20312 3068
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19524 2508 19576 2514
rect 19524 2450 19576 2456
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 19616 2304 19668 2310
rect 19616 2246 19668 2252
rect 19076 1170 19104 2246
rect 19628 1170 19656 2246
rect 19076 1142 19196 1170
rect 19628 1142 19748 1170
rect 18878 1048 18934 1057
rect 18878 983 18934 992
rect 19168 480 19196 1142
rect 19720 480 19748 1142
rect 20272 480 20300 3062
rect 20364 2514 20392 3470
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20824 480 20852 2246
rect 21376 480 21404 2858
rect 21928 480 21956 3878
rect 22468 2848 22520 2854
rect 22468 2790 22520 2796
rect 22480 480 22508 2790
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3054 0 3110 480
rect 3606 0 3662 480
rect 4158 0 4214 480
rect 4710 0 4766 480
rect 5262 0 5318 480
rect 5814 0 5870 480
rect 6366 0 6422 480
rect 6918 0 6974 480
rect 7470 0 7526 480
rect 8022 0 8078 480
rect 8574 0 8630 480
rect 9126 0 9182 480
rect 9678 0 9734 480
rect 10230 0 10286 480
rect 10782 0 10838 480
rect 11334 0 11390 480
rect 11978 0 12034 480
rect 12530 0 12586 480
rect 13082 0 13138 480
rect 13634 0 13690 480
rect 14186 0 14242 480
rect 14738 0 14794 480
rect 15290 0 15346 480
rect 15842 0 15898 480
rect 16394 0 16450 480
rect 16946 0 17002 480
rect 17498 0 17554 480
rect 18050 0 18106 480
rect 18602 0 18658 480
rect 19154 0 19210 480
rect 19706 0 19762 480
rect 20258 0 20314 480
rect 20810 0 20866 480
rect 21362 0 21418 480
rect 21914 0 21970 480
rect 22466 0 22522 480
<< via2 >>
rect 17958 22480 18014 22536
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 3422 17176 3478 17232
rect 1398 13232 1454 13288
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 8574 15816 8630 15872
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 4066 5788 4068 5808
rect 4068 5788 4120 5808
rect 4120 5788 4122 5808
rect 4066 5752 4122 5788
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 846 2896 902 2952
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 6366 3440 6422 3496
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7562 3576 7618 3632
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 9770 18028 9772 18048
rect 9772 18028 9824 18048
rect 9824 18028 9826 18048
rect 9770 17992 9826 18028
rect 10046 18028 10048 18048
rect 10048 18028 10100 18048
rect 10100 18028 10102 18048
rect 10046 17992 10102 18028
rect 9862 17040 9918 17096
rect 10046 15564 10102 15600
rect 10046 15544 10048 15564
rect 10048 15544 10100 15564
rect 10100 15544 10102 15564
rect 10138 13912 10194 13968
rect 10414 17176 10470 17232
rect 10322 16632 10378 16688
rect 10414 13912 10470 13968
rect 10138 10512 10194 10568
rect 10230 4664 10286 4720
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11518 17740 11574 17776
rect 11518 17720 11520 17740
rect 11520 17720 11572 17740
rect 11572 17720 11574 17740
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11518 16088 11574 16144
rect 12530 18128 12586 18184
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11426 12708 11482 12744
rect 11426 12688 11428 12708
rect 11428 12688 11480 12708
rect 11480 12688 11482 12708
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11150 11056 11206 11112
rect 12070 16088 12126 16144
rect 12162 15952 12218 16008
rect 11978 13232 12034 13288
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11150 9036 11206 9072
rect 11150 9016 11152 9036
rect 11152 9016 11204 9036
rect 11204 9016 11206 9036
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11702 11056 11758 11112
rect 12070 12688 12126 12744
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 10782 2760 10838 2816
rect 10966 3032 11022 3088
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 12346 15952 12402 16008
rect 12346 15852 12348 15872
rect 12348 15852 12400 15872
rect 12400 15852 12402 15872
rect 12346 15816 12402 15852
rect 12806 15952 12862 16008
rect 11794 4020 11796 4040
rect 11796 4020 11848 4040
rect 11848 4020 11850 4040
rect 11794 3984 11850 4020
rect 12806 11192 12862 11248
rect 10966 1536 11022 1592
rect 11978 2760 12034 2816
rect 12162 6296 12218 6352
rect 12162 6196 12164 6216
rect 12164 6196 12216 6216
rect 12216 6196 12218 6216
rect 12162 6160 12218 6196
rect 12346 5888 12402 5944
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 13174 5908 13230 5944
rect 13174 5888 13176 5908
rect 13176 5888 13228 5908
rect 13228 5888 13230 5908
rect 12990 4020 12992 4040
rect 12992 4020 13044 4040
rect 13044 4020 13046 4040
rect 12990 3984 13046 4020
rect 12622 3032 12678 3088
rect 13634 12824 13690 12880
rect 13634 11872 13690 11928
rect 14186 16088 14242 16144
rect 14094 11872 14150 11928
rect 13910 9016 13966 9072
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14738 16668 14740 16688
rect 14740 16668 14792 16688
rect 14792 16668 14794 16688
rect 14738 16632 14794 16668
rect 14738 16224 14794 16280
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 15658 16360 15714 16416
rect 15750 16088 15806 16144
rect 15934 15852 15936 15872
rect 15936 15852 15988 15872
rect 15988 15852 15990 15872
rect 15934 15816 15990 15852
rect 15658 13912 15714 13968
rect 15382 11872 15438 11928
rect 14738 10104 14794 10160
rect 13174 1536 13230 1592
rect 15106 9968 15162 10024
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 15750 11736 15806 11792
rect 15658 10512 15714 10568
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 16118 16668 16120 16688
rect 16120 16668 16172 16688
rect 16172 16668 16174 16688
rect 16118 16632 16174 16668
rect 16486 16768 16542 16824
rect 16486 15952 16542 16008
rect 15658 7384 15714 7440
rect 15290 4800 15346 4856
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 16394 12824 16450 12880
rect 18510 22072 18566 22128
rect 19062 21528 19118 21584
rect 18694 21120 18750 21176
rect 16302 11328 16358 11384
rect 16210 11192 16266 11248
rect 16302 10104 16358 10160
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 16670 10648 16726 10704
rect 16578 10376 16634 10432
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18970 20168 19026 20224
rect 19246 20576 19302 20632
rect 19062 19760 19118 19816
rect 18786 19216 18842 19272
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 17406 17992 17462 18048
rect 17774 17176 17830 17232
rect 17682 17040 17738 17096
rect 17590 15544 17646 15600
rect 17314 12688 17370 12744
rect 16854 9968 16910 10024
rect 16670 7656 16726 7712
rect 16670 6160 16726 6216
rect 16578 3440 16634 3496
rect 17406 11056 17462 11112
rect 17314 10648 17370 10704
rect 18694 18128 18750 18184
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 17958 16940 17960 16960
rect 17960 16940 18012 16960
rect 18012 16940 18014 16960
rect 17958 16904 18014 16940
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18510 12144 18566 12200
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18234 11772 18236 11792
rect 18236 11772 18288 11792
rect 18288 11772 18290 11792
rect 18234 11736 18290 11772
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18510 10376 18566 10432
rect 18418 10004 18420 10024
rect 18420 10004 18472 10024
rect 18472 10004 18474 10024
rect 18418 9968 18474 10004
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 17958 9172 18014 9208
rect 17958 9152 17960 9172
rect 17960 9152 18012 9172
rect 18012 9152 18014 9172
rect 18418 9444 18474 9480
rect 18418 9424 18420 9444
rect 18420 9424 18472 9444
rect 18472 9424 18474 9444
rect 17130 4664 17186 4720
rect 17498 3576 17554 3632
rect 16210 2488 16266 2544
rect 17958 8880 18014 8936
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18142 8472 18198 8528
rect 17866 7792 17922 7848
rect 18050 8084 18106 8120
rect 18050 8064 18052 8084
rect 18052 8064 18104 8084
rect 18104 8064 18106 8084
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 19246 18808 19302 18864
rect 19338 17720 19394 17776
rect 19062 16496 19118 16552
rect 19246 15816 19302 15872
rect 19246 13268 19248 13288
rect 19248 13268 19300 13288
rect 19300 13268 19302 13288
rect 19246 13232 19302 13268
rect 19246 13096 19302 13152
rect 19154 12824 19210 12880
rect 18970 12688 19026 12744
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 17774 6296 17830 6352
rect 18418 6296 18474 6352
rect 18050 5752 18106 5808
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18050 5208 18106 5264
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 17958 4156 17960 4176
rect 17960 4156 18012 4176
rect 18012 4156 18014 4176
rect 17958 4120 18014 4156
rect 17866 1944 17922 2000
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18786 3984 18842 4040
rect 18418 2916 18474 2952
rect 18418 2896 18420 2916
rect 18420 2896 18472 2916
rect 18472 2896 18474 2916
rect 18786 2932 18788 2952
rect 18788 2932 18840 2952
rect 18840 2932 18842 2952
rect 18786 2896 18842 2932
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 17590 584 17646 640
rect 18970 9016 19026 9072
rect 19706 16768 19762 16824
rect 20258 18264 20314 18320
rect 20166 17856 20222 17912
rect 20626 17312 20682 17368
rect 20442 15000 20498 15056
rect 20810 15952 20866 16008
rect 20718 15544 20774 15600
rect 20626 14592 20682 14648
rect 20902 14068 20958 14104
rect 20902 14048 20904 14068
rect 20904 14048 20956 14068
rect 20956 14048 20958 14068
rect 20442 13640 20498 13696
rect 19154 9288 19210 9344
rect 19522 10784 19578 10840
rect 19430 9424 19486 9480
rect 19246 9016 19302 9072
rect 19522 8880 19578 8936
rect 19062 7112 19118 7168
rect 19246 6160 19302 6216
rect 18970 3848 19026 3904
rect 19706 10376 19762 10432
rect 20442 13232 20498 13288
rect 20442 9968 20498 10024
rect 19246 3440 19302 3496
rect 20442 6704 20498 6760
rect 18878 992 18934 1048
<< metal3 >>
rect 17953 22538 18019 22541
rect 22320 22538 22800 22568
rect 17953 22536 22800 22538
rect 17953 22480 17958 22536
rect 18014 22480 22800 22536
rect 17953 22478 22800 22480
rect 17953 22475 18019 22478
rect 22320 22448 22800 22478
rect 18505 22130 18571 22133
rect 22320 22130 22800 22160
rect 18505 22128 22800 22130
rect 18505 22072 18510 22128
rect 18566 22072 22800 22128
rect 18505 22070 22800 22072
rect 18505 22067 18571 22070
rect 22320 22040 22800 22070
rect 19057 21586 19123 21589
rect 22320 21586 22800 21616
rect 19057 21584 22800 21586
rect 19057 21528 19062 21584
rect 19118 21528 22800 21584
rect 19057 21526 22800 21528
rect 19057 21523 19123 21526
rect 22320 21496 22800 21526
rect 18689 21178 18755 21181
rect 22320 21178 22800 21208
rect 18689 21176 22800 21178
rect 18689 21120 18694 21176
rect 18750 21120 22800 21176
rect 18689 21118 22800 21120
rect 18689 21115 18755 21118
rect 22320 21088 22800 21118
rect 19241 20634 19307 20637
rect 22320 20634 22800 20664
rect 19241 20632 22800 20634
rect 19241 20576 19246 20632
rect 19302 20576 22800 20632
rect 19241 20574 22800 20576
rect 19241 20571 19307 20574
rect 22320 20544 22800 20574
rect 18965 20226 19031 20229
rect 22320 20226 22800 20256
rect 18965 20224 22800 20226
rect 18965 20168 18970 20224
rect 19026 20168 22800 20224
rect 18965 20166 22800 20168
rect 18965 20163 19031 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 19057 19818 19123 19821
rect 22320 19818 22800 19848
rect 19057 19816 22800 19818
rect 19057 19760 19062 19816
rect 19118 19760 22800 19816
rect 19057 19758 22800 19760
rect 19057 19755 19123 19758
rect 22320 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 18781 19274 18847 19277
rect 22320 19274 22800 19304
rect 18781 19272 22800 19274
rect 18781 19216 18786 19272
rect 18842 19216 22800 19272
rect 18781 19214 22800 19216
rect 18781 19211 18847 19214
rect 22320 19184 22800 19214
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 19241 18866 19307 18869
rect 22320 18866 22800 18896
rect 19241 18864 22800 18866
rect 19241 18808 19246 18864
rect 19302 18808 22800 18864
rect 19241 18806 22800 18808
rect 19241 18803 19307 18806
rect 22320 18776 22800 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 20253 18322 20319 18325
rect 22320 18322 22800 18352
rect 20253 18320 22800 18322
rect 20253 18264 20258 18320
rect 20314 18264 22800 18320
rect 20253 18262 22800 18264
rect 20253 18259 20319 18262
rect 22320 18232 22800 18262
rect 12525 18186 12591 18189
rect 18689 18186 18755 18189
rect 12525 18184 18755 18186
rect 12525 18128 12530 18184
rect 12586 18128 18694 18184
rect 18750 18128 18755 18184
rect 12525 18126 18755 18128
rect 12525 18123 12591 18126
rect 18689 18123 18755 18126
rect 9765 18050 9831 18053
rect 10041 18050 10107 18053
rect 17401 18052 17467 18053
rect 9765 18048 10107 18050
rect 9765 17992 9770 18048
rect 9826 17992 10046 18048
rect 10102 17992 10107 18048
rect 9765 17990 10107 17992
rect 9765 17987 9831 17990
rect 10041 17987 10107 17990
rect 17350 17988 17356 18052
rect 17420 18050 17467 18052
rect 17420 18048 17512 18050
rect 17462 17992 17512 18048
rect 17420 17990 17512 17992
rect 17420 17988 17467 17990
rect 17401 17987 17467 17988
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 20161 17914 20227 17917
rect 22320 17914 22800 17944
rect 20161 17912 22800 17914
rect 20161 17856 20166 17912
rect 20222 17856 22800 17912
rect 20161 17854 22800 17856
rect 20161 17851 20227 17854
rect 22320 17824 22800 17854
rect 11513 17778 11579 17781
rect 19333 17778 19399 17781
rect 11513 17776 19399 17778
rect 11513 17720 11518 17776
rect 11574 17720 19338 17776
rect 19394 17720 19399 17776
rect 11513 17718 19399 17720
rect 11513 17715 11579 17718
rect 19333 17715 19399 17718
rect 4376 17440 4696 17441
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 20621 17370 20687 17373
rect 22320 17370 22800 17400
rect 20621 17368 22800 17370
rect 20621 17312 20626 17368
rect 20682 17312 22800 17368
rect 20621 17310 22800 17312
rect 20621 17307 20687 17310
rect 22320 17280 22800 17310
rect 0 17234 480 17264
rect 3417 17234 3483 17237
rect 0 17232 3483 17234
rect 0 17176 3422 17232
rect 3478 17176 3483 17232
rect 0 17174 3483 17176
rect 0 17144 480 17174
rect 3417 17171 3483 17174
rect 10409 17234 10475 17237
rect 17769 17234 17835 17237
rect 10409 17232 17835 17234
rect 10409 17176 10414 17232
rect 10470 17176 17774 17232
rect 17830 17176 17835 17232
rect 10409 17174 17835 17176
rect 10409 17171 10475 17174
rect 17769 17171 17835 17174
rect 9857 17098 9923 17101
rect 16798 17098 16804 17100
rect 9857 17096 16804 17098
rect 9857 17040 9862 17096
rect 9918 17040 16804 17096
rect 9857 17038 16804 17040
rect 9857 17035 9923 17038
rect 16798 17036 16804 17038
rect 16868 17098 16874 17100
rect 17677 17098 17743 17101
rect 16868 17096 17743 17098
rect 16868 17040 17682 17096
rect 17738 17040 17743 17096
rect 16868 17038 17743 17040
rect 16868 17036 16874 17038
rect 17677 17035 17743 17038
rect 17953 16962 18019 16965
rect 22320 16962 22800 16992
rect 17953 16960 22800 16962
rect 17953 16904 17958 16960
rect 18014 16904 22800 16960
rect 17953 16902 22800 16904
rect 17953 16899 18019 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 22320 16872 22800 16902
rect 14672 16831 14992 16832
rect 16481 16826 16547 16829
rect 19701 16826 19767 16829
rect 15702 16824 19767 16826
rect 15702 16768 16486 16824
rect 16542 16768 19706 16824
rect 19762 16768 19767 16824
rect 15702 16766 19767 16768
rect 10317 16690 10383 16693
rect 14733 16690 14799 16693
rect 10317 16688 14799 16690
rect 10317 16632 10322 16688
rect 10378 16632 14738 16688
rect 14794 16632 14799 16688
rect 10317 16630 14799 16632
rect 10317 16627 10383 16630
rect 14733 16627 14799 16630
rect 15702 16421 15762 16766
rect 16481 16763 16547 16766
rect 19701 16763 19767 16766
rect 16113 16690 16179 16693
rect 16246 16690 16252 16692
rect 16113 16688 16252 16690
rect 16113 16632 16118 16688
rect 16174 16632 16252 16688
rect 16113 16630 16252 16632
rect 16113 16627 16179 16630
rect 16246 16628 16252 16630
rect 16316 16628 16322 16692
rect 19057 16554 19123 16557
rect 22320 16554 22800 16584
rect 19057 16552 22800 16554
rect 19057 16496 19062 16552
rect 19118 16496 22800 16552
rect 19057 16494 22800 16496
rect 19057 16491 19123 16494
rect 22320 16464 22800 16494
rect 15653 16416 15762 16421
rect 15653 16360 15658 16416
rect 15714 16360 15762 16416
rect 15653 16358 15762 16360
rect 15653 16355 15719 16358
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 14733 16282 14799 16285
rect 15142 16282 15148 16284
rect 14733 16280 15148 16282
rect 14733 16224 14738 16280
rect 14794 16224 15148 16280
rect 14733 16222 15148 16224
rect 14733 16219 14799 16222
rect 15142 16220 15148 16222
rect 15212 16220 15218 16284
rect 11513 16146 11579 16149
rect 12065 16146 12131 16149
rect 11513 16144 12131 16146
rect 11513 16088 11518 16144
rect 11574 16088 12070 16144
rect 12126 16088 12131 16144
rect 11513 16086 12131 16088
rect 11513 16083 11579 16086
rect 12065 16083 12131 16086
rect 14181 16146 14247 16149
rect 15745 16146 15811 16149
rect 14181 16144 15811 16146
rect 14181 16088 14186 16144
rect 14242 16088 15750 16144
rect 15806 16088 15811 16144
rect 14181 16086 15811 16088
rect 14181 16083 14247 16086
rect 15745 16083 15811 16086
rect 12157 16010 12223 16013
rect 12341 16010 12407 16013
rect 12157 16008 12407 16010
rect 12157 15952 12162 16008
rect 12218 15952 12346 16008
rect 12402 15952 12407 16008
rect 12157 15950 12407 15952
rect 12157 15947 12223 15950
rect 12341 15947 12407 15950
rect 12801 16010 12867 16013
rect 16481 16010 16547 16013
rect 12801 16008 16547 16010
rect 12801 15952 12806 16008
rect 12862 15952 16486 16008
rect 16542 15952 16547 16008
rect 12801 15950 16547 15952
rect 12801 15947 12867 15950
rect 16481 15947 16547 15950
rect 20805 16010 20871 16013
rect 22320 16010 22800 16040
rect 20805 16008 22800 16010
rect 20805 15952 20810 16008
rect 20866 15952 22800 16008
rect 20805 15950 22800 15952
rect 20805 15947 20871 15950
rect 22320 15920 22800 15950
rect 8569 15874 8635 15877
rect 12341 15874 12407 15877
rect 8569 15872 12407 15874
rect 8569 15816 8574 15872
rect 8630 15816 12346 15872
rect 12402 15816 12407 15872
rect 8569 15814 12407 15816
rect 8569 15811 8635 15814
rect 12341 15811 12407 15814
rect 15929 15874 15995 15877
rect 19241 15874 19307 15877
rect 15929 15872 19307 15874
rect 15929 15816 15934 15872
rect 15990 15816 19246 15872
rect 19302 15816 19307 15872
rect 15929 15814 19307 15816
rect 15929 15811 15995 15814
rect 19241 15811 19307 15814
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 10041 15602 10107 15605
rect 17585 15602 17651 15605
rect 10041 15600 17651 15602
rect 10041 15544 10046 15600
rect 10102 15544 17590 15600
rect 17646 15544 17651 15600
rect 10041 15542 17651 15544
rect 10041 15539 10107 15542
rect 17585 15539 17651 15542
rect 20713 15602 20779 15605
rect 22320 15602 22800 15632
rect 20713 15600 22800 15602
rect 20713 15544 20718 15600
rect 20774 15544 22800 15600
rect 20713 15542 22800 15544
rect 20713 15539 20779 15542
rect 22320 15512 22800 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 20437 15058 20503 15061
rect 22320 15058 22800 15088
rect 20437 15056 22800 15058
rect 20437 15000 20442 15056
rect 20498 15000 22800 15056
rect 20437 14998 22800 15000
rect 20437 14995 20503 14998
rect 22320 14968 22800 14998
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 20621 14650 20687 14653
rect 22320 14650 22800 14680
rect 20621 14648 22800 14650
rect 20621 14592 20626 14648
rect 20682 14592 22800 14648
rect 20621 14590 22800 14592
rect 20621 14587 20687 14590
rect 22320 14560 22800 14590
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 20897 14106 20963 14109
rect 22320 14106 22800 14136
rect 20897 14104 22800 14106
rect 20897 14048 20902 14104
rect 20958 14048 22800 14104
rect 20897 14046 22800 14048
rect 20897 14043 20963 14046
rect 22320 14016 22800 14046
rect 10133 13970 10199 13973
rect 10409 13970 10475 13973
rect 15653 13970 15719 13973
rect 10133 13968 15719 13970
rect 10133 13912 10138 13968
rect 10194 13912 10414 13968
rect 10470 13912 15658 13968
rect 15714 13912 15719 13968
rect 10133 13910 15719 13912
rect 10133 13907 10199 13910
rect 10409 13907 10475 13910
rect 15653 13907 15719 13910
rect 20437 13698 20503 13701
rect 22320 13698 22800 13728
rect 20437 13696 22800 13698
rect 20437 13640 20442 13696
rect 20498 13640 22800 13696
rect 20437 13638 22800 13640
rect 20437 13635 20503 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22320 13608 22800 13638
rect 14672 13567 14992 13568
rect 1393 13290 1459 13293
rect 11973 13290 12039 13293
rect 19241 13290 19307 13293
rect 1393 13288 19307 13290
rect 1393 13232 1398 13288
rect 1454 13232 11978 13288
rect 12034 13232 19246 13288
rect 19302 13232 19307 13288
rect 1393 13230 19307 13232
rect 1393 13227 1459 13230
rect 11973 13227 12039 13230
rect 19241 13227 19307 13230
rect 20437 13290 20503 13293
rect 22320 13290 22800 13320
rect 20437 13288 22800 13290
rect 20437 13232 20442 13288
rect 20498 13232 22800 13288
rect 20437 13230 22800 13232
rect 20437 13227 20503 13230
rect 22320 13200 22800 13230
rect 19241 13156 19307 13157
rect 19190 13154 19196 13156
rect 19150 13094 19196 13154
rect 19260 13152 19307 13156
rect 19302 13096 19307 13152
rect 19190 13092 19196 13094
rect 19260 13092 19307 13096
rect 19241 13091 19307 13092
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 13629 12882 13695 12885
rect 16389 12882 16455 12885
rect 18638 12882 18644 12884
rect 13629 12880 18644 12882
rect 13629 12824 13634 12880
rect 13690 12824 16394 12880
rect 16450 12824 18644 12880
rect 13629 12822 18644 12824
rect 13629 12819 13695 12822
rect 16389 12819 16455 12822
rect 18638 12820 18644 12822
rect 18708 12882 18714 12884
rect 19149 12882 19215 12885
rect 18708 12880 19215 12882
rect 18708 12824 19154 12880
rect 19210 12824 19215 12880
rect 18708 12822 19215 12824
rect 18708 12820 18714 12822
rect 19149 12819 19215 12822
rect 11421 12746 11487 12749
rect 12065 12746 12131 12749
rect 17309 12746 17375 12749
rect 11421 12744 17375 12746
rect 11421 12688 11426 12744
rect 11482 12688 12070 12744
rect 12126 12688 17314 12744
rect 17370 12688 17375 12744
rect 11421 12686 17375 12688
rect 11421 12683 11487 12686
rect 12065 12683 12131 12686
rect 17309 12683 17375 12686
rect 18965 12746 19031 12749
rect 22320 12746 22800 12776
rect 18965 12744 22800 12746
rect 18965 12688 18970 12744
rect 19026 12688 22800 12744
rect 18965 12686 22800 12688
rect 18965 12683 19031 12686
rect 22320 12656 22800 12686
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 22320 12338 22800 12368
rect 18646 12278 22800 12338
rect 18505 12202 18571 12205
rect 18646 12202 18706 12278
rect 22320 12248 22800 12278
rect 18505 12200 18706 12202
rect 18505 12144 18510 12200
rect 18566 12144 18706 12200
rect 18505 12142 18706 12144
rect 18505 12139 18571 12142
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 13629 11930 13695 11933
rect 14089 11930 14155 11933
rect 13629 11928 14155 11930
rect 13629 11872 13634 11928
rect 13690 11872 14094 11928
rect 14150 11872 14155 11928
rect 13629 11870 14155 11872
rect 13629 11867 13695 11870
rect 14089 11867 14155 11870
rect 15377 11930 15443 11933
rect 15377 11928 15762 11930
rect 15377 11872 15382 11928
rect 15438 11872 15762 11928
rect 15377 11870 15762 11872
rect 15377 11867 15443 11870
rect 15702 11797 15762 11870
rect 15702 11792 15811 11797
rect 15702 11736 15750 11792
rect 15806 11736 15811 11792
rect 15702 11734 15811 11736
rect 15745 11731 15811 11734
rect 18229 11794 18295 11797
rect 22320 11794 22800 11824
rect 18229 11792 22800 11794
rect 18229 11736 18234 11792
rect 18290 11736 22800 11792
rect 18229 11734 22800 11736
rect 18229 11731 18295 11734
rect 22320 11704 22800 11734
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 16297 11386 16363 11389
rect 22320 11386 22800 11416
rect 16297 11384 22800 11386
rect 16297 11328 16302 11384
rect 16358 11328 22800 11384
rect 16297 11326 22800 11328
rect 16297 11323 16363 11326
rect 22320 11296 22800 11326
rect 12801 11250 12867 11253
rect 16205 11250 16271 11253
rect 12801 11248 16271 11250
rect 12801 11192 12806 11248
rect 12862 11192 16210 11248
rect 16266 11192 16271 11248
rect 12801 11190 16271 11192
rect 12801 11187 12867 11190
rect 16205 11187 16271 11190
rect 11145 11114 11211 11117
rect 11697 11114 11763 11117
rect 11145 11112 11763 11114
rect 11145 11056 11150 11112
rect 11206 11056 11702 11112
rect 11758 11056 11763 11112
rect 11145 11054 11763 11056
rect 11145 11051 11211 11054
rect 11697 11051 11763 11054
rect 16246 11052 16252 11116
rect 16316 11114 16322 11116
rect 17401 11114 17467 11117
rect 16316 11112 17467 11114
rect 16316 11056 17406 11112
rect 17462 11056 17467 11112
rect 16316 11054 17467 11056
rect 16316 11052 16322 11054
rect 17401 11051 17467 11054
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 19517 10842 19583 10845
rect 22320 10842 22800 10872
rect 19517 10840 22800 10842
rect 19517 10784 19522 10840
rect 19578 10784 22800 10840
rect 19517 10782 22800 10784
rect 19517 10779 19583 10782
rect 22320 10752 22800 10782
rect 16665 10706 16731 10709
rect 17309 10706 17375 10709
rect 16665 10704 17375 10706
rect 16665 10648 16670 10704
rect 16726 10648 17314 10704
rect 17370 10648 17375 10704
rect 16665 10646 17375 10648
rect 16665 10643 16731 10646
rect 17309 10643 17375 10646
rect 10133 10570 10199 10573
rect 15653 10570 15719 10573
rect 10133 10568 15719 10570
rect 10133 10512 10138 10568
rect 10194 10512 15658 10568
rect 15714 10512 15719 10568
rect 10133 10510 15719 10512
rect 10133 10507 10199 10510
rect 15653 10507 15719 10510
rect 16573 10434 16639 10437
rect 17350 10434 17356 10436
rect 16573 10432 17356 10434
rect 16573 10376 16578 10432
rect 16634 10376 17356 10432
rect 16573 10374 17356 10376
rect 16573 10371 16639 10374
rect 17350 10372 17356 10374
rect 17420 10434 17426 10436
rect 18505 10434 18571 10437
rect 17420 10432 18571 10434
rect 17420 10376 18510 10432
rect 18566 10376 18571 10432
rect 17420 10374 18571 10376
rect 17420 10372 17426 10374
rect 18505 10371 18571 10374
rect 19701 10434 19767 10437
rect 22320 10434 22800 10464
rect 19701 10432 22800 10434
rect 19701 10376 19706 10432
rect 19762 10376 22800 10432
rect 19701 10374 22800 10376
rect 19701 10371 19767 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22320 10344 22800 10374
rect 14672 10303 14992 10304
rect 14733 10162 14799 10165
rect 16297 10162 16363 10165
rect 14733 10160 16363 10162
rect 14733 10104 14738 10160
rect 14794 10104 16302 10160
rect 16358 10104 16363 10160
rect 14733 10102 16363 10104
rect 14733 10099 14799 10102
rect 16297 10099 16363 10102
rect 15101 10028 15167 10029
rect 16849 10028 16915 10029
rect 15101 10024 15148 10028
rect 15212 10026 15218 10028
rect 15101 9968 15106 10024
rect 15101 9964 15148 9968
rect 15212 9966 15258 10026
rect 15212 9964 15218 9966
rect 16798 9964 16804 10028
rect 16868 10026 16915 10028
rect 18413 10026 18479 10029
rect 18822 10026 18828 10028
rect 16868 10024 16960 10026
rect 16910 9968 16960 10024
rect 16868 9966 16960 9968
rect 18413 10024 18828 10026
rect 18413 9968 18418 10024
rect 18474 9968 18828 10024
rect 18413 9966 18828 9968
rect 16868 9964 16915 9966
rect 15101 9963 15167 9964
rect 16849 9963 16915 9964
rect 18413 9963 18479 9966
rect 18822 9964 18828 9966
rect 18892 9964 18898 10028
rect 20437 10026 20503 10029
rect 22320 10026 22800 10056
rect 20437 10024 22800 10026
rect 20437 9968 20442 10024
rect 20498 9968 22800 10024
rect 20437 9966 22800 9968
rect 20437 9963 20503 9966
rect 22320 9936 22800 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 18413 9482 18479 9485
rect 19425 9482 19491 9485
rect 22320 9482 22800 9512
rect 18413 9480 22800 9482
rect 18413 9424 18418 9480
rect 18474 9424 19430 9480
rect 19486 9424 22800 9480
rect 18413 9422 22800 9424
rect 18413 9419 18479 9422
rect 19425 9419 19491 9422
rect 22320 9392 22800 9422
rect 19006 9284 19012 9348
rect 19076 9346 19082 9348
rect 19149 9346 19215 9349
rect 19076 9344 19215 9346
rect 19076 9288 19154 9344
rect 19210 9288 19215 9344
rect 19076 9286 19215 9288
rect 19076 9284 19082 9286
rect 19149 9283 19215 9286
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 17953 9210 18019 9213
rect 17953 9208 19442 9210
rect 17953 9152 17958 9208
rect 18014 9152 19442 9208
rect 17953 9150 19442 9152
rect 17953 9147 18019 9150
rect 11145 9074 11211 9077
rect 13905 9074 13971 9077
rect 11145 9072 13971 9074
rect 11145 9016 11150 9072
rect 11206 9016 13910 9072
rect 13966 9016 13971 9072
rect 11145 9014 13971 9016
rect 11145 9011 11211 9014
rect 13905 9011 13971 9014
rect 18822 9012 18828 9076
rect 18892 9074 18898 9076
rect 18965 9074 19031 9077
rect 19241 9076 19307 9077
rect 19190 9074 19196 9076
rect 18892 9072 19031 9074
rect 18892 9016 18970 9072
rect 19026 9016 19031 9072
rect 18892 9014 19031 9016
rect 19150 9014 19196 9074
rect 19260 9072 19307 9076
rect 19302 9016 19307 9072
rect 18892 9012 18898 9014
rect 18965 9011 19031 9014
rect 19190 9012 19196 9014
rect 19260 9012 19307 9016
rect 19382 9074 19442 9150
rect 22320 9074 22800 9104
rect 19382 9014 22800 9074
rect 19241 9011 19307 9012
rect 22320 8984 22800 9014
rect 17953 8938 18019 8941
rect 19517 8938 19583 8941
rect 17953 8936 19583 8938
rect 17953 8880 17958 8936
rect 18014 8880 19522 8936
rect 19578 8880 19583 8936
rect 17953 8878 19583 8880
rect 17953 8875 18019 8878
rect 19517 8875 19583 8878
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 18137 8530 18203 8533
rect 22320 8530 22800 8560
rect 18137 8528 22800 8530
rect 18137 8472 18142 8528
rect 18198 8472 22800 8528
rect 18137 8470 22800 8472
rect 18137 8467 18203 8470
rect 22320 8440 22800 8470
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 18045 8122 18111 8125
rect 22320 8122 22800 8152
rect 18045 8120 22800 8122
rect 18045 8064 18050 8120
rect 18106 8064 22800 8120
rect 18045 8062 22800 8064
rect 18045 8059 18111 8062
rect 22320 8032 22800 8062
rect 17861 7848 17927 7853
rect 17861 7792 17866 7848
rect 17922 7792 17927 7848
rect 17861 7787 17927 7792
rect 16665 7714 16731 7717
rect 17864 7714 17924 7787
rect 16665 7712 17924 7714
rect 16665 7656 16670 7712
rect 16726 7656 17924 7712
rect 16665 7654 17924 7656
rect 16665 7651 16731 7654
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 22320 7578 22800 7608
rect 18508 7518 22800 7578
rect 15653 7442 15719 7445
rect 18508 7442 18568 7518
rect 22320 7488 22800 7518
rect 15653 7440 18568 7442
rect 15653 7384 15658 7440
rect 15714 7384 18568 7440
rect 15653 7382 18568 7384
rect 15653 7379 15719 7382
rect 19057 7170 19123 7173
rect 22320 7170 22800 7200
rect 19057 7168 22800 7170
rect 19057 7112 19062 7168
rect 19118 7112 22800 7168
rect 19057 7110 22800 7112
rect 19057 7107 19123 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 22320 7080 22800 7110
rect 14672 7039 14992 7040
rect 20437 6762 20503 6765
rect 22320 6762 22800 6792
rect 20437 6760 22800 6762
rect 20437 6704 20442 6760
rect 20498 6704 22800 6760
rect 20437 6702 22800 6704
rect 20437 6699 20503 6702
rect 22320 6672 22800 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 12157 6354 12223 6357
rect 17769 6354 17835 6357
rect 18413 6354 18479 6357
rect 12157 6352 18479 6354
rect 12157 6296 12162 6352
rect 12218 6296 17774 6352
rect 17830 6296 18418 6352
rect 18474 6296 18479 6352
rect 12157 6294 18479 6296
rect 12157 6291 12223 6294
rect 17769 6291 17835 6294
rect 18413 6291 18479 6294
rect 12157 6218 12223 6221
rect 16665 6218 16731 6221
rect 12157 6216 16731 6218
rect 12157 6160 12162 6216
rect 12218 6160 16670 6216
rect 16726 6160 16731 6216
rect 12157 6158 16731 6160
rect 12157 6155 12223 6158
rect 16665 6155 16731 6158
rect 19241 6218 19307 6221
rect 22320 6218 22800 6248
rect 19241 6216 22800 6218
rect 19241 6160 19246 6216
rect 19302 6160 22800 6216
rect 19241 6158 22800 6160
rect 19241 6155 19307 6158
rect 22320 6128 22800 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 12341 5946 12407 5949
rect 13169 5946 13235 5949
rect 12341 5944 13235 5946
rect 12341 5888 12346 5944
rect 12402 5888 13174 5944
rect 13230 5888 13235 5944
rect 12341 5886 13235 5888
rect 12341 5883 12407 5886
rect 13169 5883 13235 5886
rect 0 5810 480 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 480 5750
rect 4061 5747 4127 5750
rect 18045 5810 18111 5813
rect 22320 5810 22800 5840
rect 18045 5808 22800 5810
rect 18045 5752 18050 5808
rect 18106 5752 22800 5808
rect 18045 5750 22800 5752
rect 18045 5747 18111 5750
rect 22320 5720 22800 5750
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 18045 5266 18111 5269
rect 22320 5266 22800 5296
rect 18045 5264 22800 5266
rect 18045 5208 18050 5264
rect 18106 5208 22800 5264
rect 18045 5206 22800 5208
rect 18045 5203 18111 5206
rect 22320 5176 22800 5206
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 15285 4858 15351 4861
rect 22320 4858 22800 4888
rect 15285 4856 22800 4858
rect 15285 4800 15290 4856
rect 15346 4800 22800 4856
rect 15285 4798 22800 4800
rect 15285 4795 15351 4798
rect 22320 4768 22800 4798
rect 10225 4722 10291 4725
rect 17125 4722 17191 4725
rect 10225 4720 17191 4722
rect 10225 4664 10230 4720
rect 10286 4664 17130 4720
rect 17186 4664 17191 4720
rect 10225 4662 17191 4664
rect 10225 4659 10291 4662
rect 17125 4659 17191 4662
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 22320 4314 22800 4344
rect 18646 4254 22800 4314
rect 17953 4178 18019 4181
rect 18646 4178 18706 4254
rect 22320 4224 22800 4254
rect 17953 4176 18706 4178
rect 17953 4120 17958 4176
rect 18014 4120 18706 4176
rect 17953 4118 18706 4120
rect 17953 4115 18019 4118
rect 11789 4042 11855 4045
rect 12985 4042 13051 4045
rect 11789 4040 13051 4042
rect 11789 3984 11794 4040
rect 11850 3984 12990 4040
rect 13046 3984 13051 4040
rect 11789 3982 13051 3984
rect 11789 3979 11855 3982
rect 12985 3979 13051 3982
rect 18638 3980 18644 4044
rect 18708 4042 18714 4044
rect 18781 4042 18847 4045
rect 18708 4040 18847 4042
rect 18708 3984 18786 4040
rect 18842 3984 18847 4040
rect 18708 3982 18847 3984
rect 18708 3980 18714 3982
rect 18781 3979 18847 3982
rect 18965 3906 19031 3909
rect 22320 3906 22800 3936
rect 18965 3904 22800 3906
rect 18965 3848 18970 3904
rect 19026 3848 22800 3904
rect 18965 3846 22800 3848
rect 18965 3843 19031 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22320 3816 22800 3846
rect 14672 3775 14992 3776
rect 7557 3634 7623 3637
rect 17493 3634 17559 3637
rect 7557 3632 17559 3634
rect 7557 3576 7562 3632
rect 7618 3576 17498 3632
rect 17554 3576 17559 3632
rect 7557 3574 17559 3576
rect 7557 3571 7623 3574
rect 17493 3571 17559 3574
rect 6361 3498 6427 3501
rect 16573 3498 16639 3501
rect 6361 3496 16639 3498
rect 6361 3440 6366 3496
rect 6422 3440 16578 3496
rect 16634 3440 16639 3496
rect 6361 3438 16639 3440
rect 6361 3435 6427 3438
rect 16573 3435 16639 3438
rect 19241 3498 19307 3501
rect 22320 3498 22800 3528
rect 19241 3496 22800 3498
rect 19241 3440 19246 3496
rect 19302 3440 22800 3496
rect 19241 3438 22800 3440
rect 19241 3435 19307 3438
rect 22320 3408 22800 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 10961 3090 11027 3093
rect 12617 3090 12683 3093
rect 10961 3088 12683 3090
rect 10961 3032 10966 3088
rect 11022 3032 12622 3088
rect 12678 3032 12683 3088
rect 10961 3030 12683 3032
rect 10961 3027 11027 3030
rect 12617 3027 12683 3030
rect 841 2954 907 2957
rect 18413 2954 18479 2957
rect 841 2952 18479 2954
rect 841 2896 846 2952
rect 902 2896 18418 2952
rect 18474 2896 18479 2952
rect 841 2894 18479 2896
rect 841 2891 907 2894
rect 18413 2891 18479 2894
rect 18781 2954 18847 2957
rect 22320 2954 22800 2984
rect 18781 2952 22800 2954
rect 18781 2896 18786 2952
rect 18842 2896 22800 2952
rect 18781 2894 22800 2896
rect 18781 2891 18847 2894
rect 22320 2864 22800 2894
rect 10777 2818 10843 2821
rect 11973 2818 12039 2821
rect 10777 2816 12039 2818
rect 10777 2760 10782 2816
rect 10838 2760 11978 2816
rect 12034 2760 12039 2816
rect 10777 2758 12039 2760
rect 10777 2755 10843 2758
rect 11973 2755 12039 2758
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 16205 2546 16271 2549
rect 22320 2546 22800 2576
rect 16205 2544 22800 2546
rect 16205 2488 16210 2544
rect 16266 2488 22800 2544
rect 16205 2486 22800 2488
rect 16205 2483 16271 2486
rect 22320 2456 22800 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 17861 2002 17927 2005
rect 22320 2002 22800 2032
rect 17861 2000 22800 2002
rect 17861 1944 17866 2000
rect 17922 1944 22800 2000
rect 17861 1942 22800 1944
rect 17861 1939 17927 1942
rect 22320 1912 22800 1942
rect 10961 1594 11027 1597
rect 13169 1594 13235 1597
rect 22320 1594 22800 1624
rect 10961 1592 22800 1594
rect 10961 1536 10966 1592
rect 11022 1536 13174 1592
rect 13230 1536 22800 1592
rect 10961 1534 22800 1536
rect 10961 1531 11027 1534
rect 13169 1531 13235 1534
rect 22320 1504 22800 1534
rect 18873 1050 18939 1053
rect 22320 1050 22800 1080
rect 18873 1048 22800 1050
rect 18873 992 18878 1048
rect 18934 992 22800 1048
rect 18873 990 22800 992
rect 18873 987 18939 990
rect 22320 960 22800 990
rect 17585 642 17651 645
rect 22320 642 22800 672
rect 17585 640 22800 642
rect 17585 584 17590 640
rect 17646 584 22800 640
rect 17585 582 22800 584
rect 17585 579 17651 582
rect 22320 552 22800 582
rect 19006 172 19012 236
rect 19076 234 19082 236
rect 22320 234 22800 264
rect 19076 174 22800 234
rect 19076 172 19082 174
rect 22320 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 17356 18048 17420 18052
rect 17356 17992 17406 18048
rect 17406 17992 17420 18048
rect 17356 17988 17420 17992
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 16804 17036 16868 17100
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 16252 16628 16316 16692
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 15148 16220 15212 16284
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 19196 13152 19260 13156
rect 19196 13096 19246 13152
rect 19246 13096 19260 13152
rect 19196 13092 19260 13096
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 18644 12820 18708 12884
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 16252 11052 16316 11116
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 17356 10372 17420 10436
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 15148 10024 15212 10028
rect 15148 9968 15162 10024
rect 15162 9968 15212 10024
rect 15148 9964 15212 9968
rect 16804 10024 16868 10028
rect 16804 9968 16854 10024
rect 16854 9968 16868 10024
rect 16804 9964 16868 9968
rect 18828 9964 18892 10028
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 19012 9284 19076 9348
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 18828 9012 18892 9076
rect 19196 9072 19260 9076
rect 19196 9016 19246 9072
rect 19246 9016 19260 9072
rect 19196 9012 19260 9016
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 18644 3980 18708 4044
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
rect 19012 172 19076 236
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 17355 18052 17421 18053
rect 17355 17988 17356 18052
rect 17420 17988 17421 18052
rect 17355 17987 17421 17988
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 16803 17100 16869 17101
rect 16803 17036 16804 17100
rect 16868 17036 16869 17100
rect 16803 17035 16869 17036
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 16251 16692 16317 16693
rect 16251 16628 16252 16692
rect 16316 16628 16317 16692
rect 16251 16627 16317 16628
rect 15147 16284 15213 16285
rect 15147 16220 15148 16284
rect 15212 16220 15213 16284
rect 15147 16219 15213 16220
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 15150 10029 15210 16219
rect 16254 11117 16314 16627
rect 16251 11116 16317 11117
rect 16251 11052 16252 11116
rect 16316 11052 16317 11116
rect 16251 11051 16317 11052
rect 16806 10029 16866 17035
rect 17358 10437 17418 17987
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 19195 13156 19261 13157
rect 19195 13092 19196 13156
rect 19260 13092 19261 13156
rect 19195 13091 19261 13092
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18643 12884 18709 12885
rect 18643 12820 18644 12884
rect 18708 12820 18709 12884
rect 18643 12819 18709 12820
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 17355 10436 17421 10437
rect 17355 10372 17356 10436
rect 17420 10372 17421 10436
rect 17355 10371 17421 10372
rect 15147 10028 15213 10029
rect 15147 9964 15148 10028
rect 15212 9964 15213 10028
rect 15147 9963 15213 9964
rect 16803 10028 16869 10029
rect 16803 9964 16804 10028
rect 16868 9964 16869 10028
rect 16803 9963 16869 9964
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18646 4045 18706 12819
rect 18827 10028 18893 10029
rect 18827 9964 18828 10028
rect 18892 9964 18893 10028
rect 18827 9963 18893 9964
rect 18830 9077 18890 9963
rect 19011 9348 19077 9349
rect 19011 9284 19012 9348
rect 19076 9284 19077 9348
rect 19011 9283 19077 9284
rect 18827 9076 18893 9077
rect 18827 9012 18828 9076
rect 18892 9012 18893 9076
rect 18827 9011 18893 9012
rect 18643 4044 18709 4045
rect 18643 3980 18644 4044
rect 18708 3980 18709 4044
rect 18643 3979 18709 3980
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
rect 19014 237 19074 9283
rect 19198 9077 19258 13091
rect 19195 9076 19261 9077
rect 19195 9012 19196 9076
rect 19260 9012 19261 9076
rect 19195 9011 19261 9012
rect 19011 236 19077 237
rect 19011 172 19012 236
rect 19076 172 19077 236
rect 19011 171 19077 172
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1605641404
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1605641404
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1605641404
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1605641404
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1605641404
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1605641404
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1605641404
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _105_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10304 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10672 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1605641404
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1605641404
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1605641404
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1605641404
transform 1 0 11132 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1605641404
transform 1 0 11500 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1605641404
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1605641404
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1605641404
transform 1 0 11776 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1605641404
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1605641404
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1605641404
transform 1 0 11960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1605641404
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 14260 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13340 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13248 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1605641404
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_139
timestamp 1605641404
transform 1 0 13892 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_129
timestamp 1605641404
transform 1 0 12972 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_141
timestamp 1605641404
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1605641404
transform 1 0 15916 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1605641404
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1605641404
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1605641404
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1605641404
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_159
timestamp 1605641404
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_165
timestamp 1605641404
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_176
timestamp 1605641404
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_175 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 17204 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_171
timestamp 1605641404
transform 1 0 16836 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16468 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1605641404
transform 1 0 16468 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1605641404
transform 1 0 17296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1605641404
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1605641404
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _041_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 17480 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1605641404
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_191
timestamp 1605641404
transform 1 0 18676 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_195
timestamp 1605641404
transform 1 0 19044 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1605641404
transform 1 0 18952 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_202
timestamp 1605641404
transform 1 0 19688 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_198
timestamp 1605641404
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1605641404
transform 1 0 19504 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1605641404
transform 1 0 19320 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1605641404
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1605641404
transform 1 0 19964 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_208
timestamp 1605641404
transform 1 0 20240 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1605641404
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1605641404
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1605641404
transform 1 0 20332 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1605641404
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1605641404
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1605641404
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1605641404
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1605641404
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1605641404
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1605641404
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1605641404
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1605641404
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1605641404
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9936 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11592 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_112
timestamp 1605641404
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13248 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_130
timestamp 1605641404
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15548 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1605641404
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1605641404
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 17204 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 1605641404
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19044 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19780 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1605641404
transform 1 0 18676 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_201
timestamp 1605641404
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1605641404
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1605641404
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1605641404
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1605641404
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1605641404
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1605641404
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1605641404
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1605641404
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1605641404
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_74
timestamp 1605641404
transform 1 0 7912 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_82
timestamp 1605641404
transform 1 0 8648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8924 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_3_101
timestamp 1605641404
transform 1 0 10396 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1605641404
transform 1 0 10948 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1605641404
transform 1 0 11776 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_110
timestamp 1605641404
transform 1 0 11224 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1605641404
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_123
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1605641404
transform 1 0 13432 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12696 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13892 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1605641404
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_137
timestamp 1605641404
transform 1 0 13708 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15272 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16284 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_148
timestamp 1605641404
transform 1 0 14720 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_163
timestamp 1605641404
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1605641404
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18032 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_171
timestamp 1605641404
transform 1 0 16836 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1605641404
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19688 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1605641404
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1605641404
transform 1 0 20700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1605641404
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 1605641404
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1605641404
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1605641404
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1605641404
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1605641404
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1605641404
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1605641404
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1605641404
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_117
timestamp 1605641404
transform 1 0 11868 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1605641404
transform 1 0 14444 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13432 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_132
timestamp 1605641404
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_143
timestamp 1605641404
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1605641404
transform 1 0 15640 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1605641404
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18032 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_167
timestamp 1605641404
transform 1 0 16468 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_179
timestamp 1605641404
transform 1 0 17572 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_183
timestamp 1605641404
transform 1 0 17940 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1605641404
transform 1 0 19044 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19596 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_193
timestamp 1605641404
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_198
timestamp 1605641404
transform 1 0 19320 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1605641404
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1605641404
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1605641404
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1605641404
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1605641404
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1605641404
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1605641404
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1605641404
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10304 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1605641404
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_98
timestamp 1605641404
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1605641404
transform 1 0 11868 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_109
timestamp 1605641404
transform 1 0 11132 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1605641404
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14076 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_139
timestamp 1605641404
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 15916 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_157
timestamp 1605641404
transform 1 0 15548 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1605641404
transform 1 0 18216 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_177
timestamp 1605641404
transform 1 0 17388 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1605641404
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 19228 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_195
timestamp 1605641404
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_213
timestamp 1605641404
transform 1 0 20700 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1605641404
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1605641404
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1605641404
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1605641404
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1605641404
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1605641404
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6440 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1605641404
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_56
timestamp 1605641404
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1605641404
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1605641404
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7636 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1605641404
transform 1 0 7912 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1605641404
transform 1 0 7544 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1605641404
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1605641404
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_86
timestamp 1605641404
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9292 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1605641404
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_98
timestamp 1605641404
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_102
timestamp 1605641404
transform 1 0 10488 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10304 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10856 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12512 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 11316 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_122
timestamp 1605641404
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_109
timestamp 1605641404
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1605641404
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13432 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1605641404
transform 1 0 13524 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_133
timestamp 1605641404
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_144
timestamp 1605641404
transform 1 0 14352 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1605641404
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_143
timestamp 1605641404
transform 1 0 14260 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15272 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1605641404
transform 1 0 16284 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1605641404
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_151
timestamp 1605641404
transform 1 0 14996 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_163
timestamp 1605641404
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 17112 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_170
timestamp 1605641404
transform 1 0 16744 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_174
timestamp 1605641404
transform 1 0 17112 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1605641404
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18768 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1605641404
transform 1 0 20240 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1605641404
transform 1 0 19228 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_190
timestamp 1605641404
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_208
timestamp 1605641404
transform 1 0 20240 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1605641404
transform 1 0 18860 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_206
timestamp 1605641404
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1605641404
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_218
timestamp 1605641404
transform 1 0 21160 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_217
timestamp 1605641404
transform 1 0 21068 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1605641404
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1605641404
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1605641404
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1605641404
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7912 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_8_68
timestamp 1605641404
transform 1 0 7360 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1605641404
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_102
timestamp 1605641404
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11500 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10764 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_108
timestamp 1605641404
transform 1 0 11040 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_112
timestamp 1605641404
transform 1 0 11408 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13708 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_129
timestamp 1605641404
transform 1 0 12972 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1605641404
transform 1 0 16284 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_146
timestamp 1605641404
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1605641404
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1605641404
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 17112 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1605641404
transform 1 0 16744 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_168
timestamp 1605641404
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_173
timestamp 1605641404
transform 1 0 17020 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 19136 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp 1605641404
transform 1 0 18584 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1605641404
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1605641404
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1605641404
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1605641404
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1605641404
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1605641404
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1605641404
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1605641404
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1605641404
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9108 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_86
timestamp 1605641404
transform 1 0 9016 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1605641404
transform 1 0 10580 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1605641404
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_123
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1605641404
transform 1 0 12696 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1605641404
transform 1 0 14168 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13156 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_129
timestamp 1605641404
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_140
timestamp 1605641404
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 15272 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_9_151
timestamp 1605641404
transform 1 0 14996 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 16928 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_170
timestamp 1605641404
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1605641404
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1605641404
transform 1 0 19044 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1605641404
transform 1 0 20056 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1605641404
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_204
timestamp 1605641404
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1605641404
transform 1 0 20884 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1605641404
transform 1 0 21252 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1605641404
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1605641404
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1605641404
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1605641404
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1605641404
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1605641404
transform 1 0 8464 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 8832 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10120 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1605641404
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_97
timestamp 1605641404
transform 1 0 10028 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 11132 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1605641404
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_125
timestamp 1605641404
transform 1 0 12604 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13524 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_133
timestamp 1605641404
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 15640 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1605641404
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16652 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_167
timestamp 1605641404
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1605641404
transform 1 0 18124 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18860 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1605641404
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1605641404
transform 1 0 20332 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1605641404
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_218
timestamp 1605641404
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1605641404
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1605641404
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1605641404
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1605641404
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1605641404
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8556 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_74
timestamp 1605641404
transform 1 0 7912 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_80
timestamp 1605641404
transform 1 0 8464 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_90
timestamp 1605641404
transform 1 0 9384 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 12604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_109
timestamp 1605641404
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1605641404
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14168 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13156 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_128
timestamp 1605641404
transform 1 0 12880 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_140
timestamp 1605641404
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15548 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 15180 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_151
timestamp 1605641404
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_156
timestamp 1605641404
transform 1 0 15456 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1605641404
transform 1 0 17204 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1605641404
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_173
timestamp 1605641404
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1605641404
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1605641404
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19504 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_193
timestamp 1605641404
transform 1 0 18860 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_199
timestamp 1605641404
transform 1 0 19412 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_209
timestamp 1605641404
transform 1 0 20332 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_217
timestamp 1605641404
transform 1 0 21068 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1605641404
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1605641404
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1605641404
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1605641404
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1605641404
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_80
timestamp 1605641404
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10672 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1605641404
transform 1 0 10396 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1605641404
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1605641404
transform 1 0 11684 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_113
timestamp 1605641404
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_124
timestamp 1605641404
transform 1 0 12512 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12788 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_143
timestamp 1605641404
transform 1 0 14260 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1605641404
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_163
timestamp 1605641404
transform 1 0 16100 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 17020 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1605641404
transform 1 0 16744 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_169
timestamp 1605641404
transform 1 0 16652 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18676 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp 1605641404
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_207
timestamp 1605641404
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1605641404
transform 1 0 20332 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1605641404
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1605641404
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1605641404
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1605641404
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1605641404
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1605641404
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1605641404
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1605641404
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1605641404
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1605641404
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1605641404
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1605641404
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7636 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8004 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_13_74
timestamp 1605641404
transform 1 0 7912 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_68
timestamp 1605641404
transform 1 0 7360 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9752 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10396 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_91
timestamp 1605641404
transform 1 0 9476 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1605641404
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1605641404
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_96
timestamp 1605641404
transform 1 0 9936 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_100
timestamp 1605641404
transform 1 0 10304 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1605641404
transform 1 0 11408 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12328 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1605641404
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_115
timestamp 1605641404
transform 1 0 11684 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1605641404
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1605641404
transform 1 0 11868 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1605641404
transform 1 0 12236 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 13340 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 14352 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_139
timestamp 1605641404
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_144
timestamp 1605641404
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_131
timestamp 1605641404
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_142
timestamp 1605641404
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1605641404
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14536 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16192 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16376 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1605641404
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1605641404
transform 1 0 17112 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18124 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1605641404
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_173
timestamp 1605641404
transform 1 0 17020 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1605641404
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_172
timestamp 1605641404
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_183
timestamp 1605641404
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 19136 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1605641404
transform 1 0 19964 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19044 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1605641404
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_201
timestamp 1605641404
transform 1 0 19596 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1605641404
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1605641404
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_214
timestamp 1605641404
transform 1 0 20792 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1605641404
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1605641404
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1605641404
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1605641404
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1605641404
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1605641404
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1605641404
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1605641404
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8464 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_15_74
timestamp 1605641404
transform 1 0 7912 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 9476 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 10580 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1605641404
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_97
timestamp 1605641404
transform 1 0 10028 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11592 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_112
timestamp 1605641404
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1605641404
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14260 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13248 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1605641404
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 16284 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_152
timestamp 1605641404
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1605641404
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1605641404
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1605641404
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1605641404
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_187
timestamp 1605641404
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 19596 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1605641404
transform 1 0 18584 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_199
timestamp 1605641404
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_217
timestamp 1605641404
transform 1 0 21068 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1605641404
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1605641404
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1605641404
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1605641404
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7360 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1605641404
transform 1 0 9016 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9752 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1605641404
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_89
timestamp 1605641404
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_103
timestamp 1605641404
transform 1 0 10580 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1605641404
transform 1 0 12420 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10764 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp 1605641404
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 13064 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_16_126
timestamp 1605641404
transform 1 0 12696 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15548 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1605641404
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1605641404
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16560 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_184
timestamp 1605641404
transform 1 0 18032 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1605641404
transform 1 0 18768 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19780 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1605641404
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1605641404
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1605641404
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1605641404
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1605641404
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1605641404
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1605641404
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1605641404
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1605641404
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1605641404
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8280 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_74
timestamp 1605641404
transform 1 0 7912 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10212 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 9292 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1605641404
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_95
timestamp 1605641404
transform 1 0 9844 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 11316 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_108
timestamp 1605641404
transform 1 0 11040 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1605641404
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13892 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1605641404
transform 1 0 15364 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_148
timestamp 1605641404
transform 1 0 14720 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_154
timestamp 1605641404
transform 1 0 15272 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_164
timestamp 1605641404
transform 1 0 16192 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1605641404
transform 1 0 18124 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1605641404
transform 1 0 16836 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1605641404
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_170
timestamp 1605641404
transform 1 0 16744 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1605641404
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1605641404
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 19688 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1605641404
transform 1 0 18676 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_189
timestamp 1605641404
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1605641404
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1605641404
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1605641404
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1605641404
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1605641404
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1605641404
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7452 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_68
timestamp 1605641404
transform 1 0 7360 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1605641404
transform 1 0 9108 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1605641404
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1605641404
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 11408 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_109
timestamp 1605641404
transform 1 0 11132 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13432 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_128
timestamp 1605641404
transform 1 0 12880 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15732 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1605641404
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1605641404
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1605641404
transform 1 0 17388 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_175
timestamp 1605641404
transform 1 0 17204 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1605641404
transform 1 0 18216 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1605641404
transform 1 0 20240 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 18584 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1605641404
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1605641404
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1605641404
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1605641404
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_218
timestamp 1605641404
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1605641404
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1605641404
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1605641404
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1605641404
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1605641404
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1605641404
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1605641404
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1605641404
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1605641404
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1605641404
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1605641404
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1605641404
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9384 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9752 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1605641404
transform 1 0 9108 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_86
timestamp 1605641404
transform 1 0 9016 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_103
timestamp 1605641404
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10764 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11040 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11960 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_106
timestamp 1605641404
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_117
timestamp 1605641404
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_114
timestamp 1605641404
transform 1 0 11592 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 14352 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 13156 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 13340 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_129
timestamp 1605641404
transform 1 0 12972 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_142
timestamp 1605641404
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_127
timestamp 1605641404
transform 1 0 12788 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_140
timestamp 1605641404
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 15732 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1605641404
transform 1 0 16192 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_160
timestamp 1605641404
transform 1 0 15824 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1605641404
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_157
timestamp 1605641404
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_168
timestamp 1605641404
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1605641404
transform 1 0 16468 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 16744 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 16560 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp 1605641404
transform 1 0 17572 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_184
timestamp 1605641404
transform 1 0 18032 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_177
timestamp 1605641404
transform 1 0 17388 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1605641404
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 17756 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1605641404
transform 1 0 18124 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18676 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18768 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1605641404
transform 1 0 19780 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_189
timestamp 1605641404
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1605641404
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1605641404
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_201
timestamp 1605641404
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1605641404
transform 1 0 20332 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1605641404
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_218
timestamp 1605641404
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1605641404
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1605641404
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1605641404
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1605641404
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1605641404
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1605641404
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1605641404
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1605641404
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1605641404
transform 1 0 8740 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_74
timestamp 1605641404
transform 1 0 7912 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_82
timestamp 1605641404
transform 1 0 8648 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9200 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_86
timestamp 1605641404
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_104
timestamp 1605641404
transform 1 0 10672 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 11316 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_110
timestamp 1605641404
transform 1 0 11224 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1605641404
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_123
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1605641404
transform 1 0 13708 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12696 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_135
timestamp 1605641404
transform 1 0 13524 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16192 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14904 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 15916 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_146
timestamp 1605641404
transform 1 0 14536 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_159
timestamp 1605641404
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1605641404
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_180
timestamp 1605641404
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1605641404
transform 1 0 19688 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_193
timestamp 1605641404
transform 1 0 18860 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_201
timestamp 1605641404
transform 1 0 19596 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1605641404
transform 1 0 20700 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1605641404
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_217
timestamp 1605641404
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1605641404
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1605641404
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1605641404
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1605641404
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_62
timestamp 1605641404
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6900 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_79
timestamp 1605641404
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1605641404
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1605641404
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_102
timestamp 1605641404
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 11040 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 10764 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_124
timestamp 1605641404
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12696 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14352 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_142
timestamp 1605641404
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 16284 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_150
timestamp 1605641404
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_163
timestamp 1605641404
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1605641404
transform 1 0 17940 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_181
timestamp 1605641404
transform 1 0 17756 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_186
timestamp 1605641404
transform 1 0 18216 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1605641404
transform 1 0 20240 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18584 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1605641404
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1605641404
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1605641404
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1605641404
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1605641404
transform 1 0 21160 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1605641404
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1605641404
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1605641404
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_39
timestamp 1605641404
transform 1 0 4692 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1605641404
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_47
timestamp 1605641404
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1605641404
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_62
timestamp 1605641404
transform 1 0 6808 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7728 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_70
timestamp 1605641404
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 10580 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9384 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_88
timestamp 1605641404
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_99
timestamp 1605641404
transform 1 0 10212 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1605641404
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_109
timestamp 1605641404
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1605641404
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13616 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_132
timestamp 1605641404
transform 1 0 13248 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1605641404
transform 1 0 15364 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_23_152
timestamp 1605641404
transform 1 0 15088 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_164
timestamp 1605641404
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1605641404
transform 1 0 17388 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1605641404
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1605641404
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1605641404
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1605641404
transform 1 0 18032 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18400 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19412 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_197
timestamp 1605641404
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_208
timestamp 1605641404
transform 1 0 20240 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20424 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_216
timestamp 1605641404
transform 1 0 20976 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1605641404
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1605641404
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1605641404
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1605641404
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1605641404
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6440 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1605641404
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_56
timestamp 1605641404
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_74
timestamp 1605641404
transform 1 0 7912 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10672 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 9660 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1605641404
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_86
timestamp 1605641404
transform 1 0 9016 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_99
timestamp 1605641404
transform 1 0 10212 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_103
timestamp 1605641404
transform 1 0 10580 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11684 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_113
timestamp 1605641404
transform 1 0 11500 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_124
timestamp 1605641404
transform 1 0 12512 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 13524 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12788 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1605641404
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1605641404
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1605641404
transform 1 0 16284 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1605641404
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_163
timestamp 1605641404
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16560 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_184
timestamp 1605641404
transform 1 0 18032 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18400 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20056 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_204
timestamp 1605641404
transform 1 0 19872 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1605641404
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1605641404
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1605641404
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1605641404
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1605641404
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1605641404
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1605641404
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1605641404
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1605641404
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1605641404
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1605641404
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1605641404
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 8648 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_78
timestamp 1605641404
transform 1 0 8280 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9476 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_88
timestamp 1605641404
transform 1 0 9200 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11132 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1605641404
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_107
timestamp 1605641404
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1605641404
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14168 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_139
timestamp 1605641404
transform 1 0 13892 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1605641404
transform 1 0 15824 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_158
timestamp 1605641404
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18032 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16836 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1605641404
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1605641404
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1605641404
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19688 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1605641404
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1605641404
transform 1 0 20700 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1605641404
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_211
timestamp 1605641404
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_217
timestamp 1605641404
transform 1 0 21068 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1605641404
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1605641404
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1605641404
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1605641404
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1605641404
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1605641404
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1605641404
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1605641404
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1605641404
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1605641404
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1605641404
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1605641404
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1605641404
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1605641404
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_56
timestamp 1605641404
transform 1 0 6256 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1605641404
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1605641404
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1605641404
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6992 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6992 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8096 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1605641404
transform 1 0 8648 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_26_73
timestamp 1605641404
transform 1 0 7820 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_80
timestamp 1605641404
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1605641404
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1605641404
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1605641404
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1605641404
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1605641404
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9660 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1605641404
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_102
timestamp 1605641404
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1605641404
transform 1 0 10028 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1605641404
transform 1 0 10120 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10672 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10396 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1605641404
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12512 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1605641404
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_117
timestamp 1605641404
transform 1 0 11868 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1605641404
transform 1 0 11500 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1605641404
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1605641404
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1605641404
transform 1 0 13524 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1605641404
transform 1 0 13064 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_128
timestamp 1605641404
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_139
timestamp 1605641404
transform 1 0 13892 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_133
timestamp 1605641404
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_144
timestamp 1605641404
transform 1 0 14352 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_152
timestamp 1605641404
transform 1 0 15088 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_154
timestamp 1605641404
transform 1 0 15272 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1605641404
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1605641404
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15364 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15364 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_164
timestamp 1605641404
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_164
timestamp 1605641404
transform 1 0 16192 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1605641404
transform 1 0 16376 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1605641404
transform 1 0 16376 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1605641404
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1605641404
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1605641404
transform 1 0 17296 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_170
timestamp 1605641404
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1605641404
transform 1 0 16928 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1605641404
transform 1 0 16836 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1605641404
transform 1 0 17388 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1605641404
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_184
timestamp 1605641404
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1605641404
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18216 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17480 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18032 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1605641404
transform 1 0 20240 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1605641404
transform 1 0 19228 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19780 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_195
timestamp 1605641404
transform 1 0 19044 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1605641404
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_200
timestamp 1605641404
transform 1 0 19504 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1605641404
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20516 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1605641404
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1605641404
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1605641404
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1605641404
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_218
timestamp 1605641404
transform 1 0 21160 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1605641404
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_217
timestamp 1605641404
transform 1 0 21068 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1605641404
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1605641404
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1605641404
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1605641404
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1605641404
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1605641404
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1605641404
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1605641404
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7360 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10212 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1605641404
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1605641404
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_93
timestamp 1605641404
transform 1 0 9660 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11960 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11224 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_108
timestamp 1605641404
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_116
timestamp 1605641404
transform 1 0 11776 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_124
timestamp 1605641404
transform 1 0 12512 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12972 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13984 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_128
timestamp 1605641404
transform 1 0 12880 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1605641404
transform 1 0 13800 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1605641404
transform 1 0 14720 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15456 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1605641404
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_146
timestamp 1605641404
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1605641404
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_154
timestamp 1605641404
transform 1 0 15272 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_165
timestamp 1605641404
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1605641404
transform 1 0 16468 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16928 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_170
timestamp 1605641404
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1605641404
transform 1 0 18584 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19688 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_188
timestamp 1605641404
transform 1 0 18400 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_199
timestamp 1605641404
transform 1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_208
timestamp 1605641404
transform 1 0 20240 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1605641404
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1605641404
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1605641404
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1605641404
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1605641404
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1605641404
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1605641404
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1605641404
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1605641404
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1605641404
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1605641404
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1605641404
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1605641404
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_74
timestamp 1605641404
transform 1 0 7912 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_82
timestamp 1605641404
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8832 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9844 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_93
timestamp 1605641404
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_104
timestamp 1605641404
transform 1 0 10672 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11224 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1605641404
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_116
timestamp 1605641404
transform 1 0 11776 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_123
timestamp 1605641404
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13708 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12696 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_135
timestamp 1605641404
transform 1 0 13524 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15364 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_153
timestamp 1605641404
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1605641404
transform 1 0 17388 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1605641404
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_171
timestamp 1605641404
transform 1 0 16836 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1605641404
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1605641404
transform 1 0 19228 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19780 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1605641404
transform 1 0 18860 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_201
timestamp 1605641404
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1605641404
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1605641404
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1605641404
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1605641404
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1605641404
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1605641404
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1605641404
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1605641404
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1605641404
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1605641404
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1605641404
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1605641404
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1605641404
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7636 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_30_68
timestamp 1605641404
transform 1 0 7360 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1605641404
transform 1 0 10120 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10580 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1605641404
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_87
timestamp 1605641404
transform 1 0 9108 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1605641404
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_93
timestamp 1605641404
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_97
timestamp 1605641404
transform 1 0 10028 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_101
timestamp 1605641404
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12604 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_30_119
timestamp 1605641404
transform 1 0 12052 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1605641404
transform 1 0 14076 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1605641404
transform 1 0 15456 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1605641404
transform 1 0 14628 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16008 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1605641404
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1605641404
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1605641404
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_160
timestamp 1605641404
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1605641404
transform 1 0 17664 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_178
timestamp 1605641404
transform 1 0 17480 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19596 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18860 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_189
timestamp 1605641404
transform 1 0 18492 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_199
timestamp 1605641404
transform 1 0 19412 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_207
timestamp 1605641404
transform 1 0 20148 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1605641404
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1605641404
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1605641404
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1605641404
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1605641404
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1605641404
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1605641404
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1605641404
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1605641404
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1605641404
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1605641404
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1605641404
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1605641404
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1605641404
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8372 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_74
timestamp 1605641404
transform 1 0 7912 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_78
timestamp 1605641404
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 10028 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_95
timestamp 1605641404
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1605641404
transform 1 0 11684 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1605641404
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1605641404
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1605641404
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1605641404
transform 1 0 14076 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1605641404
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1605641404
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1605641404
transform 1 0 15732 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1605641404
transform 1 0 15180 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1605641404
transform 1 0 14628 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_151
timestamp 1605641404
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_157
timestamp 1605641404
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1605641404
transform 1 0 16100 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1605641404
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1605641404
transform 1 0 16468 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17112 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1605641404
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_171
timestamp 1605641404
transform 1 0 16836 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1605641404
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1605641404
transform 1 0 18860 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1605641404
transform 1 0 19412 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1605641404
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_188
timestamp 1605641404
transform 1 0 18400 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_192
timestamp 1605641404
transform 1 0 18768 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1605641404
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1605641404
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1605641404
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1605641404
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1605641404
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1605641404
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1605641404
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1605641404
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1605641404
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1605641404
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1605641404
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1605641404
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1605641404
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1605641404
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1605641404
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1605641404
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8648 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1605641404
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_75
timestamp 1605641404
transform 1 0 8004 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_81
timestamp 1605641404
transform 1 0 8556 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9752 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1605641404
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_91
timestamp 1605641404
transform 1 0 9476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_103
timestamp 1605641404
transform 1 0 10580 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1605641404
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11500 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1605641404
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_111
timestamp 1605641404
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1605641404
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1605641404
transform 1 0 13800 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1605641404
transform 1 0 14352 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1605641404
transform 1 0 13156 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_129
timestamp 1605641404
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_135
timestamp 1605641404
transform 1 0 13524 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_142
timestamp 1605641404
transform 1 0 14168 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1605641404
transform 1 0 15548 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1605641404
transform 1 0 16100 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1605641404
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_148
timestamp 1605641404
transform 1 0 14720 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1605641404
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_156
timestamp 1605641404
transform 1 0 15456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_161
timestamp 1605641404
transform 1 0 15916 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1605641404
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1605641404
transform 1 0 17204 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1605641404
transform 1 0 16652 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1605641404
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_167
timestamp 1605641404
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1605641404
transform 1 0 17020 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_179
timestamp 1605641404
transform 1 0 17572 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_185
timestamp 1605641404
transform 1 0 18124 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1605641404
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1605641404
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1605641404
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp 1605641404
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1605641404
transform 1 0 19228 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1605641404
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1605641404
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1605641404
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1605641404
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1605641404
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1605641404
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1605641404
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal3 s 0 5720 480 5840 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 17144 480 17264 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 22320 3816 22800 3936 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 22320 8440 22800 8560 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 22320 8984 22800 9104 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 22320 9392 22800 9512 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 22320 9936 22800 10056 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 22320 10344 22800 10464 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 22320 10752 22800 10872 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 22320 11296 22800 11416 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 22320 11704 22800 11824 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 22320 12248 22800 12368 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 22320 12656 22800 12776 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 22320 4224 22800 4344 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 22320 4768 22800 4888 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 22320 5176 22800 5296 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 22320 6128 22800 6248 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 22320 6672 22800 6792 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 22320 7080 22800 7200 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 22320 7488 22800 7608 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 22320 8032 22800 8152 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 22320 13200 22800 13320 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 22320 17824 22800 17944 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 22320 18776 22800 18896 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 22320 19184 22800 19304 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 22320 13608 22800 13728 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 22320 14016 22800 14136 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 22320 14560 22800 14680 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 22320 14968 22800 15088 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 22320 15512 22800 15632 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 22320 15920 22800 16040 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 22320 16464 22800 16584 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 22320 16872 22800 16992 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 22320 17280 22800 17400 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 846 0 902 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 7470 0 7526 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 8022 0 8078 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 9678 0 9734 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 10230 0 10286 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 1950 0 2006 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2502 0 2558 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3054 0 3110 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 3606 0 3662 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 17498 0 17554 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 22466 0 22522 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 14738 0 14794 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 15290 0 15346 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 16394 0 16450 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal2 s 846 22320 902 22800 6 chany_top_in[0]
port 83 nsew default input
rlabel metal2 s 6366 22320 6422 22800 6 chany_top_in[10]
port 84 nsew default input
rlabel metal2 s 6918 22320 6974 22800 6 chany_top_in[11]
port 85 nsew default input
rlabel metal2 s 7470 22320 7526 22800 6 chany_top_in[12]
port 86 nsew default input
rlabel metal2 s 8022 22320 8078 22800 6 chany_top_in[13]
port 87 nsew default input
rlabel metal2 s 8574 22320 8630 22800 6 chany_top_in[14]
port 88 nsew default input
rlabel metal2 s 9126 22320 9182 22800 6 chany_top_in[15]
port 89 nsew default input
rlabel metal2 s 9678 22320 9734 22800 6 chany_top_in[16]
port 90 nsew default input
rlabel metal2 s 10230 22320 10286 22800 6 chany_top_in[17]
port 91 nsew default input
rlabel metal2 s 10782 22320 10838 22800 6 chany_top_in[18]
port 92 nsew default input
rlabel metal2 s 11334 22320 11390 22800 6 chany_top_in[19]
port 93 nsew default input
rlabel metal2 s 1398 22320 1454 22800 6 chany_top_in[1]
port 94 nsew default input
rlabel metal2 s 1950 22320 2006 22800 6 chany_top_in[2]
port 95 nsew default input
rlabel metal2 s 2502 22320 2558 22800 6 chany_top_in[3]
port 96 nsew default input
rlabel metal2 s 3054 22320 3110 22800 6 chany_top_in[4]
port 97 nsew default input
rlabel metal2 s 3606 22320 3662 22800 6 chany_top_in[5]
port 98 nsew default input
rlabel metal2 s 4158 22320 4214 22800 6 chany_top_in[6]
port 99 nsew default input
rlabel metal2 s 4710 22320 4766 22800 6 chany_top_in[7]
port 100 nsew default input
rlabel metal2 s 5262 22320 5318 22800 6 chany_top_in[8]
port 101 nsew default input
rlabel metal2 s 5814 22320 5870 22800 6 chany_top_in[9]
port 102 nsew default input
rlabel metal2 s 11978 22320 12034 22800 6 chany_top_out[0]
port 103 nsew default tristate
rlabel metal2 s 17498 22320 17554 22800 6 chany_top_out[10]
port 104 nsew default tristate
rlabel metal2 s 18050 22320 18106 22800 6 chany_top_out[11]
port 105 nsew default tristate
rlabel metal2 s 18602 22320 18658 22800 6 chany_top_out[12]
port 106 nsew default tristate
rlabel metal2 s 19154 22320 19210 22800 6 chany_top_out[13]
port 107 nsew default tristate
rlabel metal2 s 19706 22320 19762 22800 6 chany_top_out[14]
port 108 nsew default tristate
rlabel metal2 s 20258 22320 20314 22800 6 chany_top_out[15]
port 109 nsew default tristate
rlabel metal2 s 20810 22320 20866 22800 6 chany_top_out[16]
port 110 nsew default tristate
rlabel metal2 s 21362 22320 21418 22800 6 chany_top_out[17]
port 111 nsew default tristate
rlabel metal2 s 21914 22320 21970 22800 6 chany_top_out[18]
port 112 nsew default tristate
rlabel metal2 s 22466 22320 22522 22800 6 chany_top_out[19]
port 113 nsew default tristate
rlabel metal2 s 12530 22320 12586 22800 6 chany_top_out[1]
port 114 nsew default tristate
rlabel metal2 s 13082 22320 13138 22800 6 chany_top_out[2]
port 115 nsew default tristate
rlabel metal2 s 13634 22320 13690 22800 6 chany_top_out[3]
port 116 nsew default tristate
rlabel metal2 s 14186 22320 14242 22800 6 chany_top_out[4]
port 117 nsew default tristate
rlabel metal2 s 14738 22320 14794 22800 6 chany_top_out[5]
port 118 nsew default tristate
rlabel metal2 s 15290 22320 15346 22800 6 chany_top_out[6]
port 119 nsew default tristate
rlabel metal2 s 15842 22320 15898 22800 6 chany_top_out[7]
port 120 nsew default tristate
rlabel metal2 s 16394 22320 16450 22800 6 chany_top_out[8]
port 121 nsew default tristate
rlabel metal2 s 16946 22320 17002 22800 6 chany_top_out[9]
port 122 nsew default tristate
rlabel metal3 s 22320 22448 22800 22568 6 prog_clk
port 123 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_34_
port 124 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_35_
port 125 nsew default input
rlabel metal3 s 22320 960 22800 1080 6 right_bottom_grid_pin_36_
port 126 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_37_
port 127 nsew default input
rlabel metal3 s 22320 1912 22800 2032 6 right_bottom_grid_pin_38_
port 128 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_39_
port 129 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_40_
port 130 nsew default input
rlabel metal3 s 22320 3408 22800 3528 6 right_bottom_grid_pin_41_
port 131 nsew default input
rlabel metal2 s 294 22320 350 22800 6 top_left_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 133 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
