* NGSPICE file created from cbx_1__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

.subckt cbx_1__2_ IO_ISOL_N SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP bottom_grid_pin_0_
+ bottom_grid_pin_10_ bottom_grid_pin_11_ bottom_grid_pin_12_ bottom_grid_pin_13_
+ bottom_grid_pin_14_ bottom_grid_pin_15_ bottom_grid_pin_1_ bottom_grid_pin_2_ bottom_grid_pin_3_
+ bottom_grid_pin_4_ bottom_grid_pin_5_ bottom_grid_pin_6_ bottom_grid_pin_7_ bottom_grid_pin_8_
+ bottom_grid_pin_9_ bottom_width_0_height_0__pin_0_ bottom_width_0_height_0__pin_1_lower
+ bottom_width_0_height_0__pin_1_upper ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_IN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
+ prog_clk_0_S_in prog_clk_0_W_out top_grid_pin_0_ VPWR VGND
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_7.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_13.mux_l3_in_0_ mux_top_ipin_13.mux_l2_in_1_/X mux_top_ipin_13.mux_l2_in_0_/X
+ mux_top_ipin_13.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_13.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_66_ chanx_left_in[10] VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_6.mux_l1_in_0_/X mux_top_ipin_6.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
X_49_ chanx_right_in[7] VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_13.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_top_ipin_13.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_65_ chanx_left_in[11] VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_48_ chanx_right_in[8] VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_13.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_13.mux_l1_in_0_/X mux_top_ipin_13.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_6.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_bottom_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_64_ chanx_left_in[12] VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_4.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_4_ sky130_fd_sc_hd__buf_4
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_47_ chanx_right_in[9] VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_13.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_bottom_ipin_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_63_ chanx_left_in[13] VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
Xprog_clk_0_FTB00 prog_clk_0_S_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_46_ chanx_right_in[10] VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_29_ VGND VGND VPWR VPWR _29_/HI _29_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_11.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_11_ sky130_fd_sc_hd__buf_4
Xmux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_0.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR top_grid_pin_0_ sky130_fd_sc_hd__buf_4
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_bottom_ipin_0.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_2.mux_l2_in_3_ _30_/HI chanx_right_in[15] mux_top_ipin_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_62_ chanx_left_in[14] VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_45_ chanx_right_in[11] VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_2.mux_l4_in_0_ mux_top_ipin_2.mux_l3_in_1_/X mux_top_ipin_2.mux_l3_in_0_/X
+ mux_top_ipin_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_28_ VGND VGND VPWR VPWR _28_/HI _28_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_7.mux_l2_in_3_ _18_/HI chanx_right_in[18] mux_top_ipin_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_2.mux_l3_in_1_ mux_top_ipin_2.mux_l2_in_3_/X mux_top_ipin_2.mux_l2_in_2_/X
+ mux_top_ipin_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ ccff_head VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_2.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[7] mux_top_ipin_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_7.mux_l4_in_0_ mux_top_ipin_7.mux_l3_in_1_/X mux_top_ipin_7.mux_l3_in_0_/X
+ mux_top_ipin_7.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_61_ chanx_left_in[15] VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_7.mux_l3_in_1_ mux_top_ipin_7.mux_l2_in_3_/X mux_top_ipin_7.mux_l2_in_2_/X
+ mux_top_ipin_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_44_ chanx_right_in[12] VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
XFILLER_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27_ VGND VGND VPWR VPWR _27_/HI _27_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_7.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_top_ipin_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_2.mux_l3_in_0_ mux_top_ipin_2.mux_l2_in_1_/X mux_top_ipin_2.mux_l2_in_0_/X
+ mux_top_ipin_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_14.mux_l2_in_3_ _28_/HI chanx_right_in[19] mux_top_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_4_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_2.mux_l2_in_1_ chanx_left_in[7] chanx_right_in[3] mux_top_ipin_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_14.mux_l4_in_0_ mux_top_ipin_14.mux_l3_in_1_/X mux_top_ipin_14.mux_l3_in_0_/X
+ mux_top_ipin_14.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_14.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_60_ chanx_left_in[16] VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_7.mux_l3_in_0_ mux_top_ipin_7.mux_l2_in_1_/X mux_top_ipin_7.mux_l2_in_0_/X
+ mux_top_ipin_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_43_ chanx_right_in[13] VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_7.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_7_ sky130_fd_sc_hd__buf_4
Xmux_top_ipin_14.mux_l3_in_1_ mux_top_ipin_14.mux_l2_in_3_/X mux_top_ipin_14.mux_l2_in_2_/X
+ mux_top_ipin_14.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_14.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_7.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_7.mux_l1_in_2_/X mux_top_ipin_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26_ VGND VGND VPWR VPWR _26_/HI _26_/LO sky130_fd_sc_hd__conb_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_14.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[11] mux_top_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_7.mux_l1_in_2_ chanx_right_in[8] chanx_left_in[8] mux_top_ipin_7.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_2.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_2.mux_l1_in_0_/X mux_top_ipin_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XFILLER_4_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_42_ chanx_right_in[14] VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_14.mux_l3_in_0_ mux_top_ipin_14.mux_l2_in_1_/X mux_top_ipin_14.mux_l2_in_0_/X
+ mux_top_ipin_14.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_14.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_11.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_11.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_7.mux_l2_in_0_ mux_top_ipin_7.mux_l1_in_1_/X mux_top_ipin_7.mux_l1_in_0_/X
+ mux_top_ipin_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_25_ VGND VGND VPWR VPWR _25_/HI _25_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_14.mux_l2_in_1_ chanx_left_in[11] chanx_right_in[3] mux_top_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_14.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_14_ sky130_fd_sc_hd__buf_4
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_7.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_7.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_top_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_14.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_14.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_1.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_2.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_41_ chanx_right_in[15] VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_11.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_11.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24_ VGND VGND VPWR VPWR _24_/HI _24_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_14.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_14.mux_l1_in_0_/X mux_top_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_0_ sky130_fd_sc_hd__buf_4
XFILLER_21_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_7.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_7.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_top_ipin_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_14.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_14.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_1.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_40_ chanx_right_in[16] VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_11.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_11.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
X_23_ VGND VGND VPWR VPWR _23_/HI _23_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_top_ipin_4.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_14.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_14.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_14.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_22_ VGND VGND VPWR VPWR _22_/HI _22_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_10.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_11.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_7.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN
+ logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR bottom_width_0_height_0__pin_1_lower sky130_fd_sc_hd__ebufn_4
XFILLER_21_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_top_ipin_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_13.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_14.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_3.mux_l2_in_3_ _31_/HI chanx_right_in[14] mux_top_ipin_3.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21_ VGND VGND VPWR VPWR _21_/HI _21_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_6.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_3.mux_l4_in_0_ mux_top_ipin_3.mux_l3_in_1_/X mux_top_ipin_3.mux_l3_in_0_/X
+ mux_top_ipin_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_8.mux_l2_in_3_ _19_/HI chanx_right_in[19] mux_top_ipin_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l3_in_1_ mux_top_ipin_3.mux_l2_in_3_/X mux_top_ipin_3.mux_l2_in_2_/X
+ mux_top_ipin_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_3.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[8] mux_top_ipin_3.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l4_in_0_ mux_top_ipin_8.mux_l3_in_1_/X mux_top_ipin_8.mux_l3_in_0_/X
+ mux_top_ipin_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_10.mux_l2_in_3_ _24_/HI chanx_right_in[15] mux_top_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20_ VGND VGND VPWR VPWR _20_/HI _20_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_8.mux_l3_in_1_ mux_top_ipin_8.mux_l2_in_3_/X mux_top_ipin_8.mux_l2_in_2_/X
+ mux_top_ipin_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_8.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[13] mux_top_ipin_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_3_ sky130_fd_sc_hd__buf_4
Xmux_top_ipin_10.mux_l4_in_0_ mux_top_ipin_10.mux_l3_in_1_/X mux_top_ipin_10.mux_l3_in_0_/X
+ mux_top_ipin_10.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_10.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_3.mux_l3_in_0_ mux_top_ipin_3.mux_l2_in_1_/X mux_top_ipin_3.mux_l2_in_0_/X
+ mux_top_ipin_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_15.mux_l2_in_3_ _29_/HI chanx_right_in[16] mux_top_ipin_15.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_10.mux_l3_in_1_ mux_top_ipin_10.mux_l2_in_3_/X mux_top_ipin_10.mux_l2_in_2_/X
+ mux_top_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_10.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_3.mux_l2_in_1_ chanx_left_in[8] mux_top_ipin_3.mux_l1_in_2_/X mux_top_ipin_3.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[7] mux_top_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_15.mux_l4_in_0_ mux_top_ipin_15.mux_l3_in_1_/X mux_top_ipin_15.mux_l3_in_0_/X
+ mux_top_ipin_15.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_15.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l3_in_0_ mux_top_ipin_8.mux_l2_in_1_/X mux_top_ipin_8.mux_l2_in_0_/X
+ mux_top_ipin_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_15.mux_l3_in_1_ mux_top_ipin_15.mux_l2_in_3_/X mux_top_ipin_15.mux_l2_in_2_/X
+ mux_top_ipin_15.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_15.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_8.mux_l2_in_1_ chanx_left_in[13] mux_top_ipin_8.mux_l1_in_2_/X mux_top_ipin_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_15.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_15.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l1_in_2_ chanx_right_in[9] chanx_left_in[9] mux_top_ipin_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_10.mux_l3_in_0_ mux_top_ipin_10.mux_l2_in_1_/X mux_top_ipin_10.mux_l2_in_0_/X
+ mux_top_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_10.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l2_in_0_ mux_top_ipin_3.mux_l1_in_1_/X mux_top_ipin_3.mux_l1_in_0_/X
+ mux_top_ipin_3.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_10.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_10_ sky130_fd_sc_hd__buf_4
XFILLER_1_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_10.mux_l2_in_1_ chanx_left_in[7] chanx_right_in[3] mux_top_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_15.mux_l3_in_0_ mux_top_ipin_15.mux_l2_in_1_/X mux_top_ipin_15.mux_l2_in_0_/X
+ mux_top_ipin_15.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_15.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_8.mux_l2_in_0_ mux_top_ipin_8.mux_l1_in_1_/X mux_top_ipin_8.mux_l1_in_0_/X
+ mux_top_ipin_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_15.mux_l1_in_2_/X mux_top_ipin_15.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_8.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_10.mux_l1_in_0_/X mux_top_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_3.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_15.mux_l2_in_0_ mux_top_ipin_15.mux_l1_in_1_/X mux_top_ipin_15.mux_l1_in_0_/X
+ mux_top_ipin_15.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_15.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_/CLK sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_8.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_15.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_76_ chanx_left_in[0] VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_10.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_59_ chanx_left_in[17] VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_6.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_6_ sky130_fd_sc_hd__buf_4
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_15.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_15.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_75_ chanx_left_in[1] VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_58_ chanx_left_in[18] VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_13.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_13_ sky130_fd_sc_hd__buf_4
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_74_ chanx_left_in[2] VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_3_ _32_/HI chanx_right_in[15] mux_top_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_ipin_0.mux_l2_in_3_ _21_/HI chanx_right_in[16] mux_bottom_ipin_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_57_ chanx_left_in[19] VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE bottom_width_0_height_0__pin_0_
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
+ sky130_fd_sc_hd__ebufn_4
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_4.mux_l4_in_0_ mux_top_ipin_4.mux_l3_in_1_/X mux_top_ipin_4.mux_l3_in_0_/X
+ mux_top_ipin_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_ipin_0.mux_l4_in_0_ mux_bottom_ipin_0.mux_l3_in_1_/X mux_bottom_ipin_0.mux_l3_in_0_/X
+ mux_bottom_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_9.mux_l2_in_3_ _20_/HI chanx_right_in[14] mux_top_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_4.mux_l3_in_1_ mux_top_ipin_4.mux_l2_in_3_/X mux_top_ipin_4.mux_l2_in_2_/X
+ mux_top_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_10.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_0.mux_l3_in_1_ mux_bottom_ipin_0.mux_l2_in_3_/X mux_bottom_ipin_0.mux_l2_in_2_/X
+ mux_bottom_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_73_ chanx_left_in[3] VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[9] mux_top_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_9.mux_l4_in_0_ mux_top_ipin_9.mux_l3_in_1_/X mux_top_ipin_9.mux_l3_in_0_/X
+ mux_top_ipin_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xprog_clk_0_W_FTB01 prog_clk_0_S_in VGND VGND VPWR VPWR prog_clk_0_W_out sky130_fd_sc_hd__buf_4
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_bottom_ipin_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_11.mux_l2_in_3_ _25_/HI chanx_right_in[16] mux_top_ipin_11.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_56_ chanx_right_in[0] VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
X_39_ chanx_right_in[17] VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_9.mux_l3_in_1_ mux_top_ipin_9.mux_l2_in_3_/X mux_top_ipin_9.mux_l2_in_2_/X
+ mux_top_ipin_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_13.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_13.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_0.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_11.mux_l4_in_0_ mux_top_ipin_11.mux_l3_in_1_/X mux_top_ipin_11.mux_l3_in_0_/X
+ mux_top_ipin_11.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_11.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_9.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_top_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_10.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_10.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_4.mux_l3_in_0_ mux_top_ipin_4.mux_l2_in_1_/X mux_top_ipin_4.mux_l2_in_0_/X
+ mux_top_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_ipin_0.mux_l3_in_0_ mux_bottom_ipin_0.mux_l2_in_1_/X mux_bottom_ipin_0.mux_l2_in_0_/X
+ mux_bottom_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_11.mux_l3_in_1_ mux_top_ipin_11.mux_l2_in_3_/X mux_top_ipin_11.mux_l2_in_2_/X
+ mux_top_ipin_11.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_11.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_72_ chanx_left_in[4] VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_1_ chanx_left_in[9] mux_top_ipin_4.mux_l1_in_2_/X mux_top_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_bottom_ipin_0.mux_l1_in_2_/X
+ mux_bottom_ipin_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_55_ chanx_right_in[1] VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_3.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_11.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[12] mux_top_ipin_11.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_9.mux_l3_in_0_ mux_top_ipin_9.mux_l2_in_1_/X mux_top_ipin_9.mux_l2_in_0_/X
+ mux_top_ipin_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_4.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_38_ chanx_right_in[18] VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_13.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_13.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_bottom_ipin_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_9.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_9_ sky130_fd_sc_hd__buf_4
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_9.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ VGND VGND VPWR VPWR mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_9.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_top_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_10.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_10.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK sky130_fd_sc_hd__clkbuf_1
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_6.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_11.mux_l3_in_0_ mux_top_ipin_11.mux_l2_in_1_/X mux_top_ipin_11.mux_l2_in_0_/X
+ mux_top_ipin_11.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_11.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_71_ chanx_left_in[5] VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_0_ mux_top_ipin_4.mux_l1_in_1_/X mux_top_ipin_4.mux_l1_in_0_/X
+ mux_top_ipin_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_ipin_0.mux_l2_in_0_ mux_bottom_ipin_0.mux_l1_in_1_/X mux_bottom_ipin_0.mux_l1_in_0_/X
+ mux_bottom_ipin_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_3.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
X_54_ chanx_right_in[2] VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_11.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_11.mux_l1_in_2_/X mux_top_ipin_11.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_4.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_13.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_13.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_37_ chanx_right_in[19] VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
Xmux_bottom_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_bottom_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_11.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_top_ipin_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_9.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_9.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_9.mux_l1_in_0_/X mux_top_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_10.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_6.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_70_ chanx_left_in[6] VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_53_ chanx_right_in[3] VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_11.mux_l2_in_0_ mux_top_ipin_11.mux_l1_in_1_/X mux_top_ipin_11.mux_l1_in_0_/X
+ mux_top_ipin_11.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_11.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_4.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_12.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_13.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_36_ bottom_width_0_height_0__pin_1_lower VGND VGND VPWR VPWR bottom_width_0_height_0__pin_1_upper
+ sky130_fd_sc_hd__buf_2
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_11.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19_ VGND VGND VPWR VPWR _19_/HI _19_/LO sky130_fd_sc_hd__conb_1
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_9.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_9.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_2.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_2_ sky130_fd_sc_hd__buf_4
Xmux_top_ipin_9.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_52_ chanx_right_in[4] VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_35_ SC_IN_BOT VGND VGND VPWR VPWR SC_OUT_TOP sky130_fd_sc_hd__buf_2
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_/CLK mux_top_ipin_15.mux_l4_in_0_/S VGND
+ VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_11.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18_ VGND VGND VPWR VPWR _18_/HI _18_/LO sky130_fd_sc_hd__conb_1
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_top_ipin_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_9.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_51_ chanx_right_in[5] VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
X_34_ SC_IN_TOP VGND VGND VPWR VPWR SC_OUT_BOT sky130_fd_sc_hd__buf_2
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17_ VGND VGND VPWR VPWR _17_/HI _17_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l2_in_3_ _22_/HI chanx_right_in[17] mux_top_ipin_0.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_0.mux_l4_in_0_ mux_top_ipin_0.mux_l3_in_1_/X mux_top_ipin_0.mux_l3_in_0_/X
+ mux_top_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_50_ chanx_right_in[6] VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
XFILLER_11_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_5.mux_l2_in_3_ _33_/HI chanx_right_in[18] mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_33_ VGND VGND VPWR VPWR _33_/HI _33_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_0.mux_l3_in_1_ mux_top_ipin_0.mux_l2_in_3_/X mux_top_ipin_0.mux_l2_in_2_/X
+ mux_top_ipin_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_top_ipin_0.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.mux_l4_in_0_ mux_top_ipin_5.mux_l3_in_1_/X mux_top_ipin_5.mux_l3_in_0_/X
+ mux_top_ipin_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ VGND VGND VPWR VPWR mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_5.mux_l3_in_1_ mux_top_ipin_5.mux_l2_in_3_/X mux_top_ipin_5.mux_l2_in_2_/X
+ mux_top_ipin_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_5.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_32_ VGND VGND VPWR VPWR _32_/HI _32_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_0.mux_l3_in_0_ mux_top_ipin_0.mux_l2_in_1_/X mux_top_ipin_0.mux_l2_in_0_/X
+ mux_top_ipin_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_12.mux_l2_in_3_ _26_/HI chanx_right_in[17] mux_top_ipin_12.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_0.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_0.mux_l1_in_2_/X mux_top_ipin_0.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_12.mux_l4_in_0_ mux_top_ipin_12.mux_l3_in_1_/X mux_top_ipin_12.mux_l3_in_0_/X
+ mux_top_ipin_12.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_12.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_0.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.mux_l3_in_0_ mux_top_ipin_5.mux_l2_in_1_/X mux_top_ipin_5.mux_l2_in_0_/X
+ mux_top_ipin_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_5.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_5_ sky130_fd_sc_hd__buf_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_12.mux_l3_in_1_ mux_top_ipin_12.mux_l2_in_3_/X mux_top_ipin_12.mux_l2_in_2_/X
+ mux_top_ipin_12.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_12.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_5.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_31_ VGND VGND VPWR VPWR _31_/HI _31_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_12.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[13] mux_top_ipin_12.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l2_in_0_ mux_top_ipin_0.mux_l1_in_1_/X mux_top_ipin_0.mux_l1_in_0_/X
+ mux_top_ipin_0.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_12.mux_l3_in_0_ mux_top_ipin_12.mux_l2_in_1_/X mux_top_ipin_12.mux_l2_in_0_/X
+ mux_top_ipin_12.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_12.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_5.mux_l1_in_0_/X mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
X_30_ VGND VGND VPWR VPWR _30_/HI _30_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_12.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_12_ sky130_fd_sc_hd__buf_4
Xmux_top_ipin_12.mux_l2_in_1_ chanx_left_in[13] mux_top_ipin_12.mux_l1_in_2_/X mux_top_ipin_12.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_12.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_12.mux_l2_in_0_ mux_top_ipin_12.mux_l1_in_1_/X mux_top_ipin_12.mux_l1_in_0_/X
+ mux_top_ipin_12.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_12.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_5.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_12.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_12.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/A
+ VGND VGND VPWR VPWR mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_14_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_12.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_12.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_8.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_8_ sky130_fd_sc_hd__buf_4
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE ccff_tail
+ IO_ISOL_N VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR sky130_fd_sc_hd__or2b_4
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ mux_top_ipin_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_15.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_15.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_1.mux_l2_in_3_ _23_/HI chanx_right_in[14] mux_top_ipin_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_12.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_12.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_top_ipin_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_1.mux_l4_in_0_ mux_top_ipin_1.mux_l3_in_1_/X mux_top_ipin_1.mux_l3_in_0_/X
+ mux_top_ipin_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_15.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_15_ sky130_fd_sc_hd__buf_4
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_69_ chanx_left_in[7] VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_6.mux_l2_in_3_ _17_/HI chanx_right_in[19] mux_top_ipin_6.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_1.mux_l3_in_1_ mux_top_ipin_1.mux_l2_in_3_/X mux_top_ipin_1.mux_l2_in_2_/X
+ mux_top_ipin_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_15.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_15.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_1.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_top_ipin_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_6.mux_l4_in_0_ mux_top_ipin_6.mux_l3_in_1_/X mux_top_ipin_6.mux_l3_in_0_/X
+ mux_top_ipin_6.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_12.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_ipin_12.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_6.mux_l3_in_1_ mux_top_ipin_6.mux_l2_in_3_/X mux_top_ipin_6.mux_l2_in_2_/X
+ mux_top_ipin_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_1_ sky130_fd_sc_hd__buf_4
X_68_ chanx_left_in[8] VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_top_ipin_5.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_6.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[11] mux_top_ipin_6.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.mux_l3_in_0_ mux_top_ipin_1.mux_l2_in_1_/X mux_top_ipin_1.mux_l2_in_0_/X
+ mux_top_ipin_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_15.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_15.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_13.mux_l2_in_3_ _27_/HI chanx_right_in[18] mux_top_ipin_13.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_top_ipin_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_11.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_12.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_13.mux_l4_in_0_ mux_top_ipin_13.mux_l3_in_1_/X mux_top_ipin_13.mux_l3_in_0_/X
+ mux_top_ipin_13.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_13.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_ mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_/CLK
+ mux_top_ipin_8.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_6.mux_l3_in_0_ mux_top_ipin_6.mux_l2_in_1_/X mux_top_ipin_6.mux_l2_in_0_/X
+ mux_top_ipin_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_13.mux_l3_in_1_ mux_top_ipin_13.mux_l2_in_3_/X mux_top_ipin_13.mux_l2_in_2_/X
+ mux_top_ipin_13.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_13.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_67_ chanx_left_in[9] VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_top_ipin_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_6.mux_l2_in_1_ chanx_left_in[11] chanx_right_in[3] mux_top_ipin_6.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_ mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_/CLK
+ mux_top_ipin_14.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_15.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_13.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_top_ipin_13.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_1.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_1.mux_l1_in_0_/X mux_top_ipin_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

