VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_3__0_
  CLASS BLOCK ;
  FOREIGN sb_3__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 6.160 140.000 6.760 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 137.600 4.050 140.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 2.400 ;
    END
  END address[5]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 2.400 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 137.600 11.870 140.000 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 2.400 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 18.400 140.000 19.000 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 2.400 30.560 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.400 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.400 39.400 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.400 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 2.400 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 2.400 48.240 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 137.600 20.150 140.000 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.400 57.080 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.400 65.920 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 2.400 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 2.400 74.760 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 2.400 82.920 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 2.400 ;
    END
  END chanx_left_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 2.400 91.760 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 137.600 28.430 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 137.600 36.710 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 2.400 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 2.400 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 31.320 140.000 31.920 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 2.400 109.440 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.710 137.600 44.990 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.990 137.600 53.270 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 2.400 118.280 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.240 140.000 44.840 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 56.480 140.000 57.080 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.400 127.120 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.270 137.600 61.550 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 2.400 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 2.400 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 137.600 85.930 140.000 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.930 137.600 94.210 140.000 ;
    END
  END left_bottom_grid_pin_13_
  PIN left_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.210 137.600 102.490 140.000 ;
    END
  END left_bottom_grid_pin_15_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 2.400 135.960 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 82.320 140.000 82.920 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 137.600 77.650 140.000 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 95.240 140.000 95.840 ;
    END
  END left_bottom_grid_pin_9_
  PIN left_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 2.400 ;
    END
  END left_top_grid_pin_10_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 107.480 140.000 108.080 ;
    END
  END top_left_grid_pin_13_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 2.400 ;
    END
  END top_right_grid_pin_11_
  PIN top_right_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 133.320 140.000 133.920 ;
    END
  END top_right_grid_pin_13_
  PIN top_right_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.330 137.600 135.610 140.000 ;
    END
  END top_right_grid_pin_15_
  PIN top_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 137.600 110.770 140.000 ;
    END
  END top_right_grid_pin_1_
  PIN top_right_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 120.400 140.000 121.000 ;
    END
  END top_right_grid_pin_3_
  PIN top_right_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.770 137.600 119.050 140.000 ;
    END
  END top_right_grid_pin_5_
  PIN top_right_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 137.600 127.330 140.000 ;
    END
  END top_right_grid_pin_7_
  PIN top_right_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 2.400 ;
    END
  END top_right_grid_pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.070 10.640 138.390 135.620 ;
      LAYER met2 ;
        RECT 0.100 137.320 3.490 137.770 ;
        RECT 4.330 137.320 11.310 137.770 ;
        RECT 12.150 137.320 19.590 137.770 ;
        RECT 20.430 137.320 27.870 137.770 ;
        RECT 28.710 137.320 36.150 137.770 ;
        RECT 36.990 137.320 44.430 137.770 ;
        RECT 45.270 137.320 52.710 137.770 ;
        RECT 53.550 137.320 60.990 137.770 ;
        RECT 61.830 137.320 69.270 137.770 ;
        RECT 70.110 137.320 77.090 137.770 ;
        RECT 77.930 137.320 85.370 137.770 ;
        RECT 86.210 137.320 93.650 137.770 ;
        RECT 94.490 137.320 101.930 137.770 ;
        RECT 102.770 137.320 110.210 137.770 ;
        RECT 111.050 137.320 118.490 137.770 ;
        RECT 119.330 137.320 126.770 137.770 ;
        RECT 127.610 137.320 135.050 137.770 ;
        RECT 135.890 137.320 138.370 137.770 ;
        RECT 0.100 2.680 138.370 137.320 ;
        RECT 0.100 0.155 3.490 2.680 ;
        RECT 4.330 0.155 10.850 2.680 ;
        RECT 11.690 0.155 18.670 2.680 ;
        RECT 19.510 0.155 26.490 2.680 ;
        RECT 27.330 0.155 34.310 2.680 ;
        RECT 35.150 0.155 42.130 2.680 ;
        RECT 42.970 0.155 49.950 2.680 ;
        RECT 50.790 0.155 57.770 2.680 ;
        RECT 58.610 0.155 65.590 2.680 ;
        RECT 66.430 0.155 73.410 2.680 ;
        RECT 74.250 0.155 80.770 2.680 ;
        RECT 81.610 0.155 88.590 2.680 ;
        RECT 89.430 0.155 96.410 2.680 ;
        RECT 97.250 0.155 104.230 2.680 ;
        RECT 105.070 0.155 112.050 2.680 ;
        RECT 112.890 0.155 119.870 2.680 ;
        RECT 120.710 0.155 127.690 2.680 ;
        RECT 128.530 0.155 135.510 2.680 ;
        RECT 136.350 0.155 138.370 2.680 ;
      LAYER met3 ;
        RECT 2.800 134.960 138.610 135.360 ;
        RECT 0.310 134.320 138.610 134.960 ;
        RECT 0.310 132.920 137.200 134.320 ;
        RECT 0.310 127.520 138.610 132.920 ;
        RECT 2.800 126.120 138.610 127.520 ;
        RECT 0.310 121.400 138.610 126.120 ;
        RECT 0.310 120.000 137.200 121.400 ;
        RECT 0.310 118.680 138.610 120.000 ;
        RECT 2.800 117.280 138.610 118.680 ;
        RECT 0.310 109.840 138.610 117.280 ;
        RECT 2.800 108.480 138.610 109.840 ;
        RECT 2.800 108.440 137.200 108.480 ;
        RECT 0.310 107.080 137.200 108.440 ;
        RECT 0.310 101.000 138.610 107.080 ;
        RECT 2.800 99.600 138.610 101.000 ;
        RECT 0.310 96.240 138.610 99.600 ;
        RECT 0.310 94.840 137.200 96.240 ;
        RECT 0.310 92.160 138.610 94.840 ;
        RECT 2.800 90.760 138.610 92.160 ;
        RECT 0.310 83.320 138.610 90.760 ;
        RECT 2.800 81.920 137.200 83.320 ;
        RECT 0.310 75.160 138.610 81.920 ;
        RECT 2.800 73.760 138.610 75.160 ;
        RECT 0.310 70.400 138.610 73.760 ;
        RECT 0.310 69.000 137.200 70.400 ;
        RECT 0.310 66.320 138.610 69.000 ;
        RECT 2.800 64.920 138.610 66.320 ;
        RECT 0.310 57.480 138.610 64.920 ;
        RECT 2.800 56.080 137.200 57.480 ;
        RECT 0.310 48.640 138.610 56.080 ;
        RECT 2.800 47.240 138.610 48.640 ;
        RECT 0.310 45.240 138.610 47.240 ;
        RECT 0.310 43.840 137.200 45.240 ;
        RECT 0.310 39.800 138.610 43.840 ;
        RECT 2.800 38.400 138.610 39.800 ;
        RECT 0.310 32.320 138.610 38.400 ;
        RECT 0.310 30.960 137.200 32.320 ;
        RECT 2.800 30.920 137.200 30.960 ;
        RECT 2.800 29.560 138.610 30.920 ;
        RECT 0.310 22.120 138.610 29.560 ;
        RECT 2.800 20.720 138.610 22.120 ;
        RECT 0.310 19.400 138.610 20.720 ;
        RECT 0.310 18.000 137.200 19.400 ;
        RECT 0.310 13.280 138.610 18.000 ;
        RECT 2.800 11.880 138.610 13.280 ;
        RECT 0.310 7.160 138.610 11.880 ;
        RECT 0.310 5.760 137.200 7.160 ;
        RECT 0.310 5.120 138.610 5.760 ;
        RECT 2.800 3.720 138.610 5.120 ;
        RECT 0.310 0.175 138.610 3.720 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END sb_3__0_
END LIBRARY

