magic
tech EFS8A
magscale 1 2
timestamp 1602269098
<< locali >>
rect 23247 24225 23374 24259
rect 24627 20961 24662 20995
rect 11931 19873 12058 19907
rect 8527 18785 8654 18819
rect 7711 18377 7757 18411
rect 19579 18105 19717 18139
rect 10051 16745 10057 16779
rect 19343 16745 19349 16779
rect 10051 16677 10085 16745
rect 19343 16677 19377 16745
rect 9683 14807 9717 14875
rect 9683 14773 9689 14807
rect 13455 14569 13461 14603
rect 15663 14569 15669 14603
rect 19435 14569 19441 14603
rect 13455 14501 13489 14569
rect 15663 14501 15697 14569
rect 19435 14501 19469 14569
rect 24075 14433 24110 14467
rect 18199 14025 18245 14059
rect 14013 13787 14047 14025
rect 18003 13821 18130 13855
rect 20177 12699 20211 12869
rect 20177 12665 20269 12699
rect 10879 12393 10885 12427
rect 10879 12325 10913 12393
rect 14375 11543 14409 11611
rect 14375 11509 14381 11543
rect 19435 11305 19441 11339
rect 19435 11237 19469 11305
rect 1443 10081 1478 10115
rect 9321 9911 9355 10217
rect 18699 9367 18733 9435
rect 18699 9333 18705 9367
rect 17083 8993 17118 9027
rect 14139 7905 14174 7939
rect 22511 7905 22546 7939
rect 18003 7293 18095 7327
rect 22615 6749 22661 6783
rect 6009 6307 6043 6341
rect 5917 6273 6043 6307
rect 24075 4641 24110 4675
rect 6837 4063 6871 4097
rect 6837 4029 6998 4063
rect 22017 3927 22051 4029
rect 17963 3689 17969 3723
rect 13771 3621 13816 3655
rect 17963 3621 17997 3689
rect 22511 3553 22546 3587
rect 23615 2941 23742 2975
rect 7389 2363 7423 2465
<< viali >>
rect 17785 24361 17819 24395
rect 17601 24225 17635 24259
rect 23213 24225 23247 24259
rect 23443 24021 23477 24055
rect 7021 23817 7055 23851
rect 12633 23817 12667 23851
rect 14289 23817 14323 23851
rect 16129 23817 16163 23851
rect 17601 23817 17635 23851
rect 18613 23817 18647 23851
rect 23305 23817 23339 23851
rect 25145 23817 25179 23851
rect 22477 23749 22511 23783
rect 1547 23681 1581 23715
rect 1444 23613 1478 23647
rect 1869 23613 1903 23647
rect 4328 23613 4362 23647
rect 4721 23613 4755 23647
rect 6837 23613 6871 23647
rect 12449 23613 12483 23647
rect 13001 23613 13035 23647
rect 14105 23613 14139 23647
rect 15945 23613 15979 23647
rect 16497 23613 16531 23647
rect 18429 23613 18463 23647
rect 18981 23613 19015 23647
rect 22620 23613 22654 23647
rect 24644 23613 24678 23647
rect 22707 23545 22741 23579
rect 24731 23545 24765 23579
rect 4399 23477 4433 23511
rect 7481 23477 7515 23511
rect 14749 23477 14783 23511
rect 1593 23273 1627 23307
rect 1409 23137 1443 23171
rect 25145 22729 25179 22763
rect 1685 22525 1719 22559
rect 24660 22525 24694 22559
rect 24731 22389 24765 22423
rect 24593 20961 24627 20995
rect 24731 20757 24765 20791
rect 24685 20553 24719 20587
rect 11897 19873 11931 19907
rect 12127 19669 12161 19703
rect 13921 19669 13955 19703
rect 15531 19465 15565 19499
rect 11345 19329 11379 19363
rect 10952 19261 10986 19295
rect 12576 19261 12610 19295
rect 13001 19261 13035 19295
rect 14105 19261 14139 19295
rect 14289 19261 14323 19295
rect 15460 19261 15494 19295
rect 15853 19261 15887 19295
rect 12679 19193 12713 19227
rect 14565 19193 14599 19227
rect 11023 19125 11057 19159
rect 12081 19125 12115 19159
rect 13645 19125 13679 19159
rect 10885 18921 10919 18955
rect 9873 18853 9907 18887
rect 13829 18853 13863 18887
rect 15577 18853 15611 18887
rect 8493 18785 8527 18819
rect 12392 18785 12426 18819
rect 21532 18785 21566 18819
rect 8723 18717 8757 18751
rect 9781 18717 9815 18751
rect 11253 18717 11287 18751
rect 13737 18717 13771 18751
rect 14381 18717 14415 18751
rect 15485 18717 15519 18751
rect 16129 18717 16163 18751
rect 10333 18649 10367 18683
rect 12495 18649 12529 18683
rect 13461 18649 13495 18683
rect 12817 18581 12851 18615
rect 21603 18581 21637 18615
rect 7757 18377 7791 18411
rect 8585 18377 8619 18411
rect 10241 18377 10275 18411
rect 12173 18377 12207 18411
rect 21557 18377 21591 18411
rect 22477 18377 22511 18411
rect 15393 18309 15427 18343
rect 17233 18309 17267 18343
rect 8953 18241 8987 18275
rect 10885 18241 10919 18275
rect 14565 18241 14599 18275
rect 15853 18241 15887 18275
rect 16129 18241 16163 18275
rect 7481 18173 7515 18207
rect 7608 18173 7642 18207
rect 12817 18173 12851 18207
rect 13093 18173 13127 18207
rect 19508 18173 19542 18207
rect 19901 18173 19935 18207
rect 22084 18173 22118 18207
rect 9045 18105 9079 18139
rect 9597 18105 9631 18139
rect 10701 18105 10735 18139
rect 10977 18105 11011 18139
rect 11529 18105 11563 18139
rect 13369 18105 13403 18139
rect 14289 18105 14323 18139
rect 14381 18105 14415 18139
rect 15945 18105 15979 18139
rect 19717 18105 19751 18139
rect 20545 18105 20579 18139
rect 20637 18105 20671 18139
rect 21189 18105 21223 18139
rect 8217 18037 8251 18071
rect 9873 18037 9907 18071
rect 13737 18037 13771 18071
rect 14105 18037 14139 18071
rect 16773 18037 16807 18071
rect 20269 18037 20303 18071
rect 22155 18037 22189 18071
rect 9045 17833 9079 17867
rect 14289 17833 14323 17867
rect 20545 17833 20579 17867
rect 24777 17833 24811 17867
rect 8217 17765 8251 17799
rect 10333 17765 10367 17799
rect 11805 17765 11839 17799
rect 11897 17765 11931 17799
rect 13461 17765 13495 17799
rect 15485 17765 15519 17799
rect 19441 17765 19475 17799
rect 21097 17765 21131 17799
rect 21189 17765 21223 17799
rect 22661 17765 22695 17799
rect 22753 17765 22787 17799
rect 17693 17697 17727 17731
rect 18153 17697 18187 17731
rect 24593 17697 24627 17731
rect 8125 17629 8159 17663
rect 10057 17629 10091 17663
rect 10241 17629 10275 17663
rect 12081 17629 12115 17663
rect 13185 17629 13219 17663
rect 13369 17629 13403 17663
rect 13645 17629 13679 17663
rect 15393 17629 15427 17663
rect 15853 17629 15887 17663
rect 18429 17629 18463 17663
rect 19165 17629 19199 17663
rect 19349 17629 19383 17663
rect 19993 17629 20027 17663
rect 21465 17629 21499 17663
rect 22937 17629 22971 17663
rect 8677 17561 8711 17595
rect 10793 17561 10827 17595
rect 16405 17561 16439 17595
rect 12817 17493 12851 17527
rect 14749 17493 14783 17527
rect 7481 17289 7515 17323
rect 7711 17289 7745 17323
rect 9597 17289 9631 17323
rect 11805 17289 11839 17323
rect 15393 17289 15427 17323
rect 18199 17289 18233 17323
rect 24133 17289 24167 17323
rect 15025 17221 15059 17255
rect 16865 17221 16899 17255
rect 22201 17221 22235 17255
rect 23121 17221 23155 17255
rect 10057 17153 10091 17187
rect 10609 17153 10643 17187
rect 14105 17153 14139 17187
rect 16221 17153 16255 17187
rect 17693 17153 17727 17187
rect 20637 17153 20671 17187
rect 20821 17153 20855 17187
rect 23673 17153 23707 17187
rect 7640 17085 7674 17119
rect 8033 17085 8067 17119
rect 8677 17085 8711 17119
rect 12633 17085 12667 17119
rect 12909 17085 12943 17119
rect 18128 17085 18162 17119
rect 22360 17085 22394 17119
rect 22753 17085 22787 17119
rect 8585 17017 8619 17051
rect 8998 17017 9032 17051
rect 10425 17017 10459 17051
rect 10930 17017 10964 17051
rect 12265 17017 12299 17051
rect 13185 17017 13219 17051
rect 14426 17017 14460 17051
rect 15761 17017 15795 17051
rect 15945 17017 15979 17051
rect 16037 17017 16071 17051
rect 19257 17017 19291 17051
rect 19349 17017 19383 17051
rect 19901 17017 19935 17051
rect 20913 17017 20947 17051
rect 21465 17017 21499 17051
rect 11529 16949 11563 16983
rect 13461 16949 13495 16983
rect 13921 16949 13955 16983
rect 17417 16949 17451 16983
rect 18613 16949 18647 16983
rect 18981 16949 19015 16983
rect 20177 16949 20211 16983
rect 21741 16949 21775 16983
rect 22431 16949 22465 16983
rect 24593 16949 24627 16983
rect 7941 16745 7975 16779
rect 10057 16745 10091 16779
rect 10609 16745 10643 16779
rect 10885 16745 10919 16779
rect 15025 16745 15059 16779
rect 16221 16745 16255 16779
rect 19349 16745 19383 16779
rect 19901 16745 19935 16779
rect 20729 16745 20763 16779
rect 7205 16677 7239 16711
rect 8769 16677 8803 16711
rect 9045 16677 9079 16711
rect 11621 16677 11655 16711
rect 11713 16677 11747 16711
rect 13277 16677 13311 16711
rect 13737 16677 13771 16711
rect 13829 16677 13863 16711
rect 14381 16677 14415 16711
rect 15622 16677 15656 16711
rect 21097 16677 21131 16711
rect 21649 16677 21683 16711
rect 22569 16677 22603 16711
rect 22661 16677 22695 16711
rect 6745 16609 6779 16643
rect 7021 16609 7055 16643
rect 8125 16609 8159 16643
rect 8493 16609 8527 16643
rect 17049 16609 17083 16643
rect 17509 16609 17543 16643
rect 18981 16609 19015 16643
rect 9689 16541 9723 16575
rect 11897 16541 11931 16575
rect 15301 16541 15335 16575
rect 17785 16541 17819 16575
rect 18061 16541 18095 16575
rect 21005 16541 21039 16575
rect 22845 16541 22879 16575
rect 12633 16405 12667 16439
rect 18797 16405 18831 16439
rect 8125 16201 8159 16235
rect 9413 16201 9447 16235
rect 9781 16201 9815 16235
rect 11897 16201 11931 16235
rect 14289 16201 14323 16235
rect 14933 16201 14967 16235
rect 18981 16201 19015 16235
rect 19947 16201 19981 16235
rect 20729 16201 20763 16235
rect 22201 16201 22235 16235
rect 22523 16201 22557 16235
rect 22937 16201 22971 16235
rect 23213 16201 23247 16235
rect 10517 16133 10551 16167
rect 12909 16133 12943 16167
rect 19625 16133 19659 16167
rect 6561 16065 6595 16099
rect 7757 16065 7791 16099
rect 9045 16065 9079 16099
rect 11621 16065 11655 16099
rect 13093 16065 13127 16099
rect 15577 16065 15611 16099
rect 15853 16065 15887 16099
rect 18061 16065 18095 16099
rect 20913 16065 20947 16099
rect 8309 15997 8343 16031
rect 8769 15997 8803 16031
rect 19844 15997 19878 16031
rect 20269 15997 20303 16031
rect 22452 15997 22486 16031
rect 7113 15929 7147 15963
rect 9965 15929 9999 15963
rect 10057 15929 10091 15963
rect 13414 15929 13448 15963
rect 15301 15929 15335 15963
rect 15669 15929 15703 15963
rect 17049 15929 17083 15963
rect 18382 15929 18416 15963
rect 21005 15929 21039 15963
rect 21557 15929 21591 15963
rect 10885 15861 10919 15895
rect 14013 15861 14047 15895
rect 16497 15861 16531 15895
rect 17417 15861 17451 15895
rect 17785 15861 17819 15895
rect 19349 15861 19383 15895
rect 21833 15861 21867 15895
rect 1593 15657 1627 15691
rect 13185 15657 13219 15691
rect 13553 15657 13587 15691
rect 16865 15657 16899 15691
rect 20729 15657 20763 15691
rect 22569 15657 22603 15691
rect 9873 15589 9907 15623
rect 11529 15589 11563 15623
rect 13829 15589 13863 15623
rect 15485 15589 15519 15623
rect 16313 15589 16347 15623
rect 18290 15589 18324 15623
rect 21097 15589 21131 15623
rect 1409 15521 1443 15555
rect 10425 15521 10459 15555
rect 12081 15521 12115 15555
rect 19784 15521 19818 15555
rect 9781 15453 9815 15487
rect 11437 15453 11471 15487
rect 13737 15453 13771 15487
rect 14381 15453 14415 15487
rect 15393 15453 15427 15487
rect 15853 15453 15887 15487
rect 17969 15453 18003 15487
rect 21005 15453 21039 15487
rect 21649 15453 21683 15487
rect 8769 15385 8803 15419
rect 18889 15385 18923 15419
rect 8401 15317 8435 15351
rect 9321 15317 9355 15351
rect 10793 15317 10827 15351
rect 19165 15317 19199 15351
rect 19855 15317 19889 15351
rect 9229 15113 9263 15147
rect 10241 15113 10275 15147
rect 10517 15113 10551 15147
rect 11161 15113 11195 15147
rect 13645 15113 13679 15147
rect 13921 15113 13955 15147
rect 15209 15113 15243 15147
rect 17049 15113 17083 15147
rect 17509 15113 17543 15147
rect 18199 15113 18233 15147
rect 19993 15113 20027 15147
rect 22385 15113 22419 15147
rect 8447 15045 8481 15079
rect 14749 15045 14783 15079
rect 12173 14977 12207 15011
rect 16221 14977 16255 15011
rect 19073 14977 19107 15011
rect 21097 14977 21131 15011
rect 22753 14977 22787 15011
rect 8376 14909 8410 14943
rect 9321 14909 9355 14943
rect 11396 14909 11430 14943
rect 11805 14909 11839 14943
rect 12449 14909 12483 14943
rect 12909 14909 12943 14943
rect 18096 14909 18130 14943
rect 18521 14909 18555 14943
rect 11483 14841 11517 14875
rect 13185 14841 13219 14875
rect 14197 14841 14231 14875
rect 14289 14841 14323 14875
rect 15485 14841 15519 14875
rect 15761 14841 15795 14875
rect 15853 14841 15887 14875
rect 19435 14841 19469 14875
rect 21166 14841 21200 14875
rect 21741 14841 21775 14875
rect 1685 14773 1719 14807
rect 8769 14773 8803 14807
rect 9689 14773 9723 14807
rect 16773 14773 16807 14807
rect 17785 14773 17819 14807
rect 18981 14773 19015 14807
rect 20269 14773 20303 14807
rect 20821 14773 20855 14807
rect 22017 14773 22051 14807
rect 9873 14569 9907 14603
rect 11437 14569 11471 14603
rect 11713 14569 11747 14603
rect 13001 14569 13035 14603
rect 13461 14569 13495 14603
rect 14013 14569 14047 14603
rect 15669 14569 15703 14603
rect 16221 14569 16255 14603
rect 19441 14569 19475 14603
rect 19993 14569 20027 14603
rect 20637 14569 20671 14603
rect 22569 14569 22603 14603
rect 10838 14501 10872 14535
rect 17785 14501 17819 14535
rect 21005 14501 21039 14535
rect 21097 14501 21131 14535
rect 8217 14433 8251 14467
rect 8585 14433 8619 14467
rect 17325 14433 17359 14467
rect 17509 14433 17543 14467
rect 22477 14433 22511 14467
rect 22937 14433 22971 14467
rect 24041 14433 24075 14467
rect 8769 14365 8803 14399
rect 10517 14365 10551 14399
rect 13093 14365 13127 14399
rect 15301 14365 15335 14399
rect 19073 14365 19107 14399
rect 21281 14365 21315 14399
rect 9229 14229 9263 14263
rect 12449 14229 12483 14263
rect 14289 14229 14323 14263
rect 18061 14229 18095 14263
rect 18889 14229 18923 14263
rect 24179 14229 24213 14263
rect 1593 14025 1627 14059
rect 9137 14025 9171 14059
rect 10149 14025 10183 14059
rect 11437 14025 11471 14059
rect 12173 14025 12207 14059
rect 13461 14025 13495 14059
rect 14013 14025 14047 14059
rect 14105 14025 14139 14059
rect 15209 14025 15243 14059
rect 17785 14025 17819 14059
rect 18245 14025 18279 14059
rect 20177 14025 20211 14059
rect 22385 14025 22419 14059
rect 23029 14025 23063 14059
rect 24225 14025 24259 14059
rect 10517 13957 10551 13991
rect 9229 13889 9263 13923
rect 1409 13821 1443 13855
rect 1961 13821 1995 13855
rect 7941 13821 7975 13855
rect 8125 13821 8159 13855
rect 11044 13821 11078 13855
rect 12449 13821 12483 13855
rect 13001 13821 13035 13855
rect 16221 13957 16255 13991
rect 20453 13957 20487 13991
rect 17141 13889 17175 13923
rect 14289 13821 14323 13855
rect 15945 13821 15979 13855
rect 16405 13821 16439 13855
rect 16865 13821 16899 13855
rect 17417 13821 17451 13855
rect 17969 13821 18003 13855
rect 19253 13821 19287 13855
rect 20821 13821 20855 13855
rect 21005 13821 21039 13855
rect 21465 13821 21499 13855
rect 22636 13821 22670 13855
rect 23740 13821 23774 13855
rect 7573 13753 7607 13787
rect 8401 13753 8435 13787
rect 9550 13753 9584 13787
rect 13185 13753 13219 13787
rect 14013 13753 14047 13787
rect 14651 13753 14685 13787
rect 15577 13753 15611 13787
rect 19578 13753 19612 13787
rect 22017 13753 22051 13787
rect 24501 13753 24535 13787
rect 7205 13685 7239 13719
rect 8769 13685 8803 13719
rect 11115 13685 11149 13719
rect 18797 13685 18831 13719
rect 19073 13685 19107 13719
rect 21097 13685 21131 13719
rect 22707 13685 22741 13719
rect 23811 13685 23845 13719
rect 10701 13481 10735 13515
rect 11069 13481 11103 13515
rect 13093 13481 13127 13515
rect 20177 13481 20211 13515
rect 20729 13481 20763 13515
rect 23765 13481 23799 13515
rect 7757 13413 7791 13447
rect 11345 13413 11379 13447
rect 11437 13413 11471 13447
rect 12541 13413 12575 13447
rect 18061 13413 18095 13447
rect 19251 13413 19285 13447
rect 21097 13413 21131 13447
rect 22661 13413 22695 13447
rect 22845 13413 22879 13447
rect 22937 13413 22971 13447
rect 8033 13345 8067 13379
rect 8493 13345 8527 13379
rect 9965 13345 9999 13379
rect 10149 13345 10183 13379
rect 13185 13345 13219 13379
rect 13645 13345 13679 13379
rect 16037 13345 16071 13379
rect 16313 13345 16347 13379
rect 17325 13345 17359 13379
rect 17785 13345 17819 13379
rect 24660 13345 24694 13379
rect 8769 13277 8803 13311
rect 10241 13277 10275 13311
rect 11621 13277 11655 13311
rect 13737 13277 13771 13311
rect 15485 13277 15519 13311
rect 16497 13277 16531 13311
rect 18889 13277 18923 13311
rect 21005 13277 21039 13311
rect 21649 13277 21683 13311
rect 23489 13277 23523 13311
rect 14289 13209 14323 13243
rect 24731 13209 24765 13243
rect 9229 13141 9263 13175
rect 18429 13141 18463 13175
rect 19809 13141 19843 13175
rect 1593 12937 1627 12971
rect 8125 12937 8159 12971
rect 11805 12937 11839 12971
rect 12817 12937 12851 12971
rect 13185 12937 13219 12971
rect 15945 12937 15979 12971
rect 17417 12937 17451 12971
rect 18981 12937 19015 12971
rect 22385 12937 22419 12971
rect 24777 12937 24811 12971
rect 25421 12937 25455 12971
rect 8493 12869 8527 12903
rect 12173 12869 12207 12903
rect 15485 12869 15519 12903
rect 19349 12869 19383 12903
rect 20177 12869 20211 12903
rect 10885 12801 10919 12835
rect 13645 12801 13679 12835
rect 14933 12801 14967 12835
rect 19717 12801 19751 12835
rect 1409 12733 1443 12767
rect 9505 12733 9539 12767
rect 9689 12733 9723 12767
rect 16313 12733 16347 12767
rect 16589 12733 16623 12767
rect 16865 12733 16899 12767
rect 18061 12733 18095 12767
rect 19844 12733 19878 12767
rect 21097 12801 21131 12835
rect 23029 12801 23063 12835
rect 23765 12801 23799 12835
rect 24041 12801 24075 12835
rect 20821 12733 20855 12767
rect 22604 12733 22638 12767
rect 25237 12733 25271 12767
rect 25789 12733 25823 12767
rect 9137 12665 9171 12699
rect 10241 12665 10275 12699
rect 10701 12665 10735 12699
rect 10977 12665 11011 12699
rect 11529 12665 11563 12699
rect 13369 12665 13403 12699
rect 13461 12665 13495 12699
rect 15025 12665 15059 12699
rect 17141 12665 17175 12699
rect 18382 12665 18416 12699
rect 20269 12665 20303 12699
rect 21189 12665 21223 12699
rect 21741 12665 21775 12699
rect 23397 12665 23431 12699
rect 23857 12665 23891 12699
rect 2053 12597 2087 12631
rect 9321 12597 9355 12631
rect 14749 12597 14783 12631
rect 17877 12597 17911 12631
rect 19947 12597 19981 12631
rect 22017 12597 22051 12631
rect 22707 12597 22741 12631
rect 10885 12393 10919 12427
rect 11437 12393 11471 12427
rect 14013 12393 14047 12427
rect 14335 12393 14369 12427
rect 14933 12393 14967 12427
rect 16773 12393 16807 12427
rect 17325 12393 17359 12427
rect 18613 12393 18647 12427
rect 20361 12393 20395 12427
rect 9965 12325 9999 12359
rect 12449 12325 12483 12359
rect 15485 12325 15519 12359
rect 16037 12325 16071 12359
rect 16405 12325 16439 12359
rect 18014 12325 18048 12359
rect 21005 12325 21039 12359
rect 21097 12325 21131 12359
rect 22661 12325 22695 12359
rect 24225 12325 24259 12359
rect 8620 12257 8654 12291
rect 8723 12257 8757 12291
rect 13737 12257 13771 12291
rect 14243 12257 14277 12291
rect 19876 12257 19910 12291
rect 10517 12189 10551 12223
rect 12357 12189 12391 12223
rect 12633 12189 12667 12223
rect 15393 12189 15427 12223
rect 17693 12189 17727 12223
rect 21649 12189 21683 12223
rect 22569 12189 22603 12223
rect 22845 12189 22879 12223
rect 24133 12189 24167 12223
rect 24409 12189 24443 12223
rect 9413 12121 9447 12155
rect 19947 12121 19981 12155
rect 9137 12053 9171 12087
rect 10333 12053 10367 12087
rect 13369 12053 13403 12087
rect 19625 12053 19659 12087
rect 20637 12053 20671 12087
rect 23673 12053 23707 12087
rect 10149 11849 10183 11883
rect 10517 11849 10551 11883
rect 11529 11849 11563 11883
rect 11897 11849 11931 11883
rect 13553 11849 13587 11883
rect 14933 11849 14967 11883
rect 18659 11849 18693 11883
rect 20913 11849 20947 11883
rect 21281 11849 21315 11883
rect 23029 11849 23063 11883
rect 24777 11849 24811 11883
rect 16405 11781 16439 11815
rect 19349 11781 19383 11815
rect 24317 11781 24351 11815
rect 8493 11713 8527 11747
rect 9505 11713 9539 11747
rect 10609 11713 10643 11747
rect 14013 11713 14047 11747
rect 15669 11713 15703 11747
rect 15853 11713 15887 11747
rect 19533 11713 19567 11747
rect 22385 11713 22419 11747
rect 23489 11713 23523 11747
rect 23765 11713 23799 11747
rect 25237 11713 25271 11747
rect 7665 11645 7699 11679
rect 7849 11645 7883 11679
rect 9045 11645 9079 11679
rect 9137 11645 9171 11679
rect 9321 11645 9355 11679
rect 12725 11645 12759 11679
rect 13001 11645 13035 11679
rect 13185 11645 13219 11679
rect 18588 11645 18622 11679
rect 18981 11645 19015 11679
rect 20453 11645 20487 11679
rect 21833 11645 21867 11679
rect 8217 11577 8251 11611
rect 10971 11577 11005 11611
rect 12265 11577 12299 11611
rect 15945 11577 15979 11611
rect 18337 11577 18371 11611
rect 19854 11577 19888 11611
rect 22109 11577 22143 11611
rect 22201 11577 22235 11611
rect 23857 11577 23891 11611
rect 7573 11509 7607 11543
rect 8861 11509 8895 11543
rect 13829 11509 13863 11543
rect 14381 11509 14415 11543
rect 15209 11509 15243 11543
rect 16773 11509 16807 11543
rect 17785 11509 17819 11543
rect 10057 11305 10091 11339
rect 10793 11305 10827 11339
rect 12817 11305 12851 11339
rect 16221 11305 16255 11339
rect 19441 11305 19475 11339
rect 20361 11305 20395 11339
rect 22569 11305 22603 11339
rect 24133 11305 24167 11339
rect 24409 11305 24443 11339
rect 11529 11237 11563 11271
rect 12541 11237 12575 11271
rect 13455 11237 13489 11271
rect 15622 11237 15656 11271
rect 21189 11237 21223 11271
rect 21741 11237 21775 11271
rect 22946 11237 22980 11271
rect 23489 11237 23523 11271
rect 7849 11169 7883 11203
rect 8769 11169 8803 11203
rect 10057 11169 10091 11203
rect 10333 11169 10367 11203
rect 12081 11169 12115 11203
rect 15301 11169 15335 11203
rect 17509 11169 17543 11203
rect 17969 11169 18003 11203
rect 19073 11169 19107 11203
rect 24593 11169 24627 11203
rect 24869 11169 24903 11203
rect 7757 11101 7791 11135
rect 11437 11101 11471 11135
rect 13093 11101 13127 11135
rect 15117 11101 15151 11135
rect 18245 11101 18279 11135
rect 21097 11101 21131 11135
rect 22845 11101 22879 11135
rect 14013 11033 14047 11067
rect 7297 10965 7331 10999
rect 7573 10965 7607 10999
rect 9229 10965 9263 10999
rect 11161 10965 11195 10999
rect 14289 10965 14323 10999
rect 16497 10965 16531 10999
rect 19993 10965 20027 10999
rect 22109 10965 22143 10999
rect 7021 10761 7055 10795
rect 11529 10761 11563 10795
rect 12817 10761 12851 10795
rect 13737 10761 13771 10795
rect 14841 10761 14875 10795
rect 17233 10761 17267 10795
rect 20637 10761 20671 10795
rect 22753 10761 22787 10795
rect 24685 10761 24719 10795
rect 25421 10761 25455 10795
rect 8861 10693 8895 10727
rect 21833 10693 21867 10727
rect 7757 10625 7791 10659
rect 8125 10625 8159 10659
rect 8953 10625 8987 10659
rect 9321 10625 9355 10659
rect 9689 10625 9723 10659
rect 10057 10625 10091 10659
rect 10885 10625 10919 10659
rect 13047 10625 13081 10659
rect 13921 10625 13955 10659
rect 15761 10625 15795 10659
rect 16037 10625 16071 10659
rect 18061 10625 18095 10659
rect 19441 10625 19475 10659
rect 7389 10557 7423 10591
rect 8732 10557 8766 10591
rect 10425 10557 10459 10591
rect 10701 10557 10735 10591
rect 12960 10557 12994 10591
rect 20361 10557 20395 10591
rect 21005 10557 21039 10591
rect 23949 10557 23983 10591
rect 24133 10557 24167 10591
rect 25237 10557 25271 10591
rect 25789 10557 25823 10591
rect 7205 10489 7239 10523
rect 8585 10489 8619 10523
rect 14243 10489 14277 10523
rect 15853 10489 15887 10523
rect 19762 10489 19796 10523
rect 21281 10489 21315 10523
rect 21373 10489 21407 10523
rect 8493 10421 8527 10455
rect 11161 10421 11195 10455
rect 11897 10421 11931 10455
rect 13461 10421 13495 10455
rect 15393 10421 15427 10455
rect 16681 10421 16715 10455
rect 17601 10421 17635 10455
rect 18705 10421 18739 10455
rect 19073 10421 19107 10455
rect 22385 10421 22419 10455
rect 23397 10421 23431 10455
rect 23765 10421 23799 10455
rect 25053 10421 25087 10455
rect 9321 10217 9355 10251
rect 9413 10217 9447 10251
rect 10333 10217 10367 10251
rect 13093 10217 13127 10251
rect 15117 10217 15151 10251
rect 18981 10217 19015 10251
rect 19349 10217 19383 10251
rect 19993 10217 20027 10251
rect 20729 10217 20763 10251
rect 22017 10217 22051 10251
rect 23765 10217 23799 10251
rect 5457 10149 5491 10183
rect 1409 10081 1443 10115
rect 4112 10081 4146 10115
rect 7757 10081 7791 10115
rect 7941 10081 7975 10115
rect 8309 10081 8343 10115
rect 4215 10013 4249 10047
rect 5365 10013 5399 10047
rect 6009 10013 6043 10047
rect 8769 10013 8803 10047
rect 12817 10149 12851 10183
rect 21097 10149 21131 10183
rect 9689 10081 9723 10115
rect 12357 10081 12391 10115
rect 12541 10081 12575 10115
rect 13645 10081 13679 10115
rect 14197 10081 14231 10115
rect 15945 10081 15979 10115
rect 16129 10081 16163 10115
rect 17969 10081 18003 10115
rect 18429 10081 18463 10115
rect 19533 10081 19567 10115
rect 22753 10081 22787 10115
rect 22937 10081 22971 10115
rect 10057 10013 10091 10047
rect 14381 10013 14415 10047
rect 16221 10013 16255 10047
rect 18705 10013 18739 10047
rect 21005 10013 21039 10047
rect 23029 10013 23063 10047
rect 11897 9945 11931 9979
rect 21557 9945 21591 9979
rect 1547 9877 1581 9911
rect 7297 9877 7331 9911
rect 9045 9877 9079 9911
rect 9321 9877 9355 9911
rect 9827 9877 9861 9911
rect 9965 9877 9999 9911
rect 10701 9877 10735 9911
rect 11069 9877 11103 9911
rect 15577 9877 15611 9911
rect 3985 9673 4019 9707
rect 6561 9673 6595 9707
rect 7573 9673 7607 9707
rect 8309 9673 8343 9707
rect 9689 9673 9723 9707
rect 12173 9673 12207 9707
rect 20269 9673 20303 9707
rect 20637 9673 20671 9707
rect 22523 9673 22557 9707
rect 23305 9673 23339 9707
rect 4307 9605 4341 9639
rect 9321 9605 9355 9639
rect 15393 9605 15427 9639
rect 19257 9605 19291 9639
rect 22201 9605 22235 9639
rect 5273 9537 5307 9571
rect 6193 9537 6227 9571
rect 9413 9537 9447 9571
rect 10793 9537 10827 9571
rect 11437 9537 11471 9571
rect 12541 9537 12575 9571
rect 15025 9537 15059 9571
rect 15577 9537 15611 9571
rect 16037 9537 16071 9571
rect 18337 9537 18371 9571
rect 19993 9537 20027 9571
rect 20913 9537 20947 9571
rect 21189 9537 21223 9571
rect 4236 9469 4270 9503
rect 4629 9469 4663 9503
rect 7389 9469 7423 9503
rect 9192 9469 9226 9503
rect 10701 9469 10735 9503
rect 10977 9469 11011 9503
rect 14013 9469 14047 9503
rect 14565 9469 14599 9503
rect 22420 9469 22454 9503
rect 22845 9469 22879 9503
rect 5089 9401 5123 9435
rect 5365 9401 5399 9435
rect 5917 9401 5951 9435
rect 9045 9401 9079 9435
rect 11713 9401 11747 9435
rect 12633 9401 12667 9435
rect 13185 9401 13219 9435
rect 15669 9401 15703 9435
rect 16589 9401 16623 9435
rect 21005 9401 21039 9435
rect 1593 9333 1627 9367
rect 7113 9333 7147 9367
rect 8953 9333 8987 9367
rect 10057 9333 10091 9367
rect 10517 9333 10551 9367
rect 13645 9333 13679 9367
rect 14197 9333 14231 9367
rect 17509 9333 17543 9367
rect 17785 9333 17819 9367
rect 18705 9333 18739 9367
rect 21833 9333 21867 9367
rect 7205 9129 7239 9163
rect 11069 9129 11103 9163
rect 12357 9129 12391 9163
rect 17187 9129 17221 9163
rect 19993 9129 20027 9163
rect 5911 9061 5945 9095
rect 10425 9061 10459 9095
rect 13185 9061 13219 9095
rect 15663 9061 15697 9095
rect 18791 9061 18825 9095
rect 21097 9061 21131 9095
rect 7481 8993 7515 9027
rect 9137 8993 9171 9027
rect 9689 8993 9723 9027
rect 10701 8993 10735 9027
rect 11621 8993 11655 9027
rect 11805 8993 11839 9027
rect 15301 8993 15335 9027
rect 17049 8993 17083 9027
rect 4537 8925 4571 8959
rect 5549 8925 5583 8959
rect 7297 8925 7331 8959
rect 9836 8925 9870 8959
rect 10057 8925 10091 8959
rect 12081 8925 12115 8959
rect 13093 8925 13127 8959
rect 13369 8925 13403 8959
rect 18429 8925 18463 8959
rect 21005 8925 21039 8959
rect 22477 8925 22511 8959
rect 5273 8857 5307 8891
rect 6469 8857 6503 8891
rect 14105 8857 14139 8891
rect 21557 8857 21591 8891
rect 21925 8857 21959 8891
rect 6837 8789 6871 8823
rect 8585 8789 8619 8823
rect 9505 8789 9539 8823
rect 9965 8789 9999 8823
rect 12817 8789 12851 8823
rect 16221 8789 16255 8823
rect 18061 8789 18095 8823
rect 19349 8789 19383 8823
rect 19625 8789 19659 8823
rect 8033 8585 8067 8619
rect 10701 8585 10735 8619
rect 11253 8585 11287 8619
rect 13369 8585 13403 8619
rect 15853 8585 15887 8619
rect 18475 8585 18509 8619
rect 21005 8585 21039 8619
rect 24777 8585 24811 8619
rect 8493 8517 8527 8551
rect 17601 8517 17635 8551
rect 5273 8449 5307 8483
rect 5917 8449 5951 8483
rect 7205 8449 7239 8483
rect 12449 8449 12483 8483
rect 14013 8449 14047 8483
rect 17141 8449 17175 8483
rect 19349 8449 19383 8483
rect 21465 8449 21499 8483
rect 8585 8381 8619 8415
rect 9045 8381 9079 8415
rect 9413 8381 9447 8415
rect 9873 8381 9907 8415
rect 11345 8381 11379 8415
rect 13645 8381 13679 8415
rect 14933 8381 14967 8415
rect 16748 8381 16782 8415
rect 18404 8381 18438 8415
rect 18797 8381 18831 8415
rect 24593 8381 24627 8415
rect 25145 8381 25179 8415
rect 5089 8313 5123 8347
rect 5365 8313 5399 8347
rect 6929 8313 6963 8347
rect 7021 8313 7055 8347
rect 12770 8313 12804 8347
rect 15295 8313 15329 8347
rect 19165 8313 19199 8347
rect 19670 8313 19704 8347
rect 21189 8313 21223 8347
rect 21281 8313 21315 8347
rect 6193 8245 6227 8279
rect 6653 8245 6687 8279
rect 8677 8245 8711 8279
rect 10425 8245 10459 8279
rect 11805 8245 11839 8279
rect 12173 8245 12207 8279
rect 14841 8245 14875 8279
rect 16129 8245 16163 8279
rect 16819 8245 16853 8279
rect 20269 8245 20303 8279
rect 20637 8245 20671 8279
rect 22109 8245 22143 8279
rect 5273 8041 5307 8075
rect 5595 8041 5629 8075
rect 7481 8041 7515 8075
rect 10241 8041 10275 8075
rect 13277 8041 13311 8075
rect 13553 8041 13587 8075
rect 15485 8041 15519 8075
rect 6285 7973 6319 8007
rect 6653 7973 6687 8007
rect 9965 7973 9999 8007
rect 12678 7973 12712 8007
rect 16542 7973 16576 8007
rect 19441 7973 19475 8007
rect 19993 7973 20027 8007
rect 21097 7973 21131 8007
rect 5524 7905 5558 7939
rect 8677 7905 8711 7939
rect 10517 7905 10551 7939
rect 10793 7905 10827 7939
rect 14105 7905 14139 7939
rect 16221 7905 16255 7939
rect 18004 7905 18038 7939
rect 22477 7905 22511 7939
rect 6561 7837 6595 7871
rect 7205 7837 7239 7871
rect 11253 7837 11287 7871
rect 11897 7837 11931 7871
rect 12357 7837 12391 7871
rect 19165 7837 19199 7871
rect 19349 7837 19383 7871
rect 21005 7837 21039 7871
rect 21281 7837 21315 7871
rect 5917 7769 5951 7803
rect 10609 7769 10643 7803
rect 8309 7701 8343 7735
rect 9045 7701 9079 7735
rect 12265 7701 12299 7735
rect 14243 7701 14277 7735
rect 14933 7701 14967 7735
rect 16037 7701 16071 7735
rect 17141 7701 17175 7735
rect 18107 7701 18141 7735
rect 18521 7701 18555 7735
rect 22017 7701 22051 7735
rect 22615 7701 22649 7735
rect 6193 7497 6227 7531
rect 8125 7497 8159 7531
rect 13737 7497 13771 7531
rect 15669 7497 15703 7531
rect 19165 7497 19199 7531
rect 22477 7497 22511 7531
rect 1593 7429 1627 7463
rect 14105 7429 14139 7463
rect 16773 7429 16807 7463
rect 20269 7429 20303 7463
rect 5917 7361 5951 7395
rect 6561 7361 6595 7395
rect 6929 7361 6963 7395
rect 7205 7361 7239 7395
rect 14841 7361 14875 7395
rect 16221 7361 16255 7395
rect 18613 7361 18647 7395
rect 19717 7361 19751 7395
rect 21281 7361 21315 7395
rect 21557 7361 21591 7395
rect 1409 7293 1443 7327
rect 1961 7293 1995 7327
rect 5089 7293 5123 7327
rect 5825 7293 5859 7327
rect 9045 7293 9079 7327
rect 11069 7293 11103 7327
rect 11345 7293 11379 7327
rect 12449 7293 12483 7327
rect 12909 7293 12943 7327
rect 14565 7293 14599 7327
rect 14749 7293 14783 7327
rect 17969 7293 18003 7327
rect 18521 7293 18555 7327
rect 7021 7225 7055 7259
rect 8953 7225 8987 7259
rect 10517 7225 10551 7259
rect 11529 7225 11563 7259
rect 16313 7225 16347 7259
rect 19809 7225 19843 7259
rect 21005 7225 21039 7259
rect 21373 7225 21407 7259
rect 8401 7157 8435 7191
rect 8769 7157 8803 7191
rect 10241 7157 10275 7191
rect 11805 7157 11839 7191
rect 12173 7157 12207 7191
rect 12541 7157 12575 7191
rect 15945 7157 15979 7191
rect 17417 7157 17451 7191
rect 17785 7157 17819 7191
rect 19441 7157 19475 7191
rect 6101 6953 6135 6987
rect 7573 6953 7607 6987
rect 8493 6953 8527 6987
rect 10885 6953 10919 6987
rect 16221 6953 16255 6987
rect 21005 6953 21039 6987
rect 21925 6953 21959 6987
rect 24777 6953 24811 6987
rect 6974 6885 7008 6919
rect 12449 6885 12483 6919
rect 16865 6885 16899 6919
rect 19441 6885 19475 6919
rect 19993 6885 20027 6919
rect 5549 6817 5583 6851
rect 11345 6817 11379 6851
rect 11713 6817 11747 6851
rect 12725 6817 12759 6851
rect 13185 6817 13219 6851
rect 15577 6817 15611 6851
rect 17417 6817 17451 6851
rect 18153 6817 18187 6851
rect 18280 6817 18314 6851
rect 20913 6817 20947 6851
rect 21373 6817 21407 6851
rect 22512 6817 22546 6851
rect 23556 6817 23590 6851
rect 24593 6817 24627 6851
rect 6653 6749 6687 6783
rect 11897 6749 11931 6783
rect 13461 6749 13495 6783
rect 16773 6749 16807 6783
rect 19349 6749 19383 6783
rect 22661 6749 22695 6783
rect 10425 6681 10459 6715
rect 14381 6681 14415 6715
rect 18383 6681 18417 6715
rect 19073 6681 19107 6715
rect 20729 6681 20763 6715
rect 23627 6681 23661 6715
rect 5273 6613 5307 6647
rect 5733 6613 5767 6647
rect 6561 6613 6595 6647
rect 8861 6613 8895 6647
rect 15761 6613 15795 6647
rect 18797 6613 18831 6647
rect 20361 6613 20395 6647
rect 16037 6409 16071 6443
rect 16727 6409 16761 6443
rect 17141 6409 17175 6443
rect 17509 6409 17543 6443
rect 19073 6409 19107 6443
rect 19441 6409 19475 6443
rect 20913 6409 20947 6443
rect 22477 6409 22511 6443
rect 25513 6409 25547 6443
rect 6009 6341 6043 6375
rect 6653 6273 6687 6307
rect 10701 6273 10735 6307
rect 13277 6273 13311 6307
rect 15117 6273 15151 6307
rect 15485 6273 15519 6307
rect 19809 6273 19843 6307
rect 21373 6273 21407 6307
rect 22845 6273 22879 6307
rect 24823 6273 24857 6307
rect 5089 6205 5123 6239
rect 5181 6205 5215 6239
rect 5273 6205 5307 6239
rect 5457 6205 5491 6239
rect 6837 6205 6871 6239
rect 6929 6205 6963 6239
rect 7113 6205 7147 6239
rect 8309 6205 8343 6239
rect 8585 6205 8619 6239
rect 9137 6205 9171 6239
rect 9229 6205 9263 6239
rect 9781 6205 9815 6239
rect 10793 6205 10827 6239
rect 11253 6205 11287 6239
rect 11805 6205 11839 6239
rect 12725 6205 12759 6239
rect 16624 6205 16658 6239
rect 17785 6205 17819 6239
rect 18153 6205 18187 6239
rect 23740 6205 23774 6239
rect 24501 6205 24535 6239
rect 24720 6205 24754 6239
rect 7573 6137 7607 6171
rect 11529 6137 11563 6171
rect 13598 6137 13632 6171
rect 15209 6137 15243 6171
rect 18061 6137 18095 6171
rect 19901 6137 19935 6171
rect 20453 6137 20487 6171
rect 21465 6137 21499 6171
rect 22017 6137 22051 6171
rect 25145 6137 25179 6171
rect 6193 6069 6227 6103
rect 7941 6069 7975 6103
rect 8493 6069 8527 6103
rect 10149 6069 10183 6103
rect 12173 6069 12207 6103
rect 13185 6069 13219 6103
rect 14197 6069 14231 6103
rect 14841 6069 14875 6103
rect 16405 6069 16439 6103
rect 23811 6069 23845 6103
rect 24133 6069 24167 6103
rect 5549 5865 5583 5899
rect 6377 5865 6411 5899
rect 8493 5865 8527 5899
rect 13277 5865 13311 5899
rect 15025 5865 15059 5899
rect 22569 5865 22603 5899
rect 24133 5865 24167 5899
rect 7573 5797 7607 5831
rect 10425 5797 10459 5831
rect 12259 5797 12293 5831
rect 13737 5797 13771 5831
rect 13829 5797 13863 5831
rect 15622 5797 15656 5831
rect 17554 5797 17588 5831
rect 19343 5797 19377 5831
rect 21097 5797 21131 5831
rect 21649 5797 21683 5831
rect 6469 5729 6503 5763
rect 6745 5729 6779 5763
rect 7205 5729 7239 5763
rect 8033 5729 8067 5763
rect 8309 5729 8343 5763
rect 9689 5729 9723 5763
rect 9965 5729 9999 5763
rect 10793 5729 10827 5763
rect 11253 5729 11287 5763
rect 11897 5729 11931 5763
rect 15301 5729 15335 5763
rect 18981 5729 19015 5763
rect 22477 5729 22511 5763
rect 22937 5729 22971 5763
rect 24041 5729 24075 5763
rect 24501 5729 24535 5763
rect 8125 5661 8159 5695
rect 9045 5661 9079 5695
rect 14013 5661 14047 5695
rect 17233 5661 17267 5695
rect 21005 5661 21039 5695
rect 5273 5593 5307 5627
rect 6561 5593 6595 5627
rect 9413 5593 9447 5627
rect 9781 5593 9815 5627
rect 18153 5593 18187 5627
rect 20269 5593 20303 5627
rect 7941 5525 7975 5559
rect 11805 5525 11839 5559
rect 12817 5525 12851 5559
rect 14749 5525 14783 5559
rect 16221 5525 16255 5559
rect 18705 5525 18739 5559
rect 19901 5525 19935 5559
rect 20729 5525 20763 5559
rect 21925 5525 21959 5559
rect 6193 5321 6227 5355
rect 7021 5321 7055 5355
rect 7389 5321 7423 5355
rect 9045 5321 9079 5355
rect 14381 5321 14415 5355
rect 20177 5321 20211 5355
rect 23397 5321 23431 5355
rect 24501 5321 24535 5355
rect 9229 5253 9263 5287
rect 15485 5253 15519 5287
rect 15853 5253 15887 5287
rect 10701 5185 10735 5219
rect 13093 5185 13127 5219
rect 16773 5185 16807 5219
rect 18613 5185 18647 5219
rect 20453 5185 20487 5219
rect 20729 5185 20763 5219
rect 22477 5185 22511 5219
rect 7665 5117 7699 5151
rect 8585 5117 8619 5151
rect 9137 5117 9171 5151
rect 9413 5117 9447 5151
rect 10241 5117 10275 5151
rect 10609 5117 10643 5151
rect 11345 5117 11379 5151
rect 14013 5117 14047 5151
rect 14657 5117 14691 5151
rect 19533 5117 19567 5151
rect 21925 5117 21959 5151
rect 22385 5117 22419 5151
rect 23740 5117 23774 5151
rect 24133 5117 24167 5151
rect 24720 5117 24754 5151
rect 25145 5117 25179 5151
rect 7573 5049 7607 5083
rect 9873 5049 9907 5083
rect 13414 5049 13448 5083
rect 14933 5049 14967 5083
rect 15025 5049 15059 5083
rect 16497 5049 16531 5083
rect 16589 5049 16623 5083
rect 17877 5049 17911 5083
rect 18975 5049 19009 5083
rect 20545 5049 20579 5083
rect 24823 5049 24857 5083
rect 6561 4981 6595 5015
rect 11897 4981 11931 5015
rect 12909 4981 12943 5015
rect 16313 4981 16347 5015
rect 17417 4981 17451 5015
rect 18429 4981 18463 5015
rect 19809 4981 19843 5015
rect 21373 4981 21407 5015
rect 21741 4981 21775 5015
rect 22937 4981 22971 5015
rect 23811 4981 23845 5015
rect 7941 4777 7975 4811
rect 8493 4777 8527 4811
rect 11897 4777 11931 4811
rect 13093 4777 13127 4811
rect 15485 4777 15519 4811
rect 16497 4777 16531 4811
rect 19533 4777 19567 4811
rect 20361 4777 20395 4811
rect 20729 4777 20763 4811
rect 21005 4777 21039 4811
rect 21925 4777 21959 4811
rect 22293 4777 22327 4811
rect 22569 4777 22603 4811
rect 7159 4709 7193 4743
rect 12173 4709 12207 4743
rect 13737 4709 13771 4743
rect 14289 4709 14323 4743
rect 17094 4709 17128 4743
rect 18705 4709 18739 4743
rect 7056 4641 7090 4675
rect 8033 4641 8067 4675
rect 8309 4641 8343 4675
rect 9137 4641 9171 4675
rect 9689 4641 9723 4675
rect 10149 4641 10183 4675
rect 10517 4641 10551 4675
rect 11069 4641 11103 4675
rect 14933 4641 14967 4675
rect 15669 4641 15703 4675
rect 16773 4641 16807 4675
rect 20913 4641 20947 4675
rect 21373 4641 21407 4675
rect 22477 4641 22511 4675
rect 22937 4641 22971 4675
rect 24041 4641 24075 4675
rect 25120 4641 25154 4675
rect 11161 4573 11195 4607
rect 12081 4573 12115 4607
rect 12725 4573 12759 4607
rect 13645 4573 13679 4607
rect 18613 4573 18647 4607
rect 18889 4573 18923 4607
rect 8125 4505 8159 4539
rect 15853 4505 15887 4539
rect 25191 4505 25225 4539
rect 11529 4437 11563 4471
rect 14565 4437 14599 4471
rect 17693 4437 17727 4471
rect 24179 4437 24213 4471
rect 7067 4233 7101 4267
rect 13461 4233 13495 4267
rect 15485 4233 15519 4267
rect 17233 4233 17267 4267
rect 18521 4233 18555 4267
rect 20637 4233 20671 4267
rect 21741 4233 21775 4267
rect 22753 4233 22787 4267
rect 23121 4233 23155 4267
rect 24041 4233 24075 4267
rect 25145 4233 25179 4267
rect 7481 4165 7515 4199
rect 7849 4165 7883 4199
rect 14657 4165 14691 4199
rect 24731 4165 24765 4199
rect 6285 4097 6319 4131
rect 6837 4097 6871 4131
rect 8677 4097 8711 4131
rect 12173 4097 12207 4131
rect 12817 4097 12851 4131
rect 14105 4097 14139 4131
rect 16773 4097 16807 4131
rect 17877 4097 17911 4131
rect 18981 4097 19015 4131
rect 20177 4097 20211 4131
rect 25513 4097 25547 4131
rect 8585 4029 8619 4063
rect 9505 4029 9539 4063
rect 10149 4029 10183 4063
rect 10517 4029 10551 4063
rect 10885 4029 10919 4063
rect 20729 4029 20763 4063
rect 21005 4029 21039 4063
rect 22017 4029 22051 4063
rect 22328 4029 22362 4063
rect 24660 4029 24694 4063
rect 25672 4029 25706 4063
rect 26065 4029 26099 4063
rect 6561 3961 6595 3995
rect 8953 3961 8987 3995
rect 10977 3961 11011 3995
rect 12541 3961 12575 3995
rect 12633 3961 12667 3995
rect 13921 3961 13955 3995
rect 14197 3961 14231 3995
rect 15117 3961 15151 3995
rect 15669 3961 15703 3995
rect 15761 3961 15795 3995
rect 16313 3961 16347 3995
rect 19302 3961 19336 3995
rect 9413 3893 9447 3927
rect 11253 3893 11287 3927
rect 11621 3893 11655 3927
rect 18797 3893 18831 3927
rect 19901 3893 19935 3927
rect 22017 3893 22051 3927
rect 22109 3893 22143 3927
rect 22431 3893 22465 3927
rect 25743 3893 25777 3927
rect 7757 3689 7791 3723
rect 16773 3689 16807 3723
rect 17969 3689 18003 3723
rect 19073 3689 19107 3723
rect 19993 3689 20027 3723
rect 24639 3689 24673 3723
rect 9045 3621 9079 3655
rect 9413 3621 9447 3655
rect 13737 3621 13771 3655
rect 15485 3621 15519 3655
rect 16037 3621 16071 3655
rect 20729 3621 20763 3655
rect 21005 3621 21039 3655
rect 21097 3621 21131 3655
rect 22017 3621 22051 3655
rect 6929 3553 6963 3587
rect 8217 3553 8251 3587
rect 9689 3553 9723 3587
rect 10425 3553 10459 3587
rect 10609 3553 10643 3587
rect 11069 3553 11103 3587
rect 11989 3553 12023 3587
rect 13461 3553 13495 3587
rect 14381 3553 14415 3587
rect 19349 3553 19383 3587
rect 22477 3553 22511 3587
rect 23556 3553 23590 3587
rect 24568 3553 24602 3587
rect 5917 3485 5951 3519
rect 11161 3485 11195 3519
rect 15393 3485 15427 3519
rect 17601 3485 17635 3519
rect 21649 3485 21683 3519
rect 7113 3417 7147 3451
rect 12173 3417 12207 3451
rect 22615 3417 22649 3451
rect 8033 3349 8067 3383
rect 8401 3349 8435 3383
rect 11437 3349 11471 3383
rect 11805 3349 11839 3383
rect 12633 3349 12667 3383
rect 12909 3349 12943 3383
rect 13277 3349 13311 3383
rect 14657 3349 14691 3383
rect 15117 3349 15151 3383
rect 16497 3349 16531 3383
rect 18521 3349 18555 3383
rect 19533 3349 19567 3383
rect 23627 3349 23661 3383
rect 7021 3145 7055 3179
rect 8861 3145 8895 3179
rect 9229 3145 9263 3179
rect 11437 3145 11471 3179
rect 11989 3145 12023 3179
rect 15485 3145 15519 3179
rect 15945 3145 15979 3179
rect 17601 3145 17635 3179
rect 18429 3145 18463 3179
rect 19993 3145 20027 3179
rect 21557 3145 21591 3179
rect 24823 3145 24857 3179
rect 6285 3077 6319 3111
rect 13369 3077 13403 3111
rect 19165 3077 19199 3111
rect 22661 3077 22695 3111
rect 24133 3077 24167 3111
rect 4721 3009 4755 3043
rect 11069 3009 11103 3043
rect 16497 3009 16531 3043
rect 17141 3009 17175 3043
rect 18613 3009 18647 3043
rect 19533 3009 19567 3043
rect 20453 3009 20487 3043
rect 21741 3009 21775 3043
rect 22017 3009 22051 3043
rect 5800 2941 5834 2975
rect 6653 2941 6687 2975
rect 7849 2941 7883 2975
rect 9321 2941 9355 2975
rect 9873 2941 9907 2975
rect 10333 2941 10367 2975
rect 10701 2941 10735 2975
rect 12449 2941 12483 2975
rect 14289 2941 14323 2975
rect 15209 2941 15243 2975
rect 23397 2941 23431 2975
rect 23581 2941 23615 2975
rect 24752 2941 24786 2975
rect 25145 2941 25179 2975
rect 8493 2873 8527 2907
rect 10793 2873 10827 2907
rect 12770 2873 12804 2907
rect 13645 2873 13679 2907
rect 14105 2873 14139 2907
rect 14610 2873 14644 2907
rect 16313 2873 16347 2907
rect 16589 2873 16623 2907
rect 18705 2873 18739 2907
rect 20177 2873 20211 2907
rect 20269 2873 20303 2907
rect 21833 2873 21867 2907
rect 5871 2805 5905 2839
rect 7665 2805 7699 2839
rect 21097 2805 21131 2839
rect 23811 2805 23845 2839
rect 24593 2805 24627 2839
rect 5963 2601 5997 2635
rect 7941 2601 7975 2635
rect 13001 2601 13035 2635
rect 14197 2601 14231 2635
rect 14565 2601 14599 2635
rect 15209 2601 15243 2635
rect 17601 2601 17635 2635
rect 18797 2601 18831 2635
rect 20177 2601 20211 2635
rect 23397 2601 23431 2635
rect 25191 2601 25225 2635
rect 6745 2533 6779 2567
rect 8861 2533 8895 2567
rect 10654 2533 10688 2567
rect 11621 2533 11655 2567
rect 13369 2533 13403 2567
rect 15669 2533 15703 2567
rect 18153 2533 18187 2567
rect 19073 2533 19107 2567
rect 20637 2533 20671 2567
rect 21281 2533 21315 2567
rect 21373 2533 21407 2567
rect 4880 2465 4914 2499
rect 5860 2465 5894 2499
rect 6285 2465 6319 2499
rect 6929 2465 6963 2499
rect 7389 2465 7423 2499
rect 8217 2465 8251 2499
rect 9321 2465 9355 2499
rect 10149 2465 10183 2499
rect 10333 2465 10367 2499
rect 11897 2465 11931 2499
rect 17049 2465 17083 2499
rect 22753 2465 22787 2499
rect 24076 2465 24110 2499
rect 24501 2465 24535 2499
rect 25088 2465 25122 2499
rect 5365 2397 5399 2431
rect 13277 2397 13311 2431
rect 15577 2397 15611 2431
rect 16497 2397 16531 2431
rect 18981 2397 19015 2431
rect 19257 2397 19291 2431
rect 21005 2397 21039 2431
rect 24179 2397 24213 2431
rect 4951 2329 4985 2363
rect 7389 2329 7423 2363
rect 7573 2329 7607 2363
rect 12357 2329 12391 2363
rect 13829 2329 13863 2363
rect 16129 2329 16163 2363
rect 17233 2329 17267 2363
rect 21833 2329 21867 2363
rect 25513 2329 25547 2363
rect 7113 2261 7147 2295
rect 11253 2261 11287 2295
rect 16865 2261 16899 2295
rect 22937 2261 22971 2295
<< metal1 >>
rect 14 27480 20 27532
rect 72 27520 78 27532
rect 658 27520 664 27532
rect 72 27492 664 27520
rect 72 27480 78 27492
rect 658 27480 664 27492
rect 716 27480 722 27532
rect 2774 27480 2780 27532
rect 2832 27520 2838 27532
rect 3418 27520 3424 27532
rect 2832 27492 3424 27520
rect 2832 27480 2838 27492
rect 3418 27480 3424 27492
rect 3476 27480 3482 27532
rect 19518 27480 19524 27532
rect 19576 27520 19582 27532
rect 21634 27520 21640 27532
rect 19576 27492 21640 27520
rect 19576 27480 19582 27492
rect 21634 27480 21640 27492
rect 21692 27480 21698 27532
rect 22462 27480 22468 27532
rect 22520 27520 22526 27532
rect 23014 27520 23020 27532
rect 22520 27492 23020 27520
rect 22520 27480 22526 27492
rect 23014 27480 23020 27492
rect 23072 27480 23078 27532
rect 24854 27480 24860 27532
rect 24912 27520 24918 27532
rect 25774 27520 25780 27532
rect 24912 27492 25780 27520
rect 24912 27480 24918 27492
rect 25774 27480 25780 27492
rect 25832 27480 25838 27532
rect 26234 27480 26240 27532
rect 26292 27520 26298 27532
rect 27154 27520 27160 27532
rect 26292 27492 27160 27520
rect 26292 27480 26298 27492
rect 27154 27480 27160 27492
rect 27212 27480 27218 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 17773 24395 17831 24401
rect 17773 24361 17785 24395
rect 17819 24392 17831 24395
rect 18782 24392 18788 24404
rect 17819 24364 18788 24392
rect 17819 24361 17831 24364
rect 17773 24355 17831 24361
rect 18782 24352 18788 24364
rect 18840 24352 18846 24404
rect 10778 24216 10784 24268
rect 10836 24256 10842 24268
rect 17586 24256 17592 24268
rect 10836 24228 17592 24256
rect 10836 24216 10842 24228
rect 17586 24216 17592 24228
rect 17644 24216 17650 24268
rect 23201 24259 23259 24265
rect 23201 24225 23213 24259
rect 23247 24256 23259 24259
rect 23290 24256 23296 24268
rect 23247 24228 23296 24256
rect 23247 24225 23259 24228
rect 23201 24219 23259 24225
rect 23290 24216 23296 24228
rect 23348 24216 23354 24268
rect 22922 24012 22928 24064
rect 22980 24052 22986 24064
rect 23431 24055 23489 24061
rect 23431 24052 23443 24055
rect 22980 24024 23443 24052
rect 22980 24012 22986 24024
rect 23431 24021 23443 24024
rect 23477 24021 23489 24055
rect 23431 24015 23489 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 6178 23808 6184 23860
rect 6236 23848 6242 23860
rect 7009 23851 7067 23857
rect 7009 23848 7021 23851
rect 6236 23820 7021 23848
rect 6236 23808 6242 23820
rect 7009 23817 7021 23820
rect 7055 23817 7067 23851
rect 7009 23811 7067 23817
rect 12621 23851 12679 23857
rect 12621 23817 12633 23851
rect 12667 23848 12679 23851
rect 13170 23848 13176 23860
rect 12667 23820 13176 23848
rect 12667 23817 12679 23820
rect 12621 23811 12679 23817
rect 13170 23808 13176 23820
rect 13228 23808 13234 23860
rect 14277 23851 14335 23857
rect 14277 23817 14289 23851
rect 14323 23848 14335 23851
rect 14642 23848 14648 23860
rect 14323 23820 14648 23848
rect 14323 23817 14335 23820
rect 14277 23811 14335 23817
rect 14642 23808 14648 23820
rect 14700 23808 14706 23860
rect 16117 23851 16175 23857
rect 16117 23817 16129 23851
rect 16163 23848 16175 23851
rect 17402 23848 17408 23860
rect 16163 23820 17408 23848
rect 16163 23817 16175 23820
rect 16117 23811 16175 23817
rect 17402 23808 17408 23820
rect 17460 23808 17466 23860
rect 17586 23848 17592 23860
rect 17547 23820 17592 23848
rect 17586 23808 17592 23820
rect 17644 23808 17650 23860
rect 18601 23851 18659 23857
rect 18601 23817 18613 23851
rect 18647 23848 18659 23851
rect 20162 23848 20168 23860
rect 18647 23820 20168 23848
rect 18647 23817 18659 23820
rect 18601 23811 18659 23817
rect 20162 23808 20168 23820
rect 20220 23808 20226 23860
rect 23290 23848 23296 23860
rect 23251 23820 23296 23848
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 25130 23848 25136 23860
rect 25091 23820 25136 23848
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 22465 23783 22523 23789
rect 22465 23749 22477 23783
rect 22511 23780 22523 23783
rect 24210 23780 24216 23792
rect 22511 23752 24216 23780
rect 22511 23749 22523 23752
rect 22465 23743 22523 23749
rect 1535 23715 1593 23721
rect 1535 23681 1547 23715
rect 1581 23712 1593 23715
rect 8018 23712 8024 23724
rect 1581 23684 8024 23712
rect 1581 23681 1593 23684
rect 1535 23675 1593 23681
rect 8018 23672 8024 23684
rect 8076 23672 8082 23724
rect 1210 23604 1216 23656
rect 1268 23644 1274 23656
rect 1432 23647 1490 23653
rect 1432 23644 1444 23647
rect 1268 23616 1444 23644
rect 1268 23604 1274 23616
rect 1432 23613 1444 23616
rect 1478 23644 1490 23647
rect 1857 23647 1915 23653
rect 1857 23644 1869 23647
rect 1478 23616 1869 23644
rect 1478 23613 1490 23616
rect 1432 23607 1490 23613
rect 1857 23613 1869 23616
rect 1903 23613 1915 23647
rect 1857 23607 1915 23613
rect 4316 23647 4374 23653
rect 4316 23613 4328 23647
rect 4362 23644 4374 23647
rect 4706 23644 4712 23656
rect 4362 23616 4712 23644
rect 4362 23613 4374 23616
rect 4316 23607 4374 23613
rect 4706 23604 4712 23616
rect 4764 23604 4770 23656
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23644 6883 23647
rect 12434 23644 12440 23656
rect 6871 23616 7512 23644
rect 12347 23616 12440 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 4062 23468 4068 23520
rect 4120 23508 4126 23520
rect 7484 23517 7512 23616
rect 12434 23604 12440 23616
rect 12492 23644 12498 23656
rect 12989 23647 13047 23653
rect 12989 23644 13001 23647
rect 12492 23616 13001 23644
rect 12492 23604 12498 23616
rect 12989 23613 13001 23616
rect 13035 23613 13047 23647
rect 12989 23607 13047 23613
rect 14093 23647 14151 23653
rect 14093 23613 14105 23647
rect 14139 23644 14151 23647
rect 15930 23644 15936 23656
rect 14139 23616 14780 23644
rect 15891 23616 15936 23644
rect 14139 23613 14151 23616
rect 14093 23607 14151 23613
rect 4387 23511 4445 23517
rect 4387 23508 4399 23511
rect 4120 23480 4399 23508
rect 4120 23468 4126 23480
rect 4387 23477 4399 23480
rect 4433 23477 4445 23511
rect 4387 23471 4445 23477
rect 7469 23511 7527 23517
rect 7469 23477 7481 23511
rect 7515 23508 7527 23511
rect 7742 23508 7748 23520
rect 7515 23480 7748 23508
rect 7515 23477 7527 23480
rect 7469 23471 7527 23477
rect 7742 23468 7748 23480
rect 7800 23468 7806 23520
rect 14752 23517 14780 23616
rect 15930 23604 15936 23616
rect 15988 23644 15994 23656
rect 16485 23647 16543 23653
rect 16485 23644 16497 23647
rect 15988 23616 16497 23644
rect 15988 23604 15994 23616
rect 16485 23613 16497 23616
rect 16531 23644 16543 23647
rect 16942 23644 16948 23656
rect 16531 23616 16948 23644
rect 16531 23613 16543 23616
rect 16485 23607 16543 23613
rect 16942 23604 16948 23616
rect 17000 23604 17006 23656
rect 17218 23604 17224 23656
rect 17276 23644 17282 23656
rect 22623 23653 22651 23752
rect 24210 23740 24216 23752
rect 24268 23740 24274 23792
rect 18417 23647 18475 23653
rect 18417 23644 18429 23647
rect 17276 23616 18429 23644
rect 17276 23604 17282 23616
rect 18417 23613 18429 23616
rect 18463 23644 18475 23647
rect 18969 23647 19027 23653
rect 18969 23644 18981 23647
rect 18463 23616 18981 23644
rect 18463 23613 18475 23616
rect 18417 23607 18475 23613
rect 18969 23613 18981 23616
rect 19015 23613 19027 23647
rect 18969 23607 19027 23613
rect 22608 23647 22666 23653
rect 22608 23613 22620 23647
rect 22654 23613 22666 23647
rect 22608 23607 22666 23613
rect 24632 23647 24690 23653
rect 24632 23613 24644 23647
rect 24678 23644 24690 23647
rect 25130 23644 25136 23656
rect 24678 23616 25136 23644
rect 24678 23613 24690 23616
rect 24632 23607 24690 23613
rect 25130 23604 25136 23616
rect 25188 23604 25194 23656
rect 21450 23536 21456 23588
rect 21508 23576 21514 23588
rect 22695 23579 22753 23585
rect 22695 23576 22707 23579
rect 21508 23548 22707 23576
rect 21508 23536 21514 23548
rect 22695 23545 22707 23548
rect 22741 23545 22753 23579
rect 22695 23539 22753 23545
rect 22830 23536 22836 23588
rect 22888 23576 22894 23588
rect 24719 23579 24777 23585
rect 24719 23576 24731 23579
rect 22888 23548 24731 23576
rect 22888 23536 22894 23548
rect 24719 23545 24731 23548
rect 24765 23545 24777 23579
rect 24719 23539 24777 23545
rect 14737 23511 14795 23517
rect 14737 23477 14749 23511
rect 14783 23508 14795 23511
rect 14826 23508 14832 23520
rect 14783 23480 14832 23508
rect 14783 23477 14795 23480
rect 14737 23471 14795 23477
rect 14826 23468 14832 23480
rect 14884 23468 14890 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 106 23264 112 23316
rect 164 23304 170 23316
rect 1581 23307 1639 23313
rect 1581 23304 1593 23307
rect 164 23276 1593 23304
rect 164 23264 170 23276
rect 1581 23273 1593 23276
rect 1627 23273 1639 23307
rect 1581 23267 1639 23273
rect 1394 23168 1400 23180
rect 1355 23140 1400 23168
rect 1394 23128 1400 23140
rect 1452 23128 1458 23180
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 25130 22760 25136 22772
rect 25091 22732 25136 22760
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 11974 22652 11980 22704
rect 12032 22692 12038 22704
rect 12434 22692 12440 22704
rect 12032 22664 12440 22692
rect 12032 22652 12038 22664
rect 12434 22652 12440 22664
rect 12492 22652 12498 22704
rect 1394 22516 1400 22568
rect 1452 22556 1458 22568
rect 1673 22559 1731 22565
rect 1673 22556 1685 22559
rect 1452 22528 1685 22556
rect 1452 22516 1458 22528
rect 1673 22525 1685 22528
rect 1719 22556 1731 22559
rect 11974 22556 11980 22568
rect 1719 22528 11980 22556
rect 1719 22525 1731 22528
rect 1673 22519 1731 22525
rect 11974 22516 11980 22528
rect 12032 22516 12038 22568
rect 24648 22559 24706 22565
rect 24648 22525 24660 22559
rect 24694 22556 24706 22559
rect 25130 22556 25136 22568
rect 24694 22528 25136 22556
rect 24694 22525 24706 22528
rect 24648 22519 24706 22525
rect 25130 22516 25136 22528
rect 25188 22516 25194 22568
rect 22002 22380 22008 22432
rect 22060 22420 22066 22432
rect 24719 22423 24777 22429
rect 24719 22420 24731 22423
rect 22060 22392 24731 22420
rect 22060 22380 22066 22392
rect 24719 22389 24731 22392
rect 24765 22389 24777 22423
rect 24719 22383 24777 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 24581 20995 24639 21001
rect 24581 20961 24593 20995
rect 24627 20992 24639 20995
rect 24670 20992 24676 21004
rect 24627 20964 24676 20992
rect 24627 20961 24639 20964
rect 24581 20955 24639 20961
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 18598 20748 18604 20800
rect 18656 20788 18662 20800
rect 24719 20791 24777 20797
rect 24719 20788 24731 20791
rect 18656 20760 24731 20788
rect 18656 20748 18662 20760
rect 24719 20757 24731 20760
rect 24765 20757 24777 20791
rect 24719 20751 24777 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 24670 20584 24676 20596
rect 24631 20556 24676 20584
rect 24670 20544 24676 20556
rect 24728 20544 24734 20596
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19904 11943 19907
rect 12066 19904 12072 19916
rect 11931 19876 12072 19904
rect 11931 19873 11943 19876
rect 11885 19867 11943 19873
rect 12066 19864 12072 19876
rect 12124 19864 12130 19916
rect 11606 19660 11612 19712
rect 11664 19700 11670 19712
rect 12115 19703 12173 19709
rect 12115 19700 12127 19703
rect 11664 19672 12127 19700
rect 11664 19660 11670 19672
rect 12115 19669 12127 19672
rect 12161 19669 12173 19703
rect 13906 19700 13912 19712
rect 13867 19672 13912 19700
rect 12115 19663 12173 19669
rect 13906 19660 13912 19672
rect 13964 19660 13970 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 14826 19456 14832 19508
rect 14884 19496 14890 19508
rect 15519 19499 15577 19505
rect 15519 19496 15531 19499
rect 14884 19468 15531 19496
rect 14884 19456 14890 19468
rect 15519 19465 15531 19468
rect 15565 19465 15577 19499
rect 15519 19459 15577 19465
rect 11330 19360 11336 19372
rect 11291 19332 11336 19360
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 13906 19320 13912 19372
rect 13964 19360 13970 19372
rect 17678 19360 17684 19372
rect 13964 19332 17684 19360
rect 13964 19320 13970 19332
rect 10940 19295 10998 19301
rect 10940 19261 10952 19295
rect 10986 19292 10998 19295
rect 11348 19292 11376 19320
rect 14108 19301 14136 19332
rect 17678 19320 17684 19332
rect 17736 19320 17742 19372
rect 10986 19264 11376 19292
rect 12564 19295 12622 19301
rect 10986 19261 10998 19264
rect 10940 19255 10998 19261
rect 12564 19261 12576 19295
rect 12610 19292 12622 19295
rect 12989 19295 13047 19301
rect 12989 19292 13001 19295
rect 12610 19264 13001 19292
rect 12610 19261 12622 19264
rect 12564 19255 12622 19261
rect 12989 19261 13001 19264
rect 13035 19261 13047 19295
rect 12989 19255 13047 19261
rect 14093 19295 14151 19301
rect 14093 19261 14105 19295
rect 14139 19261 14151 19295
rect 14093 19255 14151 19261
rect 14277 19295 14335 19301
rect 14277 19261 14289 19295
rect 14323 19261 14335 19295
rect 14277 19255 14335 19261
rect 15448 19295 15506 19301
rect 15448 19261 15460 19295
rect 15494 19292 15506 19295
rect 15838 19292 15844 19304
rect 15494 19264 15844 19292
rect 15494 19261 15506 19264
rect 15448 19255 15506 19261
rect 8570 19184 8576 19236
rect 8628 19224 8634 19236
rect 12579 19224 12607 19255
rect 8628 19196 12607 19224
rect 12667 19227 12725 19233
rect 8628 19184 8634 19196
rect 12667 19193 12679 19227
rect 12713 19224 12725 19227
rect 13538 19224 13544 19236
rect 12713 19196 13544 19224
rect 12713 19193 12725 19196
rect 12667 19187 12725 19193
rect 13538 19184 13544 19196
rect 13596 19184 13602 19236
rect 14292 19224 14320 19255
rect 15838 19252 15844 19264
rect 15896 19252 15902 19304
rect 13786 19196 14320 19224
rect 14553 19227 14611 19233
rect 10870 19116 10876 19168
rect 10928 19156 10934 19168
rect 11011 19159 11069 19165
rect 11011 19156 11023 19159
rect 10928 19128 11023 19156
rect 10928 19116 10934 19128
rect 11011 19125 11023 19128
rect 11057 19125 11069 19159
rect 12066 19156 12072 19168
rect 12027 19128 12072 19156
rect 11011 19119 11069 19125
rect 12066 19116 12072 19128
rect 12124 19116 12130 19168
rect 12894 19116 12900 19168
rect 12952 19156 12958 19168
rect 13633 19159 13691 19165
rect 13633 19156 13645 19159
rect 12952 19128 13645 19156
rect 12952 19116 12958 19128
rect 13633 19125 13645 19128
rect 13679 19156 13691 19159
rect 13786 19156 13814 19196
rect 14553 19193 14565 19227
rect 14599 19224 14611 19227
rect 14826 19224 14832 19236
rect 14599 19196 14832 19224
rect 14599 19193 14611 19196
rect 14553 19187 14611 19193
rect 14826 19184 14832 19196
rect 14884 19184 14890 19236
rect 13679 19128 13814 19156
rect 13679 19125 13691 19128
rect 13633 19119 13691 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 10870 18952 10876 18964
rect 10831 18924 10876 18952
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 12066 18912 12072 18964
rect 12124 18952 12130 18964
rect 16758 18952 16764 18964
rect 12124 18924 16764 18952
rect 12124 18912 12130 18924
rect 16758 18912 16764 18924
rect 16816 18912 16822 18964
rect 9858 18884 9864 18896
rect 9819 18856 9864 18884
rect 9858 18844 9864 18856
rect 9916 18844 9922 18896
rect 13722 18844 13728 18896
rect 13780 18884 13786 18896
rect 13817 18887 13875 18893
rect 13817 18884 13829 18887
rect 13780 18856 13829 18884
rect 13780 18844 13786 18856
rect 13817 18853 13829 18856
rect 13863 18853 13875 18887
rect 15562 18884 15568 18896
rect 15523 18856 15568 18884
rect 13817 18847 13875 18853
rect 15562 18844 15568 18856
rect 15620 18844 15626 18896
rect 8481 18819 8539 18825
rect 8481 18785 8493 18819
rect 8527 18816 8539 18819
rect 8570 18816 8576 18828
rect 8527 18788 8576 18816
rect 8527 18785 8539 18788
rect 8481 18779 8539 18785
rect 8570 18776 8576 18788
rect 8628 18776 8634 18828
rect 11330 18776 11336 18828
rect 11388 18816 11394 18828
rect 12158 18816 12164 18828
rect 11388 18788 12164 18816
rect 11388 18776 11394 18788
rect 12158 18776 12164 18788
rect 12216 18816 12222 18828
rect 21542 18825 21548 18828
rect 12380 18819 12438 18825
rect 12380 18816 12392 18819
rect 12216 18788 12392 18816
rect 12216 18776 12222 18788
rect 12380 18785 12392 18788
rect 12426 18785 12438 18819
rect 21520 18819 21548 18825
rect 21520 18816 21532 18819
rect 21455 18788 21532 18816
rect 12380 18779 12438 18785
rect 21520 18785 21532 18788
rect 21600 18816 21606 18828
rect 22094 18816 22100 18828
rect 21600 18788 22100 18816
rect 21520 18779 21548 18785
rect 21542 18776 21548 18779
rect 21600 18776 21606 18788
rect 22094 18776 22100 18788
rect 22152 18776 22158 18828
rect 8711 18751 8769 18757
rect 8711 18717 8723 18751
rect 8757 18748 8769 18751
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 8757 18720 9781 18748
rect 8757 18717 8769 18720
rect 8711 18711 8769 18717
rect 9769 18717 9781 18720
rect 9815 18748 9827 18751
rect 10226 18748 10232 18760
rect 9815 18720 10232 18748
rect 9815 18717 9827 18720
rect 9769 18711 9827 18717
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 11238 18748 11244 18760
rect 11199 18720 11244 18748
rect 11238 18708 11244 18720
rect 11296 18708 11302 18760
rect 13725 18751 13783 18757
rect 13725 18717 13737 18751
rect 13771 18717 13783 18751
rect 13725 18711 13783 18717
rect 14369 18751 14427 18757
rect 14369 18717 14381 18751
rect 14415 18748 14427 18751
rect 14550 18748 14556 18760
rect 14415 18720 14556 18748
rect 14415 18717 14427 18720
rect 14369 18711 14427 18717
rect 10042 18640 10048 18692
rect 10100 18680 10106 18692
rect 10321 18683 10379 18689
rect 10321 18680 10333 18683
rect 10100 18652 10333 18680
rect 10100 18640 10106 18652
rect 10321 18649 10333 18652
rect 10367 18649 10379 18683
rect 10321 18643 10379 18649
rect 12483 18683 12541 18689
rect 12483 18649 12495 18683
rect 12529 18680 12541 18683
rect 13449 18683 13507 18689
rect 13449 18680 13461 18683
rect 12529 18652 13461 18680
rect 12529 18649 12541 18652
rect 12483 18643 12541 18649
rect 13449 18649 13461 18652
rect 13495 18680 13507 18683
rect 13740 18680 13768 18711
rect 14550 18708 14556 18720
rect 14608 18708 14614 18760
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18748 15531 18751
rect 15654 18748 15660 18760
rect 15519 18720 15660 18748
rect 15519 18717 15531 18720
rect 15473 18711 15531 18717
rect 15654 18708 15660 18720
rect 15712 18708 15718 18760
rect 16114 18748 16120 18760
rect 16075 18720 16120 18748
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 13495 18652 13768 18680
rect 13495 18649 13507 18652
rect 13449 18643 13507 18649
rect 12802 18612 12808 18624
rect 12763 18584 12808 18612
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 21591 18615 21649 18621
rect 21591 18581 21603 18615
rect 21637 18612 21649 18615
rect 22646 18612 22652 18624
rect 21637 18584 22652 18612
rect 21637 18581 21649 18584
rect 21591 18575 21649 18581
rect 22646 18572 22652 18584
rect 22704 18572 22710 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 7742 18408 7748 18420
rect 7703 18380 7748 18408
rect 7742 18368 7748 18380
rect 7800 18368 7806 18420
rect 8570 18408 8576 18420
rect 8531 18380 8576 18408
rect 8570 18368 8576 18380
rect 8628 18368 8634 18420
rect 10226 18408 10232 18420
rect 10187 18380 10232 18408
rect 10226 18368 10232 18380
rect 10284 18368 10290 18420
rect 12158 18408 12164 18420
rect 12119 18380 12164 18408
rect 12158 18368 12164 18380
rect 12216 18368 12222 18420
rect 21542 18408 21548 18420
rect 21503 18380 21548 18408
rect 21542 18368 21548 18380
rect 21600 18368 21606 18420
rect 22462 18408 22468 18420
rect 22423 18380 22468 18408
rect 22462 18368 22468 18380
rect 22520 18368 22526 18420
rect 13722 18300 13728 18352
rect 13780 18340 13786 18352
rect 15381 18343 15439 18349
rect 15381 18340 15393 18343
rect 13780 18312 15393 18340
rect 13780 18300 13786 18312
rect 15381 18309 15393 18312
rect 15427 18340 15439 18343
rect 15562 18340 15568 18352
rect 15427 18312 15568 18340
rect 15427 18309 15439 18312
rect 15381 18303 15439 18309
rect 15562 18300 15568 18312
rect 15620 18300 15626 18352
rect 15654 18300 15660 18352
rect 15712 18340 15718 18352
rect 17221 18343 17279 18349
rect 17221 18340 17233 18343
rect 15712 18312 17233 18340
rect 15712 18300 15718 18312
rect 17221 18309 17233 18312
rect 17267 18340 17279 18343
rect 21450 18340 21456 18352
rect 17267 18312 21456 18340
rect 17267 18309 17279 18312
rect 17221 18303 17279 18309
rect 21450 18300 21456 18312
rect 21508 18300 21514 18352
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 8941 18275 8999 18281
rect 8941 18272 8953 18275
rect 8076 18244 8953 18272
rect 8076 18232 8082 18244
rect 8941 18241 8953 18244
rect 8987 18272 8999 18275
rect 9030 18272 9036 18284
rect 8987 18244 9036 18272
rect 8987 18241 8999 18244
rect 8941 18235 8999 18241
rect 9030 18232 9036 18244
rect 9088 18232 9094 18284
rect 10870 18272 10876 18284
rect 10831 18244 10876 18272
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 14550 18272 14556 18284
rect 14511 18244 14556 18272
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 15841 18275 15899 18281
rect 15841 18241 15853 18275
rect 15887 18272 15899 18275
rect 15930 18272 15936 18284
rect 15887 18244 15936 18272
rect 15887 18241 15899 18244
rect 15841 18235 15899 18241
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 16114 18272 16120 18284
rect 16075 18244 16120 18272
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 7469 18207 7527 18213
rect 7469 18173 7481 18207
rect 7515 18204 7527 18207
rect 7596 18207 7654 18213
rect 7596 18204 7608 18207
rect 7515 18176 7608 18204
rect 7515 18173 7527 18176
rect 7469 18167 7527 18173
rect 7596 18173 7608 18176
rect 7642 18204 7654 18207
rect 8754 18204 8760 18216
rect 7642 18176 8760 18204
rect 7642 18173 7654 18176
rect 7596 18167 7654 18173
rect 8754 18164 8760 18176
rect 8812 18164 8818 18216
rect 12802 18204 12808 18216
rect 12763 18176 12808 18204
rect 12802 18164 12808 18176
rect 12860 18164 12866 18216
rect 12894 18164 12900 18216
rect 12952 18204 12958 18216
rect 19518 18213 19524 18216
rect 13081 18207 13139 18213
rect 13081 18204 13093 18207
rect 12952 18176 13093 18204
rect 12952 18164 12958 18176
rect 13081 18173 13093 18176
rect 13127 18173 13139 18207
rect 19496 18207 19524 18213
rect 19496 18204 19508 18207
rect 19431 18176 19508 18204
rect 13081 18167 13139 18173
rect 19496 18173 19508 18176
rect 19576 18204 19582 18216
rect 19889 18207 19947 18213
rect 19889 18204 19901 18207
rect 19576 18176 19901 18204
rect 19496 18167 19524 18173
rect 19518 18164 19524 18167
rect 19576 18164 19582 18176
rect 19889 18173 19901 18176
rect 19935 18173 19947 18207
rect 19889 18167 19947 18173
rect 22072 18207 22130 18213
rect 22072 18173 22084 18207
rect 22118 18204 22130 18207
rect 22462 18204 22468 18216
rect 22118 18176 22468 18204
rect 22118 18173 22130 18176
rect 22072 18167 22130 18173
rect 22462 18164 22468 18176
rect 22520 18164 22526 18216
rect 9033 18139 9091 18145
rect 9033 18136 9045 18139
rect 8220 18108 9045 18136
rect 8220 18080 8248 18108
rect 9033 18105 9045 18108
rect 9079 18105 9091 18139
rect 9582 18136 9588 18148
rect 9543 18108 9588 18136
rect 9033 18099 9091 18105
rect 8202 18068 8208 18080
rect 8163 18040 8208 18068
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 9048 18068 9076 18099
rect 9582 18096 9588 18108
rect 9640 18096 9646 18148
rect 10689 18139 10747 18145
rect 10689 18105 10701 18139
rect 10735 18136 10747 18139
rect 10962 18136 10968 18148
rect 10735 18108 10968 18136
rect 10735 18105 10747 18108
rect 10689 18099 10747 18105
rect 10962 18096 10968 18108
rect 11020 18096 11026 18148
rect 11517 18139 11575 18145
rect 11517 18105 11529 18139
rect 11563 18136 11575 18139
rect 11882 18136 11888 18148
rect 11563 18108 11888 18136
rect 11563 18105 11575 18108
rect 11517 18099 11575 18105
rect 11882 18096 11888 18108
rect 11940 18096 11946 18148
rect 13354 18136 13360 18148
rect 13315 18108 13360 18136
rect 13354 18096 13360 18108
rect 13412 18096 13418 18148
rect 14274 18136 14280 18148
rect 14235 18108 14280 18136
rect 14274 18096 14280 18108
rect 14332 18096 14338 18148
rect 14369 18139 14427 18145
rect 14369 18105 14381 18139
rect 14415 18105 14427 18139
rect 14369 18099 14427 18105
rect 15933 18139 15991 18145
rect 15933 18105 15945 18139
rect 15979 18105 15991 18139
rect 15933 18099 15991 18105
rect 19705 18139 19763 18145
rect 19705 18105 19717 18139
rect 19751 18136 19763 18139
rect 20530 18136 20536 18148
rect 19751 18108 20536 18136
rect 19751 18105 19763 18108
rect 19705 18099 19763 18105
rect 9490 18068 9496 18080
rect 9048 18040 9496 18068
rect 9490 18028 9496 18040
rect 9548 18068 9554 18080
rect 9858 18068 9864 18080
rect 9548 18040 9864 18068
rect 9548 18028 9554 18040
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 13722 18068 13728 18080
rect 13683 18040 13728 18068
rect 13722 18028 13728 18040
rect 13780 18028 13786 18080
rect 14093 18071 14151 18077
rect 14093 18037 14105 18071
rect 14139 18068 14151 18071
rect 14384 18068 14412 18099
rect 15378 18068 15384 18080
rect 14139 18040 15384 18068
rect 14139 18037 14151 18040
rect 14093 18031 14151 18037
rect 15378 18028 15384 18040
rect 15436 18068 15442 18080
rect 15948 18068 15976 18099
rect 20530 18096 20536 18108
rect 20588 18096 20594 18148
rect 20625 18139 20683 18145
rect 20625 18105 20637 18139
rect 20671 18105 20683 18139
rect 20625 18099 20683 18105
rect 21177 18139 21235 18145
rect 21177 18105 21189 18139
rect 21223 18136 21235 18139
rect 21450 18136 21456 18148
rect 21223 18108 21456 18136
rect 21223 18105 21235 18108
rect 21177 18099 21235 18105
rect 16761 18071 16819 18077
rect 16761 18068 16773 18071
rect 15436 18040 16773 18068
rect 15436 18028 15442 18040
rect 16761 18037 16773 18040
rect 16807 18037 16819 18071
rect 16761 18031 16819 18037
rect 19426 18028 19432 18080
rect 19484 18068 19490 18080
rect 20257 18071 20315 18077
rect 20257 18068 20269 18071
rect 19484 18040 20269 18068
rect 19484 18028 19490 18040
rect 20257 18037 20269 18040
rect 20303 18068 20315 18071
rect 20640 18068 20668 18099
rect 21450 18096 21456 18108
rect 21508 18096 21514 18148
rect 20303 18040 20668 18068
rect 20303 18037 20315 18040
rect 20257 18031 20315 18037
rect 21082 18028 21088 18080
rect 21140 18068 21146 18080
rect 22143 18071 22201 18077
rect 22143 18068 22155 18071
rect 21140 18040 22155 18068
rect 21140 18028 21146 18040
rect 22143 18037 22155 18040
rect 22189 18037 22201 18071
rect 22143 18031 22201 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 9030 17864 9036 17876
rect 8991 17836 9036 17864
rect 9030 17824 9036 17836
rect 9088 17824 9094 17876
rect 11698 17824 11704 17876
rect 11756 17864 11762 17876
rect 11756 17836 11928 17864
rect 11756 17824 11762 17836
rect 7466 17756 7472 17808
rect 7524 17796 7530 17808
rect 8202 17796 8208 17808
rect 7524 17768 8208 17796
rect 7524 17756 7530 17768
rect 8202 17756 8208 17768
rect 8260 17756 8266 17808
rect 10321 17799 10379 17805
rect 10321 17765 10333 17799
rect 10367 17796 10379 17799
rect 10686 17796 10692 17808
rect 10367 17768 10692 17796
rect 10367 17765 10379 17768
rect 10321 17759 10379 17765
rect 10686 17756 10692 17768
rect 10744 17756 10750 17808
rect 11238 17756 11244 17808
rect 11296 17796 11302 17808
rect 11790 17796 11796 17808
rect 11296 17768 11796 17796
rect 11296 17756 11302 17768
rect 11790 17756 11796 17768
rect 11848 17756 11854 17808
rect 11900 17805 11928 17836
rect 13354 17824 13360 17876
rect 13412 17864 13418 17876
rect 14090 17864 14096 17876
rect 13412 17836 14096 17864
rect 13412 17824 13418 17836
rect 14090 17824 14096 17836
rect 14148 17864 14154 17876
rect 14277 17867 14335 17873
rect 14277 17864 14289 17867
rect 14148 17836 14289 17864
rect 14148 17824 14154 17836
rect 14277 17833 14289 17836
rect 14323 17833 14335 17867
rect 20530 17864 20536 17876
rect 20491 17836 20536 17864
rect 14277 17827 14335 17833
rect 20530 17824 20536 17836
rect 20588 17824 20594 17876
rect 24762 17864 24768 17876
rect 24723 17836 24768 17864
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 11885 17799 11943 17805
rect 11885 17765 11897 17799
rect 11931 17796 11943 17799
rect 13449 17799 13507 17805
rect 13449 17796 13461 17799
rect 11931 17768 13461 17796
rect 11931 17765 11943 17768
rect 11885 17759 11943 17765
rect 13449 17765 13461 17768
rect 13495 17765 13507 17799
rect 15470 17796 15476 17808
rect 15431 17768 15476 17796
rect 13449 17759 13507 17765
rect 15470 17756 15476 17768
rect 15528 17756 15534 17808
rect 19426 17796 19432 17808
rect 19387 17768 19432 17796
rect 19426 17756 19432 17768
rect 19484 17756 19490 17808
rect 21082 17796 21088 17808
rect 21043 17768 21088 17796
rect 21082 17756 21088 17768
rect 21140 17756 21146 17808
rect 21177 17799 21235 17805
rect 21177 17765 21189 17799
rect 21223 17796 21235 17799
rect 21542 17796 21548 17808
rect 21223 17768 21548 17796
rect 21223 17765 21235 17768
rect 21177 17759 21235 17765
rect 21542 17756 21548 17768
rect 21600 17756 21606 17808
rect 22646 17796 22652 17808
rect 22607 17768 22652 17796
rect 22646 17756 22652 17768
rect 22704 17756 22710 17808
rect 22741 17799 22799 17805
rect 22741 17765 22753 17799
rect 22787 17796 22799 17799
rect 23106 17796 23112 17808
rect 22787 17768 23112 17796
rect 22787 17765 22799 17768
rect 22741 17759 22799 17765
rect 23106 17756 23112 17768
rect 23164 17756 23170 17808
rect 17678 17728 17684 17740
rect 17639 17700 17684 17728
rect 17678 17688 17684 17700
rect 17736 17688 17742 17740
rect 17954 17688 17960 17740
rect 18012 17728 18018 17740
rect 18141 17731 18199 17737
rect 18141 17728 18153 17731
rect 18012 17700 18153 17728
rect 18012 17688 18018 17700
rect 18141 17697 18153 17700
rect 18187 17697 18199 17731
rect 18141 17691 18199 17697
rect 24210 17688 24216 17740
rect 24268 17728 24274 17740
rect 24581 17731 24639 17737
rect 24581 17728 24593 17731
rect 24268 17700 24593 17728
rect 24268 17688 24274 17700
rect 24581 17697 24593 17700
rect 24627 17697 24639 17731
rect 24581 17691 24639 17697
rect 8110 17660 8116 17672
rect 8071 17632 8116 17660
rect 8110 17620 8116 17632
rect 8168 17620 8174 17672
rect 10042 17660 10048 17672
rect 9955 17632 10048 17660
rect 10042 17620 10048 17632
rect 10100 17660 10106 17672
rect 10229 17663 10287 17669
rect 10229 17660 10241 17663
rect 10100 17632 10241 17660
rect 10100 17620 10106 17632
rect 10229 17629 10241 17632
rect 10275 17660 10287 17663
rect 11882 17660 11888 17672
rect 10275 17632 11888 17660
rect 10275 17629 10287 17632
rect 10229 17623 10287 17629
rect 11882 17620 11888 17632
rect 11940 17620 11946 17672
rect 12066 17660 12072 17672
rect 12027 17632 12072 17660
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 13173 17663 13231 17669
rect 13173 17629 13185 17663
rect 13219 17660 13231 17663
rect 13354 17660 13360 17672
rect 13219 17632 13360 17660
rect 13219 17629 13231 17632
rect 13173 17623 13231 17629
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 13633 17663 13691 17669
rect 13633 17660 13645 17663
rect 13464 17632 13645 17660
rect 8665 17595 8723 17601
rect 8665 17561 8677 17595
rect 8711 17561 8723 17595
rect 8665 17555 8723 17561
rect 8680 17524 8708 17555
rect 8754 17552 8760 17604
rect 8812 17592 8818 17604
rect 10778 17592 10784 17604
rect 8812 17564 10784 17592
rect 8812 17552 8818 17564
rect 10778 17552 10784 17564
rect 10836 17552 10842 17604
rect 13464 17592 13492 17632
rect 13633 17629 13645 17632
rect 13679 17629 13691 17663
rect 13633 17623 13691 17629
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 15381 17663 15439 17669
rect 15381 17660 15393 17663
rect 14608 17632 15393 17660
rect 14608 17620 14614 17632
rect 15381 17629 15393 17632
rect 15427 17629 15439 17663
rect 15838 17660 15844 17672
rect 15799 17632 15844 17660
rect 15381 17623 15439 17629
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 18414 17660 18420 17672
rect 18375 17632 18420 17660
rect 18414 17620 18420 17632
rect 18472 17620 18478 17672
rect 19153 17663 19211 17669
rect 19153 17629 19165 17663
rect 19199 17660 19211 17663
rect 19334 17660 19340 17672
rect 19199 17632 19340 17660
rect 19199 17629 19211 17632
rect 19153 17623 19211 17629
rect 19334 17620 19340 17632
rect 19392 17620 19398 17672
rect 19981 17663 20039 17669
rect 19981 17629 19993 17663
rect 20027 17660 20039 17663
rect 21174 17660 21180 17672
rect 20027 17632 21180 17660
rect 20027 17629 20039 17632
rect 19981 17623 20039 17629
rect 21174 17620 21180 17632
rect 21232 17620 21238 17672
rect 21450 17660 21456 17672
rect 21411 17632 21456 17660
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 22370 17620 22376 17672
rect 22428 17660 22434 17672
rect 22925 17663 22983 17669
rect 22925 17660 22937 17663
rect 22428 17632 22937 17660
rect 22428 17620 22434 17632
rect 22925 17629 22937 17632
rect 22971 17629 22983 17663
rect 22925 17623 22983 17629
rect 10888 17564 13492 17592
rect 9858 17524 9864 17536
rect 8680 17496 9864 17524
rect 9858 17484 9864 17496
rect 9916 17524 9922 17536
rect 10888 17524 10916 17564
rect 15930 17552 15936 17604
rect 15988 17592 15994 17604
rect 16393 17595 16451 17601
rect 16393 17592 16405 17595
rect 15988 17564 16405 17592
rect 15988 17552 15994 17564
rect 16393 17561 16405 17564
rect 16439 17592 16451 17595
rect 22738 17592 22744 17604
rect 16439 17564 22744 17592
rect 16439 17561 16451 17564
rect 16393 17555 16451 17561
rect 22738 17552 22744 17564
rect 22796 17552 22802 17604
rect 9916 17496 10916 17524
rect 12805 17527 12863 17533
rect 9916 17484 9922 17496
rect 12805 17493 12817 17527
rect 12851 17524 12863 17527
rect 12894 17524 12900 17536
rect 12851 17496 12900 17524
rect 12851 17493 12863 17496
rect 12805 17487 12863 17493
rect 12894 17484 12900 17496
rect 12952 17484 12958 17536
rect 14274 17484 14280 17536
rect 14332 17524 14338 17536
rect 14737 17527 14795 17533
rect 14737 17524 14749 17527
rect 14332 17496 14749 17524
rect 14332 17484 14338 17496
rect 14737 17493 14749 17496
rect 14783 17524 14795 17527
rect 15562 17524 15568 17536
rect 14783 17496 15568 17524
rect 14783 17493 14795 17496
rect 14737 17487 14795 17493
rect 15562 17484 15568 17496
rect 15620 17484 15626 17536
rect 17586 17484 17592 17536
rect 17644 17524 17650 17536
rect 22462 17524 22468 17536
rect 17644 17496 22468 17524
rect 17644 17484 17650 17496
rect 22462 17484 22468 17496
rect 22520 17484 22526 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 7466 17320 7472 17332
rect 7427 17292 7472 17320
rect 7466 17280 7472 17292
rect 7524 17280 7530 17332
rect 7699 17323 7757 17329
rect 7699 17289 7711 17323
rect 7745 17320 7757 17323
rect 8110 17320 8116 17332
rect 7745 17292 8116 17320
rect 7745 17289 7757 17292
rect 7699 17283 7757 17289
rect 8110 17280 8116 17292
rect 8168 17280 8174 17332
rect 9490 17280 9496 17332
rect 9548 17320 9554 17332
rect 9585 17323 9643 17329
rect 9585 17320 9597 17323
rect 9548 17292 9597 17320
rect 9548 17280 9554 17292
rect 9585 17289 9597 17292
rect 9631 17289 9643 17323
rect 11790 17320 11796 17332
rect 11751 17292 11796 17320
rect 9585 17283 9643 17289
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 15378 17320 15384 17332
rect 15339 17292 15384 17320
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 15562 17280 15568 17332
rect 15620 17320 15626 17332
rect 18187 17323 18245 17329
rect 18187 17320 18199 17323
rect 15620 17292 18199 17320
rect 15620 17280 15626 17292
rect 18187 17289 18199 17292
rect 18233 17289 18245 17323
rect 18187 17283 18245 17289
rect 22646 17280 22652 17332
rect 22704 17320 22710 17332
rect 24121 17323 24179 17329
rect 24121 17320 24133 17323
rect 22704 17292 24133 17320
rect 22704 17280 22710 17292
rect 24121 17289 24133 17292
rect 24167 17289 24179 17323
rect 24121 17283 24179 17289
rect 15013 17255 15071 17261
rect 15013 17221 15025 17255
rect 15059 17252 15071 17255
rect 15470 17252 15476 17264
rect 15059 17224 15476 17252
rect 15059 17221 15071 17224
rect 15013 17215 15071 17221
rect 15470 17212 15476 17224
rect 15528 17252 15534 17264
rect 16853 17255 16911 17261
rect 16853 17252 16865 17255
rect 15528 17224 16865 17252
rect 15528 17212 15534 17224
rect 16853 17221 16865 17224
rect 16899 17221 16911 17255
rect 16853 17215 16911 17221
rect 20898 17212 20904 17264
rect 20956 17252 20962 17264
rect 22189 17255 22247 17261
rect 22189 17252 22201 17255
rect 20956 17224 22201 17252
rect 20956 17212 20962 17224
rect 22189 17221 22201 17224
rect 22235 17252 22247 17255
rect 23106 17252 23112 17264
rect 22235 17224 23112 17252
rect 22235 17221 22247 17224
rect 22189 17215 22247 17221
rect 23106 17212 23112 17224
rect 23164 17212 23170 17264
rect 7190 17144 7196 17196
rect 7248 17184 7254 17196
rect 10045 17187 10103 17193
rect 10045 17184 10057 17187
rect 7248 17156 10057 17184
rect 7248 17144 7254 17156
rect 10045 17153 10057 17156
rect 10091 17184 10103 17187
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10091 17156 10609 17184
rect 10091 17153 10103 17156
rect 10045 17147 10103 17153
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 14090 17184 14096 17196
rect 14051 17156 14096 17184
rect 10597 17147 10655 17153
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 15562 17144 15568 17196
rect 15620 17184 15626 17196
rect 16209 17187 16267 17193
rect 16209 17184 16221 17187
rect 15620 17156 16221 17184
rect 15620 17144 15626 17156
rect 16209 17153 16221 17156
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 17402 17144 17408 17196
rect 17460 17184 17466 17196
rect 17681 17187 17739 17193
rect 17681 17184 17693 17187
rect 17460 17156 17693 17184
rect 17460 17144 17466 17156
rect 17681 17153 17693 17156
rect 17727 17184 17739 17187
rect 17954 17184 17960 17196
rect 17727 17156 17960 17184
rect 17727 17153 17739 17156
rect 17681 17147 17739 17153
rect 17954 17144 17960 17156
rect 18012 17144 18018 17196
rect 20625 17187 20683 17193
rect 20625 17153 20637 17187
rect 20671 17184 20683 17187
rect 20809 17187 20867 17193
rect 20809 17184 20821 17187
rect 20671 17156 20821 17184
rect 20671 17153 20683 17156
rect 20625 17147 20683 17153
rect 20809 17153 20821 17156
rect 20855 17184 20867 17187
rect 23661 17187 23719 17193
rect 23661 17184 23673 17187
rect 20855 17156 23673 17184
rect 20855 17153 20867 17156
rect 20809 17147 20867 17153
rect 23661 17153 23673 17156
rect 23707 17153 23719 17187
rect 23661 17147 23719 17153
rect 6086 17076 6092 17128
rect 6144 17116 6150 17128
rect 7650 17125 7656 17128
rect 7628 17119 7656 17125
rect 7628 17116 7640 17119
rect 6144 17088 7640 17116
rect 6144 17076 6150 17088
rect 7628 17085 7640 17088
rect 7708 17116 7714 17128
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7708 17088 8033 17116
rect 7628 17079 7656 17085
rect 7650 17076 7656 17079
rect 7708 17076 7714 17088
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8662 17116 8668 17128
rect 8623 17088 8668 17116
rect 8021 17079 8079 17085
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 12618 17116 12624 17128
rect 12579 17088 12624 17116
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 12894 17116 12900 17128
rect 12855 17088 12900 17116
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 16758 17076 16764 17128
rect 16816 17116 16822 17128
rect 18116 17119 18174 17125
rect 18116 17116 18128 17119
rect 16816 17088 18128 17116
rect 16816 17076 16822 17088
rect 18116 17085 18128 17088
rect 18162 17116 18174 17119
rect 22348 17119 22406 17125
rect 18162 17088 18644 17116
rect 18162 17085 18174 17088
rect 18116 17079 18174 17085
rect 8573 17051 8631 17057
rect 8573 17017 8585 17051
rect 8619 17048 8631 17051
rect 8986 17051 9044 17057
rect 8986 17048 8998 17051
rect 8619 17020 8998 17048
rect 8619 17017 8631 17020
rect 8573 17011 8631 17017
rect 8986 17017 8998 17020
rect 9032 17048 9044 17051
rect 10042 17048 10048 17060
rect 9032 17020 10048 17048
rect 9032 17017 9044 17020
rect 8986 17011 9044 17017
rect 10042 17008 10048 17020
rect 10100 17048 10106 17060
rect 10413 17051 10471 17057
rect 10413 17048 10425 17051
rect 10100 17020 10425 17048
rect 10100 17008 10106 17020
rect 10413 17017 10425 17020
rect 10459 17048 10471 17051
rect 10918 17051 10976 17057
rect 10918 17048 10930 17051
rect 10459 17020 10930 17048
rect 10459 17017 10471 17020
rect 10413 17011 10471 17017
rect 10918 17017 10930 17020
rect 10964 17017 10976 17051
rect 10918 17011 10976 17017
rect 12253 17051 12311 17057
rect 12253 17017 12265 17051
rect 12299 17048 12311 17051
rect 12912 17048 12940 17076
rect 13170 17048 13176 17060
rect 12299 17020 12940 17048
rect 13131 17020 13176 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 13170 17008 13176 17020
rect 13228 17008 13234 17060
rect 14414 17051 14472 17057
rect 14414 17017 14426 17051
rect 14460 17017 14472 17051
rect 14414 17011 14472 17017
rect 15749 17051 15807 17057
rect 15749 17017 15761 17051
rect 15795 17048 15807 17051
rect 15930 17048 15936 17060
rect 15795 17020 15936 17048
rect 15795 17017 15807 17020
rect 15749 17011 15807 17017
rect 11517 16983 11575 16989
rect 11517 16949 11529 16983
rect 11563 16980 11575 16983
rect 11698 16980 11704 16992
rect 11563 16952 11704 16980
rect 11563 16949 11575 16952
rect 11517 16943 11575 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 13446 16980 13452 16992
rect 13407 16952 13452 16980
rect 13446 16940 13452 16952
rect 13504 16940 13510 16992
rect 13906 16980 13912 16992
rect 13867 16952 13912 16980
rect 13906 16940 13912 16952
rect 13964 16980 13970 16992
rect 14429 16980 14457 17011
rect 15930 17008 15936 17020
rect 15988 17008 15994 17060
rect 16025 17051 16083 17057
rect 16025 17017 16037 17051
rect 16071 17017 16083 17051
rect 16025 17011 16083 17017
rect 13964 16952 14457 16980
rect 13964 16940 13970 16952
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 16040 16980 16068 17011
rect 16206 16980 16212 16992
rect 15436 16952 16212 16980
rect 15436 16940 15442 16952
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 17405 16983 17463 16989
rect 17405 16949 17417 16983
rect 17451 16980 17463 16983
rect 17586 16980 17592 16992
rect 17451 16952 17592 16980
rect 17451 16949 17463 16952
rect 17405 16943 17463 16949
rect 17586 16940 17592 16952
rect 17644 16940 17650 16992
rect 18616 16989 18644 17088
rect 22348 17085 22360 17119
rect 22394 17116 22406 17119
rect 22462 17116 22468 17128
rect 22394 17088 22468 17116
rect 22394 17085 22406 17088
rect 22348 17079 22406 17085
rect 22462 17076 22468 17088
rect 22520 17116 22526 17128
rect 22741 17119 22799 17125
rect 22741 17116 22753 17119
rect 22520 17088 22753 17116
rect 22520 17076 22526 17088
rect 22741 17085 22753 17088
rect 22787 17116 22799 17119
rect 23842 17116 23848 17128
rect 22787 17088 23848 17116
rect 22787 17085 22799 17088
rect 22741 17079 22799 17085
rect 23842 17076 23848 17088
rect 23900 17076 23906 17128
rect 18782 17008 18788 17060
rect 18840 17048 18846 17060
rect 19245 17051 19303 17057
rect 19245 17048 19257 17051
rect 18840 17020 19257 17048
rect 18840 17008 18846 17020
rect 19245 17017 19257 17020
rect 19291 17017 19303 17051
rect 19245 17011 19303 17017
rect 19337 17051 19395 17057
rect 19337 17017 19349 17051
rect 19383 17048 19395 17051
rect 19426 17048 19432 17060
rect 19383 17020 19432 17048
rect 19383 17017 19395 17020
rect 19337 17011 19395 17017
rect 18601 16983 18659 16989
rect 18601 16949 18613 16983
rect 18647 16980 18659 16983
rect 18690 16980 18696 16992
rect 18647 16952 18696 16980
rect 18647 16949 18659 16952
rect 18601 16943 18659 16949
rect 18690 16940 18696 16952
rect 18748 16940 18754 16992
rect 18966 16980 18972 16992
rect 18927 16952 18972 16980
rect 18966 16940 18972 16952
rect 19024 16980 19030 16992
rect 19352 16980 19380 17011
rect 19426 17008 19432 17020
rect 19484 17008 19490 17060
rect 19889 17051 19947 17057
rect 19889 17017 19901 17051
rect 19935 17048 19947 17051
rect 20622 17048 20628 17060
rect 19935 17020 20628 17048
rect 19935 17017 19947 17020
rect 19889 17011 19947 17017
rect 20622 17008 20628 17020
rect 20680 17008 20686 17060
rect 20898 17048 20904 17060
rect 20859 17020 20904 17048
rect 20898 17008 20904 17020
rect 20956 17008 20962 17060
rect 21450 17048 21456 17060
rect 21411 17020 21456 17048
rect 21450 17008 21456 17020
rect 21508 17008 21514 17060
rect 20165 16983 20223 16989
rect 20165 16980 20177 16983
rect 19024 16952 20177 16980
rect 19024 16940 19030 16952
rect 20165 16949 20177 16952
rect 20211 16949 20223 16983
rect 20165 16943 20223 16949
rect 21542 16940 21548 16992
rect 21600 16980 21606 16992
rect 21729 16983 21787 16989
rect 21729 16980 21741 16983
rect 21600 16952 21741 16980
rect 21600 16940 21606 16952
rect 21729 16949 21741 16952
rect 21775 16949 21787 16983
rect 21729 16943 21787 16949
rect 22419 16983 22477 16989
rect 22419 16949 22431 16983
rect 22465 16980 22477 16983
rect 22554 16980 22560 16992
rect 22465 16952 22560 16980
rect 22465 16949 22477 16952
rect 22419 16943 22477 16949
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 24210 16940 24216 16992
rect 24268 16980 24274 16992
rect 24581 16983 24639 16989
rect 24581 16980 24593 16983
rect 24268 16952 24593 16980
rect 24268 16940 24274 16952
rect 24581 16949 24593 16952
rect 24627 16949 24639 16983
rect 24581 16943 24639 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 7929 16779 7987 16785
rect 7929 16745 7941 16779
rect 7975 16776 7987 16779
rect 8110 16776 8116 16788
rect 7975 16748 8116 16776
rect 7975 16745 7987 16748
rect 7929 16739 7987 16745
rect 8110 16736 8116 16748
rect 8168 16736 8174 16788
rect 10042 16776 10048 16788
rect 10003 16748 10048 16776
rect 10042 16736 10048 16748
rect 10100 16736 10106 16788
rect 10597 16779 10655 16785
rect 10597 16745 10609 16779
rect 10643 16776 10655 16779
rect 10686 16776 10692 16788
rect 10643 16748 10692 16776
rect 10643 16745 10655 16748
rect 10597 16739 10655 16745
rect 10686 16736 10692 16748
rect 10744 16776 10750 16788
rect 10873 16779 10931 16785
rect 10873 16776 10885 16779
rect 10744 16748 10885 16776
rect 10744 16736 10750 16748
rect 10873 16745 10885 16748
rect 10919 16745 10931 16779
rect 10873 16739 10931 16745
rect 14550 16736 14556 16788
rect 14608 16776 14614 16788
rect 15013 16779 15071 16785
rect 15013 16776 15025 16779
rect 14608 16748 15025 16776
rect 14608 16736 14614 16748
rect 15013 16745 15025 16748
rect 15059 16745 15071 16779
rect 16206 16776 16212 16788
rect 16167 16748 16212 16776
rect 15013 16739 15071 16745
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 19242 16736 19248 16788
rect 19300 16776 19306 16788
rect 19337 16779 19395 16785
rect 19337 16776 19349 16779
rect 19300 16748 19349 16776
rect 19300 16736 19306 16748
rect 19337 16745 19349 16748
rect 19383 16745 19395 16779
rect 19337 16739 19395 16745
rect 19889 16779 19947 16785
rect 19889 16745 19901 16779
rect 19935 16745 19947 16779
rect 19889 16739 19947 16745
rect 20717 16779 20775 16785
rect 20717 16745 20729 16779
rect 20763 16776 20775 16779
rect 20990 16776 20996 16788
rect 20763 16748 20996 16776
rect 20763 16745 20775 16748
rect 20717 16739 20775 16745
rect 7190 16708 7196 16720
rect 7151 16680 7196 16708
rect 7190 16668 7196 16680
rect 7248 16668 7254 16720
rect 8662 16668 8668 16720
rect 8720 16708 8726 16720
rect 8757 16711 8815 16717
rect 8757 16708 8769 16711
rect 8720 16680 8769 16708
rect 8720 16668 8726 16680
rect 8757 16677 8769 16680
rect 8803 16708 8815 16711
rect 9033 16711 9091 16717
rect 9033 16708 9045 16711
rect 8803 16680 9045 16708
rect 8803 16677 8815 16680
rect 8757 16671 8815 16677
rect 9033 16677 9045 16680
rect 9079 16677 9091 16711
rect 11606 16708 11612 16720
rect 11567 16680 11612 16708
rect 9033 16671 9091 16677
rect 11606 16668 11612 16680
rect 11664 16668 11670 16720
rect 11698 16668 11704 16720
rect 11756 16708 11762 16720
rect 13265 16711 13323 16717
rect 13265 16708 13277 16711
rect 11756 16680 13277 16708
rect 11756 16668 11762 16680
rect 13265 16677 13277 16680
rect 13311 16708 13323 16711
rect 13446 16708 13452 16720
rect 13311 16680 13452 16708
rect 13311 16677 13323 16680
rect 13265 16671 13323 16677
rect 13446 16668 13452 16680
rect 13504 16668 13510 16720
rect 13538 16668 13544 16720
rect 13596 16708 13602 16720
rect 13725 16711 13783 16717
rect 13725 16708 13737 16711
rect 13596 16680 13737 16708
rect 13596 16668 13602 16680
rect 13725 16677 13737 16680
rect 13771 16677 13783 16711
rect 13725 16671 13783 16677
rect 13814 16668 13820 16720
rect 13872 16708 13878 16720
rect 14369 16711 14427 16717
rect 13872 16680 13917 16708
rect 13872 16668 13878 16680
rect 14369 16677 14381 16711
rect 14415 16708 14427 16711
rect 14568 16708 14596 16736
rect 14415 16680 14596 16708
rect 14415 16677 14427 16680
rect 14369 16671 14427 16677
rect 15286 16668 15292 16720
rect 15344 16708 15350 16720
rect 15610 16711 15668 16717
rect 15610 16708 15622 16711
rect 15344 16680 15622 16708
rect 15344 16668 15350 16680
rect 15610 16677 15622 16680
rect 15656 16677 15668 16711
rect 19904 16708 19932 16739
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 21542 16736 21548 16788
rect 21600 16776 21606 16788
rect 21600 16748 22692 16776
rect 21600 16736 21606 16748
rect 20806 16708 20812 16720
rect 19904 16680 20812 16708
rect 15610 16671 15668 16677
rect 20806 16668 20812 16680
rect 20864 16708 20870 16720
rect 21085 16711 21143 16717
rect 21085 16708 21097 16711
rect 20864 16680 21097 16708
rect 20864 16668 20870 16680
rect 21085 16677 21097 16680
rect 21131 16677 21143 16711
rect 21085 16671 21143 16677
rect 21174 16668 21180 16720
rect 21232 16708 21238 16720
rect 21637 16711 21695 16717
rect 21637 16708 21649 16711
rect 21232 16680 21649 16708
rect 21232 16668 21238 16680
rect 21637 16677 21649 16680
rect 21683 16677 21695 16711
rect 22554 16708 22560 16720
rect 22515 16680 22560 16708
rect 21637 16671 21695 16677
rect 22554 16668 22560 16680
rect 22612 16668 22618 16720
rect 22664 16717 22692 16748
rect 22649 16711 22707 16717
rect 22649 16677 22661 16711
rect 22695 16708 22707 16711
rect 23198 16708 23204 16720
rect 22695 16680 23204 16708
rect 22695 16677 22707 16680
rect 22649 16671 22707 16677
rect 23198 16668 23204 16680
rect 23256 16668 23262 16720
rect 6730 16640 6736 16652
rect 6691 16612 6736 16640
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 7009 16643 7067 16649
rect 7009 16609 7021 16643
rect 7055 16609 7067 16643
rect 8110 16640 8116 16652
rect 8071 16612 8116 16640
rect 7009 16603 7067 16609
rect 7024 16572 7052 16603
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 8386 16600 8392 16652
rect 8444 16640 8450 16652
rect 8481 16643 8539 16649
rect 8481 16640 8493 16643
rect 8444 16612 8493 16640
rect 8444 16600 8450 16612
rect 8481 16609 8493 16612
rect 8527 16609 8539 16643
rect 17034 16640 17040 16652
rect 16995 16612 17040 16640
rect 8481 16603 8539 16609
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 17402 16600 17408 16652
rect 17460 16640 17466 16652
rect 17497 16643 17555 16649
rect 17497 16640 17509 16643
rect 17460 16612 17509 16640
rect 17460 16600 17466 16612
rect 17497 16609 17509 16612
rect 17543 16609 17555 16643
rect 17497 16603 17555 16609
rect 18414 16600 18420 16652
rect 18472 16640 18478 16652
rect 18969 16643 19027 16649
rect 18969 16640 18981 16643
rect 18472 16612 18981 16640
rect 18472 16600 18478 16612
rect 18969 16609 18981 16612
rect 19015 16640 19027 16643
rect 19610 16640 19616 16652
rect 19015 16612 19616 16640
rect 19015 16609 19027 16612
rect 18969 16603 19027 16609
rect 19610 16600 19616 16612
rect 19668 16600 19674 16652
rect 8404 16572 8432 16600
rect 9674 16572 9680 16584
rect 7024 16544 8432 16572
rect 9635 16544 9680 16572
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 11882 16572 11888 16584
rect 11843 16544 11888 16572
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 14826 16532 14832 16584
rect 14884 16572 14890 16584
rect 15289 16575 15347 16581
rect 15289 16572 15301 16575
rect 14884 16544 15301 16572
rect 14884 16532 14890 16544
rect 15289 16541 15301 16544
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 17773 16575 17831 16581
rect 17773 16541 17785 16575
rect 17819 16572 17831 16575
rect 18046 16572 18052 16584
rect 17819 16544 18052 16572
rect 17819 16541 17831 16544
rect 17773 16535 17831 16541
rect 18046 16532 18052 16544
rect 18104 16532 18110 16584
rect 20993 16575 21051 16581
rect 20993 16541 21005 16575
rect 21039 16572 21051 16575
rect 22186 16572 22192 16584
rect 21039 16544 22192 16572
rect 21039 16541 21051 16544
rect 20993 16535 21051 16541
rect 22186 16532 22192 16544
rect 22244 16532 22250 16584
rect 22370 16532 22376 16584
rect 22428 16572 22434 16584
rect 22833 16575 22891 16581
rect 22833 16572 22845 16575
rect 22428 16544 22845 16572
rect 22428 16532 22434 16544
rect 22833 16541 22845 16544
rect 22879 16541 22891 16575
rect 22833 16535 22891 16541
rect 12618 16436 12624 16448
rect 12579 16408 12624 16436
rect 12618 16396 12624 16408
rect 12676 16396 12682 16448
rect 18782 16436 18788 16448
rect 18743 16408 18788 16436
rect 18782 16396 18788 16408
rect 18840 16396 18846 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 8110 16232 8116 16244
rect 8071 16204 8116 16232
rect 8110 16192 8116 16204
rect 8168 16192 8174 16244
rect 9401 16235 9459 16241
rect 9401 16201 9413 16235
rect 9447 16232 9459 16235
rect 9674 16232 9680 16244
rect 9447 16204 9680 16232
rect 9447 16201 9459 16204
rect 9401 16195 9459 16201
rect 6549 16099 6607 16105
rect 6549 16065 6561 16099
rect 6595 16096 6607 16099
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 6595 16068 7757 16096
rect 6595 16065 6607 16068
rect 6549 16059 6607 16065
rect 7745 16065 7757 16068
rect 7791 16096 7803 16099
rect 9033 16099 9091 16105
rect 7791 16068 8432 16096
rect 7791 16065 7803 16068
rect 7745 16059 7803 16065
rect 8404 16040 8432 16068
rect 9033 16065 9045 16099
rect 9079 16096 9091 16099
rect 9416 16096 9444 16195
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 9766 16192 9772 16244
rect 9824 16232 9830 16244
rect 10042 16232 10048 16244
rect 9824 16204 10048 16232
rect 9824 16192 9830 16204
rect 10042 16192 10048 16204
rect 10100 16232 10106 16244
rect 10100 16204 11146 16232
rect 10100 16192 10106 16204
rect 10505 16167 10563 16173
rect 10505 16133 10517 16167
rect 10551 16164 10563 16167
rect 10778 16164 10784 16176
rect 10551 16136 10784 16164
rect 10551 16133 10563 16136
rect 10505 16127 10563 16133
rect 10778 16124 10784 16136
rect 10836 16124 10842 16176
rect 11118 16164 11146 16204
rect 11606 16192 11612 16244
rect 11664 16232 11670 16244
rect 11885 16235 11943 16241
rect 11885 16232 11897 16235
rect 11664 16204 11897 16232
rect 11664 16192 11670 16204
rect 11885 16201 11897 16204
rect 11931 16201 11943 16235
rect 11885 16195 11943 16201
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 14277 16235 14335 16241
rect 14277 16232 14289 16235
rect 13872 16204 14289 16232
rect 13872 16192 13878 16204
rect 14277 16201 14289 16204
rect 14323 16201 14335 16235
rect 14277 16195 14335 16201
rect 14826 16192 14832 16244
rect 14884 16232 14890 16244
rect 14921 16235 14979 16241
rect 14921 16232 14933 16235
rect 14884 16204 14933 16232
rect 14884 16192 14890 16204
rect 14921 16201 14933 16204
rect 14967 16201 14979 16235
rect 14921 16195 14979 16201
rect 16022 16192 16028 16244
rect 16080 16232 16086 16244
rect 18966 16232 18972 16244
rect 16080 16204 18413 16232
rect 18927 16204 18972 16232
rect 16080 16192 16086 16204
rect 12897 16167 12955 16173
rect 12897 16164 12909 16167
rect 11118 16136 12909 16164
rect 12897 16133 12909 16136
rect 12943 16133 12955 16167
rect 16114 16164 16120 16176
rect 12897 16127 12955 16133
rect 15580 16136 16120 16164
rect 9079 16068 9444 16096
rect 9079 16065 9091 16068
rect 9033 16059 9091 16065
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 11609 16099 11667 16105
rect 9640 16056 9674 16096
rect 11609 16065 11621 16099
rect 11655 16096 11667 16099
rect 11698 16096 11704 16108
rect 11655 16068 11704 16096
rect 11655 16065 11667 16068
rect 11609 16059 11667 16065
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 8294 16028 8300 16040
rect 8255 16000 8300 16028
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 8757 16031 8815 16037
rect 8757 16028 8769 16031
rect 8444 16000 8769 16028
rect 8444 15988 8450 16000
rect 8757 15997 8769 16000
rect 8803 15997 8815 16031
rect 8757 15991 8815 15997
rect 6730 15920 6736 15972
rect 6788 15960 6794 15972
rect 7101 15963 7159 15969
rect 7101 15960 7113 15963
rect 6788 15932 7113 15960
rect 6788 15920 6794 15932
rect 7101 15929 7113 15932
rect 7147 15960 7159 15963
rect 8938 15960 8944 15972
rect 7147 15932 8944 15960
rect 7147 15929 7159 15932
rect 7101 15923 7159 15929
rect 8938 15920 8944 15932
rect 8996 15920 9002 15972
rect 9646 15960 9674 16056
rect 9950 15960 9956 15972
rect 9646 15932 9956 15960
rect 9950 15920 9956 15932
rect 10008 15920 10014 15972
rect 10045 15963 10103 15969
rect 10045 15929 10057 15963
rect 10091 15929 10103 15963
rect 12912 15960 12940 16127
rect 13081 16099 13139 16105
rect 13081 16065 13093 16099
rect 13127 16096 13139 16099
rect 13170 16096 13176 16108
rect 13127 16068 13176 16096
rect 13127 16065 13139 16068
rect 13081 16059 13139 16065
rect 13170 16056 13176 16068
rect 13228 16056 13234 16108
rect 15580 16105 15608 16136
rect 16114 16124 16120 16136
rect 16172 16124 16178 16176
rect 15565 16099 15623 16105
rect 15565 16065 15577 16099
rect 15611 16065 15623 16099
rect 15838 16096 15844 16108
rect 15799 16068 15844 16096
rect 15565 16059 15623 16065
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 18046 16096 18052 16108
rect 18007 16068 18052 16096
rect 18046 16056 18052 16068
rect 18104 16056 18110 16108
rect 18385 16096 18413 16204
rect 18966 16192 18972 16204
rect 19024 16192 19030 16244
rect 19334 16192 19340 16244
rect 19392 16232 19398 16244
rect 19935 16235 19993 16241
rect 19935 16232 19947 16235
rect 19392 16204 19947 16232
rect 19392 16192 19398 16204
rect 19935 16201 19947 16204
rect 19981 16201 19993 16235
rect 19935 16195 19993 16201
rect 20717 16235 20775 16241
rect 20717 16201 20729 16235
rect 20763 16232 20775 16235
rect 20806 16232 20812 16244
rect 20763 16204 20812 16232
rect 20763 16201 20775 16204
rect 20717 16195 20775 16201
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 22186 16232 22192 16244
rect 22147 16204 22192 16232
rect 22186 16192 22192 16204
rect 22244 16232 22250 16244
rect 22511 16235 22569 16241
rect 22511 16232 22523 16235
rect 22244 16204 22523 16232
rect 22244 16192 22250 16204
rect 22511 16201 22523 16204
rect 22557 16201 22569 16235
rect 22922 16232 22928 16244
rect 22883 16204 22928 16232
rect 22511 16195 22569 16201
rect 22922 16192 22928 16204
rect 22980 16192 22986 16244
rect 23198 16232 23204 16244
rect 23159 16204 23204 16232
rect 23198 16192 23204 16204
rect 23256 16192 23262 16244
rect 19610 16164 19616 16176
rect 19571 16136 19616 16164
rect 19610 16124 19616 16136
rect 19668 16124 19674 16176
rect 18598 16096 18604 16108
rect 18385 16068 18604 16096
rect 18598 16056 18604 16068
rect 18656 16096 18662 16108
rect 20901 16099 20959 16105
rect 18656 16068 19104 16096
rect 18656 16056 18662 16068
rect 17218 15988 17224 16040
rect 17276 16028 17282 16040
rect 18966 16028 18972 16040
rect 17276 16000 18972 16028
rect 17276 15988 17282 16000
rect 18966 15988 18972 16000
rect 19024 15988 19030 16040
rect 19076 16028 19104 16068
rect 20901 16065 20913 16099
rect 20947 16096 20959 16099
rect 21174 16096 21180 16108
rect 20947 16068 21180 16096
rect 20947 16065 20959 16068
rect 20901 16059 20959 16065
rect 21174 16056 21180 16068
rect 21232 16056 21238 16108
rect 19832 16031 19890 16037
rect 19832 16028 19844 16031
rect 19076 16000 19844 16028
rect 19832 15997 19844 16000
rect 19878 16028 19890 16031
rect 20257 16031 20315 16037
rect 20257 16028 20269 16031
rect 19878 16000 20269 16028
rect 19878 15997 19890 16000
rect 19832 15991 19890 15997
rect 20257 15997 20269 16000
rect 20303 15997 20315 16031
rect 20257 15991 20315 15997
rect 22440 16031 22498 16037
rect 22440 15997 22452 16031
rect 22486 16028 22498 16031
rect 22922 16028 22928 16040
rect 22486 16000 22928 16028
rect 22486 15997 22498 16000
rect 22440 15991 22498 15997
rect 22922 15988 22928 16000
rect 22980 15988 22986 16040
rect 13446 15969 13452 15972
rect 13402 15963 13452 15969
rect 13402 15960 13414 15963
rect 12912 15932 13414 15960
rect 10045 15923 10103 15929
rect 13402 15929 13414 15932
rect 13448 15929 13452 15963
rect 13402 15923 13452 15929
rect 10060 15892 10088 15923
rect 13446 15920 13452 15923
rect 13504 15960 13510 15972
rect 13906 15960 13912 15972
rect 13504 15932 13912 15960
rect 13504 15920 13510 15932
rect 13906 15920 13912 15932
rect 13964 15960 13970 15972
rect 15286 15960 15292 15972
rect 13964 15932 15292 15960
rect 13964 15920 13970 15932
rect 15286 15920 15292 15932
rect 15344 15920 15350 15972
rect 15657 15963 15715 15969
rect 15657 15929 15669 15963
rect 15703 15929 15715 15963
rect 15657 15923 15715 15929
rect 10134 15892 10140 15904
rect 10047 15864 10140 15892
rect 10134 15852 10140 15864
rect 10192 15892 10198 15904
rect 10873 15895 10931 15901
rect 10873 15892 10885 15895
rect 10192 15864 10885 15892
rect 10192 15852 10198 15864
rect 10873 15861 10885 15864
rect 10919 15861 10931 15895
rect 10873 15855 10931 15861
rect 13722 15852 13728 15904
rect 13780 15892 13786 15904
rect 14001 15895 14059 15901
rect 14001 15892 14013 15895
rect 13780 15864 14013 15892
rect 13780 15852 13786 15864
rect 14001 15861 14013 15864
rect 14047 15861 14059 15895
rect 15672 15892 15700 15923
rect 16022 15920 16028 15972
rect 16080 15960 16086 15972
rect 17034 15960 17040 15972
rect 16080 15932 17040 15960
rect 16080 15920 16086 15932
rect 17034 15920 17040 15932
rect 17092 15920 17098 15972
rect 18370 15963 18428 15969
rect 18370 15960 18382 15963
rect 17788 15932 18382 15960
rect 17788 15904 17816 15932
rect 18370 15929 18382 15932
rect 18416 15929 18428 15963
rect 18370 15923 18428 15929
rect 20990 15920 20996 15972
rect 21048 15960 21054 15972
rect 21545 15963 21603 15969
rect 21048 15932 21093 15960
rect 21048 15920 21054 15932
rect 21545 15929 21557 15963
rect 21591 15960 21603 15963
rect 21726 15960 21732 15972
rect 21591 15932 21732 15960
rect 21591 15929 21603 15932
rect 21545 15923 21603 15929
rect 21726 15920 21732 15932
rect 21784 15920 21790 15972
rect 16114 15892 16120 15904
rect 15672 15864 16120 15892
rect 14001 15855 14059 15861
rect 16114 15852 16120 15864
rect 16172 15892 16178 15904
rect 16485 15895 16543 15901
rect 16485 15892 16497 15895
rect 16172 15864 16497 15892
rect 16172 15852 16178 15864
rect 16485 15861 16497 15864
rect 16531 15861 16543 15895
rect 17402 15892 17408 15904
rect 17363 15864 17408 15892
rect 16485 15855 16543 15861
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 17770 15892 17776 15904
rect 17731 15864 17776 15892
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 19334 15852 19340 15904
rect 19392 15892 19398 15904
rect 21008 15892 21036 15920
rect 21821 15895 21879 15901
rect 21821 15892 21833 15895
rect 19392 15864 19437 15892
rect 21008 15864 21833 15892
rect 19392 15852 19398 15864
rect 21821 15861 21833 15864
rect 21867 15861 21879 15895
rect 21821 15855 21879 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1578 15688 1584 15700
rect 1539 15660 1584 15688
rect 1578 15648 1584 15660
rect 1636 15648 1642 15700
rect 13170 15688 13176 15700
rect 13131 15660 13176 15688
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 13538 15688 13544 15700
rect 13499 15660 13544 15688
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 15930 15648 15936 15700
rect 15988 15688 15994 15700
rect 16853 15691 16911 15697
rect 16853 15688 16865 15691
rect 15988 15660 16865 15688
rect 15988 15648 15994 15660
rect 16853 15657 16865 15660
rect 16899 15657 16911 15691
rect 16853 15651 16911 15657
rect 20717 15691 20775 15697
rect 20717 15657 20729 15691
rect 20763 15688 20775 15691
rect 21174 15688 21180 15700
rect 20763 15660 21180 15688
rect 20763 15657 20775 15660
rect 20717 15651 20775 15657
rect 21174 15648 21180 15660
rect 21232 15648 21238 15700
rect 22554 15688 22560 15700
rect 22515 15660 22560 15688
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 9861 15623 9919 15629
rect 9861 15589 9873 15623
rect 9907 15620 9919 15623
rect 10042 15620 10048 15632
rect 9907 15592 10048 15620
rect 9907 15589 9919 15592
rect 9861 15583 9919 15589
rect 10042 15580 10048 15592
rect 10100 15620 10106 15632
rect 10502 15620 10508 15632
rect 10100 15592 10508 15620
rect 10100 15580 10106 15592
rect 10502 15580 10508 15592
rect 10560 15580 10566 15632
rect 10962 15580 10968 15632
rect 11020 15620 11026 15632
rect 11517 15623 11575 15629
rect 11517 15620 11529 15623
rect 11020 15592 11529 15620
rect 11020 15580 11026 15592
rect 11517 15589 11529 15592
rect 11563 15589 11575 15623
rect 11517 15583 11575 15589
rect 13722 15580 13728 15632
rect 13780 15620 13786 15632
rect 13817 15623 13875 15629
rect 13817 15620 13829 15623
rect 13780 15592 13829 15620
rect 13780 15580 13786 15592
rect 13817 15589 13829 15592
rect 13863 15589 13875 15623
rect 15470 15620 15476 15632
rect 15431 15592 15476 15620
rect 13817 15583 13875 15589
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 16206 15580 16212 15632
rect 16264 15620 16270 15632
rect 16301 15623 16359 15629
rect 16301 15620 16313 15623
rect 16264 15592 16313 15620
rect 16264 15580 16270 15592
rect 16301 15589 16313 15592
rect 16347 15589 16359 15623
rect 16301 15583 16359 15589
rect 17770 15580 17776 15632
rect 17828 15620 17834 15632
rect 18278 15623 18336 15629
rect 18278 15620 18290 15623
rect 17828 15592 18290 15620
rect 17828 15580 17834 15592
rect 18278 15589 18290 15592
rect 18324 15589 18336 15623
rect 18278 15583 18336 15589
rect 20806 15580 20812 15632
rect 20864 15620 20870 15632
rect 21085 15623 21143 15629
rect 21085 15620 21097 15623
rect 20864 15592 21097 15620
rect 20864 15580 20870 15592
rect 21085 15589 21097 15592
rect 21131 15589 21143 15623
rect 21085 15583 21143 15589
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 10413 15555 10471 15561
rect 10413 15521 10425 15555
rect 10459 15552 10471 15555
rect 10778 15552 10784 15564
rect 10459 15524 10784 15552
rect 10459 15521 10471 15524
rect 10413 15515 10471 15521
rect 10778 15512 10784 15524
rect 10836 15512 10842 15564
rect 12066 15512 12072 15564
rect 12124 15552 12130 15564
rect 19772 15555 19830 15561
rect 12124 15524 12169 15552
rect 12124 15512 12130 15524
rect 19772 15521 19784 15555
rect 19818 15552 19830 15555
rect 20254 15552 20260 15564
rect 19818 15524 20260 15552
rect 19818 15521 19830 15524
rect 19772 15515 19830 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 9769 15487 9827 15493
rect 9769 15453 9781 15487
rect 9815 15484 9827 15487
rect 9858 15484 9864 15496
rect 9815 15456 9864 15484
rect 9815 15453 9827 15456
rect 9769 15447 9827 15453
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 11425 15487 11483 15493
rect 11425 15453 11437 15487
rect 11471 15484 11483 15487
rect 11698 15484 11704 15496
rect 11471 15456 11704 15484
rect 11471 15453 11483 15456
rect 11425 15447 11483 15453
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 12986 15444 12992 15496
rect 13044 15484 13050 15496
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 13044 15456 13737 15484
rect 13044 15444 13050 15456
rect 13725 15453 13737 15456
rect 13771 15453 13783 15487
rect 13725 15447 13783 15453
rect 14369 15487 14427 15493
rect 14369 15453 14381 15487
rect 14415 15484 14427 15487
rect 15381 15487 15439 15493
rect 15381 15484 15393 15487
rect 14415 15456 15393 15484
rect 14415 15453 14427 15456
rect 14369 15447 14427 15453
rect 15381 15453 15393 15456
rect 15427 15484 15439 15487
rect 15562 15484 15568 15496
rect 15427 15456 15568 15484
rect 15427 15453 15439 15456
rect 15381 15447 15439 15453
rect 15562 15444 15568 15456
rect 15620 15444 15626 15496
rect 15838 15484 15844 15496
rect 15799 15456 15844 15484
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 17954 15484 17960 15496
rect 17915 15456 17960 15484
rect 17954 15444 17960 15456
rect 18012 15444 18018 15496
rect 20622 15444 20628 15496
rect 20680 15484 20686 15496
rect 20993 15487 21051 15493
rect 20993 15484 21005 15487
rect 20680 15456 21005 15484
rect 20680 15444 20686 15456
rect 20993 15453 21005 15456
rect 21039 15484 21051 15487
rect 21358 15484 21364 15496
rect 21039 15456 21364 15484
rect 21039 15453 21051 15456
rect 20993 15447 21051 15453
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15484 21695 15487
rect 21726 15484 21732 15496
rect 21683 15456 21732 15484
rect 21683 15453 21695 15456
rect 21637 15447 21695 15453
rect 21726 15444 21732 15456
rect 21784 15444 21790 15496
rect 1486 15376 1492 15428
rect 1544 15416 1550 15428
rect 2038 15416 2044 15428
rect 1544 15388 2044 15416
rect 1544 15376 1550 15388
rect 2038 15376 2044 15388
rect 2096 15376 2102 15428
rect 8294 15376 8300 15428
rect 8352 15416 8358 15428
rect 8757 15419 8815 15425
rect 8757 15416 8769 15419
rect 8352 15388 8769 15416
rect 8352 15376 8358 15388
rect 8757 15385 8769 15388
rect 8803 15416 8815 15419
rect 12802 15416 12808 15428
rect 8803 15388 12808 15416
rect 8803 15385 8815 15388
rect 8757 15379 8815 15385
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 18877 15419 18935 15425
rect 18877 15385 18889 15419
rect 18923 15416 18935 15419
rect 21082 15416 21088 15428
rect 18923 15388 21088 15416
rect 18923 15385 18935 15388
rect 18877 15379 18935 15385
rect 21082 15376 21088 15388
rect 21140 15416 21146 15428
rect 21542 15416 21548 15428
rect 21140 15388 21548 15416
rect 21140 15376 21146 15388
rect 21542 15376 21548 15388
rect 21600 15376 21606 15428
rect 8386 15348 8392 15360
rect 8347 15320 8392 15348
rect 8386 15308 8392 15320
rect 8444 15308 8450 15360
rect 9306 15348 9312 15360
rect 9267 15320 9312 15348
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 9950 15308 9956 15360
rect 10008 15348 10014 15360
rect 10781 15351 10839 15357
rect 10781 15348 10793 15351
rect 10008 15320 10793 15348
rect 10008 15308 10014 15320
rect 10781 15317 10793 15320
rect 10827 15348 10839 15351
rect 12066 15348 12072 15360
rect 10827 15320 12072 15348
rect 10827 15317 10839 15320
rect 10781 15311 10839 15317
rect 12066 15308 12072 15320
rect 12124 15308 12130 15360
rect 19150 15348 19156 15360
rect 19111 15320 19156 15348
rect 19150 15308 19156 15320
rect 19208 15308 19214 15360
rect 19843 15351 19901 15357
rect 19843 15317 19855 15351
rect 19889 15348 19901 15351
rect 20438 15348 20444 15360
rect 19889 15320 20444 15348
rect 19889 15317 19901 15320
rect 19843 15311 19901 15317
rect 20438 15308 20444 15320
rect 20496 15308 20502 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 9217 15147 9275 15153
rect 9217 15113 9229 15147
rect 9263 15144 9275 15147
rect 9766 15144 9772 15156
rect 9263 15116 9772 15144
rect 9263 15113 9275 15116
rect 9217 15107 9275 15113
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 10134 15104 10140 15156
rect 10192 15144 10198 15156
rect 10229 15147 10287 15153
rect 10229 15144 10241 15147
rect 10192 15116 10241 15144
rect 10192 15104 10198 15116
rect 10229 15113 10241 15116
rect 10275 15113 10287 15147
rect 10502 15144 10508 15156
rect 10463 15116 10508 15144
rect 10229 15107 10287 15113
rect 10502 15104 10508 15116
rect 10560 15104 10566 15156
rect 10962 15104 10968 15156
rect 11020 15144 11026 15156
rect 11149 15147 11207 15153
rect 11149 15144 11161 15147
rect 11020 15116 11161 15144
rect 11020 15104 11026 15116
rect 11149 15113 11161 15116
rect 11195 15113 11207 15147
rect 11149 15107 11207 15113
rect 13633 15147 13691 15153
rect 13633 15113 13645 15147
rect 13679 15144 13691 15147
rect 13722 15144 13728 15156
rect 13679 15116 13728 15144
rect 13679 15113 13691 15116
rect 13633 15107 13691 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 13909 15147 13967 15153
rect 13909 15144 13921 15147
rect 13872 15116 13921 15144
rect 13872 15104 13878 15116
rect 13909 15113 13921 15116
rect 13955 15113 13967 15147
rect 13909 15107 13967 15113
rect 15197 15147 15255 15153
rect 15197 15113 15209 15147
rect 15243 15144 15255 15147
rect 15470 15144 15476 15156
rect 15243 15116 15476 15144
rect 15243 15113 15255 15116
rect 15197 15107 15255 15113
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 15562 15104 15568 15156
rect 15620 15144 15626 15156
rect 17037 15147 17095 15153
rect 17037 15144 17049 15147
rect 15620 15116 17049 15144
rect 15620 15104 15626 15116
rect 17037 15113 17049 15116
rect 17083 15113 17095 15147
rect 17037 15107 17095 15113
rect 17497 15147 17555 15153
rect 17497 15113 17509 15147
rect 17543 15144 17555 15147
rect 17954 15144 17960 15156
rect 17543 15116 17960 15144
rect 17543 15113 17555 15116
rect 17497 15107 17555 15113
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 18187 15147 18245 15153
rect 18187 15113 18199 15147
rect 18233 15144 18245 15147
rect 18782 15144 18788 15156
rect 18233 15116 18788 15144
rect 18233 15113 18245 15116
rect 18187 15107 18245 15113
rect 18782 15104 18788 15116
rect 18840 15104 18846 15156
rect 19981 15147 20039 15153
rect 19981 15113 19993 15147
rect 20027 15144 20039 15147
rect 20990 15144 20996 15156
rect 20027 15116 20996 15144
rect 20027 15113 20039 15116
rect 19981 15107 20039 15113
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 21358 15104 21364 15156
rect 21416 15144 21422 15156
rect 22370 15144 22376 15156
rect 21416 15116 22376 15144
rect 21416 15104 21422 15116
rect 22370 15104 22376 15116
rect 22428 15104 22434 15156
rect 8435 15079 8493 15085
rect 8435 15045 8447 15079
rect 8481 15076 8493 15079
rect 9122 15076 9128 15088
rect 8481 15048 9128 15076
rect 8481 15045 8493 15048
rect 8435 15039 8493 15045
rect 9122 15036 9128 15048
rect 9180 15036 9186 15088
rect 14737 15079 14795 15085
rect 14737 15045 14749 15079
rect 14783 15076 14795 15079
rect 15580 15076 15608 15104
rect 22278 15076 22284 15088
rect 14783 15048 15608 15076
rect 16040 15048 22284 15076
rect 14783 15045 14795 15048
rect 14737 15039 14795 15045
rect 16040 15020 16068 15048
rect 22278 15036 22284 15048
rect 22336 15036 22342 15088
rect 8110 14968 8116 15020
rect 8168 15008 8174 15020
rect 12158 15008 12164 15020
rect 8168 14980 12164 15008
rect 8168 14968 8174 14980
rect 12158 14968 12164 14980
rect 12216 15008 12222 15020
rect 16022 15008 16028 15020
rect 12216 14980 16028 15008
rect 12216 14968 12222 14980
rect 8364 14943 8422 14949
rect 8364 14909 8376 14943
rect 8410 14940 8422 14943
rect 9306 14940 9312 14952
rect 8410 14912 8616 14940
rect 9267 14912 9312 14940
rect 8410 14909 8422 14912
rect 8364 14903 8422 14909
rect 8588 14816 8616 14912
rect 9306 14900 9312 14912
rect 9364 14900 9370 14952
rect 9766 14900 9772 14952
rect 9824 14940 9830 14952
rect 12452 14949 12480 14980
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 16206 15008 16212 15020
rect 16167 14980 16212 15008
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 19061 15011 19119 15017
rect 19061 14977 19073 15011
rect 19107 15008 19119 15011
rect 19150 15008 19156 15020
rect 19107 14980 19156 15008
rect 19107 14977 19119 14980
rect 19061 14971 19119 14977
rect 19150 14968 19156 14980
rect 19208 14968 19214 15020
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 15008 21143 15011
rect 21450 15008 21456 15020
rect 21131 14980 21456 15008
rect 21131 14977 21143 14980
rect 21085 14971 21143 14977
rect 21450 14968 21456 14980
rect 21508 15008 21514 15020
rect 22741 15011 22799 15017
rect 22741 15008 22753 15011
rect 21508 14980 22753 15008
rect 21508 14968 21514 14980
rect 22741 14977 22753 14980
rect 22787 14977 22799 15011
rect 22741 14971 22799 14977
rect 11384 14943 11442 14949
rect 11384 14940 11396 14943
rect 9824 14912 11396 14940
rect 9824 14900 9830 14912
rect 11384 14909 11396 14912
rect 11430 14940 11442 14943
rect 11793 14943 11851 14949
rect 11793 14940 11805 14943
rect 11430 14912 11805 14940
rect 11430 14909 11442 14912
rect 11384 14903 11442 14909
rect 11793 14909 11805 14912
rect 11839 14909 11851 14943
rect 11793 14903 11851 14909
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 12526 14900 12532 14952
rect 12584 14940 12590 14952
rect 12894 14940 12900 14952
rect 12584 14912 12900 14940
rect 12584 14900 12590 14912
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 17678 14900 17684 14952
rect 17736 14940 17742 14952
rect 18084 14943 18142 14949
rect 18084 14940 18096 14943
rect 17736 14912 18096 14940
rect 17736 14900 17742 14912
rect 18084 14909 18096 14912
rect 18130 14940 18142 14943
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18130 14912 18521 14940
rect 18130 14909 18142 14912
rect 18084 14903 18142 14909
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 19334 14940 19340 14952
rect 18509 14903 18567 14909
rect 19306 14900 19340 14940
rect 19392 14940 19398 14952
rect 19392 14912 19472 14940
rect 19392 14900 19398 14912
rect 11471 14875 11529 14881
rect 11471 14841 11483 14875
rect 11517 14872 11529 14875
rect 12986 14872 12992 14884
rect 11517 14844 12992 14872
rect 11517 14841 11529 14844
rect 11471 14835 11529 14841
rect 12986 14832 12992 14844
rect 13044 14832 13050 14884
rect 13170 14872 13176 14884
rect 13131 14844 13176 14872
rect 13170 14832 13176 14844
rect 13228 14832 13234 14884
rect 14182 14872 14188 14884
rect 14143 14844 14188 14872
rect 14182 14832 14188 14844
rect 14240 14832 14246 14884
rect 14277 14875 14335 14881
rect 14277 14841 14289 14875
rect 14323 14872 14335 14875
rect 15473 14875 15531 14881
rect 15473 14872 15485 14875
rect 14323 14844 15485 14872
rect 14323 14841 14335 14844
rect 14277 14835 14335 14841
rect 15473 14841 15485 14844
rect 15519 14841 15531 14875
rect 15746 14872 15752 14884
rect 15707 14844 15752 14872
rect 15473 14835 15531 14841
rect 1394 14764 1400 14816
rect 1452 14804 1458 14816
rect 1673 14807 1731 14813
rect 1673 14804 1685 14807
rect 1452 14776 1685 14804
rect 1452 14764 1458 14776
rect 1673 14773 1685 14776
rect 1719 14804 1731 14807
rect 5258 14804 5264 14816
rect 1719 14776 5264 14804
rect 1719 14773 1731 14776
rect 1673 14767 1731 14773
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 8570 14764 8576 14816
rect 8628 14804 8634 14816
rect 8757 14807 8815 14813
rect 8757 14804 8769 14807
rect 8628 14776 8769 14804
rect 8628 14764 8634 14776
rect 8757 14773 8769 14776
rect 8803 14773 8815 14807
rect 9674 14804 9680 14816
rect 9635 14776 9680 14804
rect 8757 14767 8815 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 14292 14804 14320 14835
rect 13872 14776 14320 14804
rect 15488 14804 15516 14835
rect 15746 14832 15752 14844
rect 15804 14832 15810 14884
rect 15841 14875 15899 14881
rect 15841 14841 15853 14875
rect 15887 14841 15899 14875
rect 15841 14835 15899 14841
rect 15856 14804 15884 14835
rect 15488 14776 15884 14804
rect 13872 14764 13878 14776
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 16761 14807 16819 14813
rect 16761 14804 16773 14807
rect 15988 14776 16773 14804
rect 15988 14764 15994 14776
rect 16761 14773 16773 14776
rect 16807 14804 16819 14807
rect 16850 14804 16856 14816
rect 16807 14776 16856 14804
rect 16807 14773 16819 14776
rect 16761 14767 16819 14773
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 17770 14804 17776 14816
rect 17731 14776 17776 14804
rect 17770 14764 17776 14776
rect 17828 14764 17834 14816
rect 18969 14807 19027 14813
rect 18969 14773 18981 14807
rect 19015 14804 19027 14807
rect 19306 14804 19334 14900
rect 19444 14881 19472 14912
rect 19423 14875 19481 14881
rect 19423 14841 19435 14875
rect 19469 14841 19481 14875
rect 19423 14835 19481 14841
rect 20162 14832 20168 14884
rect 20220 14872 20226 14884
rect 21154 14875 21212 14881
rect 21154 14872 21166 14875
rect 20220 14844 21166 14872
rect 20220 14832 20226 14844
rect 21154 14841 21166 14844
rect 21200 14872 21212 14875
rect 21726 14872 21732 14884
rect 21200 14844 21312 14872
rect 21639 14844 21732 14872
rect 21200 14841 21212 14844
rect 21154 14835 21212 14841
rect 20254 14804 20260 14816
rect 19015 14776 19334 14804
rect 20215 14776 20260 14804
rect 19015 14773 19027 14776
rect 18969 14767 19027 14773
rect 20254 14764 20260 14776
rect 20312 14764 20318 14816
rect 20346 14764 20352 14816
rect 20404 14804 20410 14816
rect 20806 14804 20812 14816
rect 20404 14776 20812 14804
rect 20404 14764 20410 14776
rect 20806 14764 20812 14776
rect 20864 14764 20870 14816
rect 21284 14804 21312 14844
rect 21726 14832 21732 14844
rect 21784 14872 21790 14884
rect 24026 14872 24032 14884
rect 21784 14844 24032 14872
rect 21784 14832 21790 14844
rect 24026 14832 24032 14844
rect 24084 14832 24090 14884
rect 22005 14807 22063 14813
rect 22005 14804 22017 14807
rect 21284 14776 22017 14804
rect 22005 14773 22017 14776
rect 22051 14773 22063 14807
rect 22005 14767 22063 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 9858 14600 9864 14612
rect 9819 14572 9864 14600
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 10962 14560 10968 14612
rect 11020 14600 11026 14612
rect 11425 14603 11483 14609
rect 11425 14600 11437 14603
rect 11020 14572 11437 14600
rect 11020 14560 11026 14572
rect 11425 14569 11437 14572
rect 11471 14600 11483 14603
rect 11514 14600 11520 14612
rect 11471 14572 11520 14600
rect 11471 14569 11483 14572
rect 11425 14563 11483 14569
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 11698 14600 11704 14612
rect 11659 14572 11704 14600
rect 11698 14560 11704 14572
rect 11756 14600 11762 14612
rect 12250 14600 12256 14612
rect 11756 14572 12256 14600
rect 11756 14560 11762 14572
rect 12250 14560 12256 14572
rect 12308 14560 12314 14612
rect 12986 14600 12992 14612
rect 12947 14572 12992 14600
rect 12986 14560 12992 14572
rect 13044 14560 13050 14612
rect 13446 14600 13452 14612
rect 13407 14572 13452 14600
rect 13446 14560 13452 14572
rect 13504 14560 13510 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 14001 14603 14059 14609
rect 14001 14600 14013 14603
rect 13872 14572 14013 14600
rect 13872 14560 13878 14572
rect 14001 14569 14013 14572
rect 14047 14569 14059 14603
rect 15654 14600 15660 14612
rect 15615 14572 15660 14600
rect 14001 14563 14059 14569
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 16114 14560 16120 14612
rect 16172 14600 16178 14612
rect 16209 14603 16267 14609
rect 16209 14600 16221 14603
rect 16172 14572 16221 14600
rect 16172 14560 16178 14572
rect 16209 14569 16221 14572
rect 16255 14569 16267 14603
rect 16209 14563 16267 14569
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19429 14603 19487 14609
rect 19429 14600 19441 14603
rect 19392 14572 19441 14600
rect 19392 14560 19398 14572
rect 19429 14569 19441 14572
rect 19475 14569 19487 14603
rect 19429 14563 19487 14569
rect 19981 14603 20039 14609
rect 19981 14569 19993 14603
rect 20027 14600 20039 14603
rect 20346 14600 20352 14612
rect 20027 14572 20352 14600
rect 20027 14569 20039 14572
rect 19981 14563 20039 14569
rect 20346 14560 20352 14572
rect 20404 14560 20410 14612
rect 20438 14560 20444 14612
rect 20496 14600 20502 14612
rect 20625 14603 20683 14609
rect 20625 14600 20637 14603
rect 20496 14572 20637 14600
rect 20496 14560 20502 14572
rect 20625 14569 20637 14572
rect 20671 14600 20683 14603
rect 20671 14572 21036 14600
rect 20671 14569 20683 14572
rect 20625 14563 20683 14569
rect 9674 14492 9680 14544
rect 9732 14532 9738 14544
rect 10826 14535 10884 14541
rect 10826 14532 10838 14535
rect 9732 14504 10838 14532
rect 9732 14492 9738 14504
rect 10826 14501 10838 14504
rect 10872 14501 10884 14535
rect 10826 14495 10884 14501
rect 17773 14535 17831 14541
rect 17773 14501 17785 14535
rect 17819 14532 17831 14535
rect 17954 14532 17960 14544
rect 17819 14504 17960 14532
rect 17819 14501 17831 14504
rect 17773 14495 17831 14501
rect 17954 14492 17960 14504
rect 18012 14492 18018 14544
rect 21008 14541 21036 14572
rect 21358 14560 21364 14612
rect 21416 14600 21422 14612
rect 22557 14603 22615 14609
rect 22557 14600 22569 14603
rect 21416 14572 22569 14600
rect 21416 14560 21422 14572
rect 22557 14569 22569 14572
rect 22603 14569 22615 14603
rect 22557 14563 22615 14569
rect 20993 14535 21051 14541
rect 20993 14501 21005 14535
rect 21039 14501 21051 14535
rect 20993 14495 21051 14501
rect 21082 14492 21088 14544
rect 21140 14532 21146 14544
rect 21140 14504 21185 14532
rect 21140 14492 21146 14504
rect 22278 14492 22284 14544
rect 22336 14532 22342 14544
rect 22336 14504 22968 14532
rect 22336 14492 22342 14504
rect 8202 14464 8208 14476
rect 8163 14436 8208 14464
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 8386 14424 8392 14476
rect 8444 14464 8450 14476
rect 8573 14467 8631 14473
rect 8573 14464 8585 14467
rect 8444 14436 8585 14464
rect 8444 14424 8450 14436
rect 8573 14433 8585 14436
rect 8619 14464 8631 14467
rect 9030 14464 9036 14476
rect 8619 14436 9036 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 9030 14424 9036 14436
rect 9088 14424 9094 14476
rect 17310 14464 17316 14476
rect 17271 14436 17316 14464
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 17402 14424 17408 14476
rect 17460 14464 17466 14476
rect 17497 14467 17555 14473
rect 17497 14464 17509 14467
rect 17460 14436 17509 14464
rect 17460 14424 17466 14436
rect 17497 14433 17509 14436
rect 17543 14464 17555 14467
rect 20806 14464 20812 14476
rect 17543 14436 20812 14464
rect 17543 14433 17555 14436
rect 17497 14427 17555 14433
rect 20806 14424 20812 14436
rect 20864 14424 20870 14476
rect 21910 14424 21916 14476
rect 21968 14464 21974 14476
rect 22940 14473 22968 14504
rect 22465 14467 22523 14473
rect 22465 14464 22477 14467
rect 21968 14436 22477 14464
rect 21968 14424 21974 14436
rect 22465 14433 22477 14436
rect 22511 14433 22523 14467
rect 22465 14427 22523 14433
rect 22925 14467 22983 14473
rect 22925 14433 22937 14467
rect 22971 14433 22983 14467
rect 24026 14464 24032 14476
rect 23987 14436 24032 14464
rect 22925 14427 22983 14433
rect 24026 14424 24032 14436
rect 24084 14424 24090 14476
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14396 8815 14399
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 8803 14368 10517 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 10505 14365 10517 14368
rect 10551 14396 10563 14399
rect 10686 14396 10692 14408
rect 10551 14368 10692 14396
rect 10551 14365 10563 14368
rect 10505 14359 10563 14365
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 13081 14399 13139 14405
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 13170 14396 13176 14408
rect 13127 14368 13176 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 13170 14356 13176 14368
rect 13228 14356 13234 14408
rect 15289 14399 15347 14405
rect 15289 14365 15301 14399
rect 15335 14396 15347 14399
rect 15378 14396 15384 14408
rect 15335 14368 15384 14396
rect 15335 14365 15347 14368
rect 15289 14359 15347 14365
rect 15378 14356 15384 14368
rect 15436 14356 15442 14408
rect 19061 14399 19119 14405
rect 19061 14365 19073 14399
rect 19107 14365 19119 14399
rect 21266 14396 21272 14408
rect 21227 14368 21272 14396
rect 19061 14359 19119 14365
rect 9214 14260 9220 14272
rect 9175 14232 9220 14260
rect 9214 14220 9220 14232
rect 9272 14220 9278 14272
rect 12434 14260 12440 14272
rect 12395 14232 12440 14260
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 14182 14220 14188 14272
rect 14240 14260 14246 14272
rect 14277 14263 14335 14269
rect 14277 14260 14289 14263
rect 14240 14232 14289 14260
rect 14240 14220 14246 14232
rect 14277 14229 14289 14232
rect 14323 14229 14335 14263
rect 18046 14260 18052 14272
rect 18007 14232 18052 14260
rect 14277 14223 14335 14229
rect 18046 14220 18052 14232
rect 18104 14220 18110 14272
rect 18874 14260 18880 14272
rect 18835 14232 18880 14260
rect 18874 14220 18880 14232
rect 18932 14260 18938 14272
rect 19076 14260 19104 14359
rect 21266 14356 21272 14368
rect 21324 14356 21330 14408
rect 18932 14232 19104 14260
rect 18932 14220 18938 14232
rect 23750 14220 23756 14272
rect 23808 14260 23814 14272
rect 24167 14263 24225 14269
rect 24167 14260 24179 14263
rect 23808 14232 24179 14260
rect 23808 14220 23814 14232
rect 24167 14229 24179 14232
rect 24213 14229 24225 14263
rect 24167 14223 24225 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 9125 14059 9183 14065
rect 9125 14025 9137 14059
rect 9171 14056 9183 14059
rect 9674 14056 9680 14068
rect 9171 14028 9680 14056
rect 9171 14025 9183 14028
rect 9125 14019 9183 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 10042 14016 10048 14068
rect 10100 14056 10106 14068
rect 10137 14059 10195 14065
rect 10137 14056 10149 14059
rect 10100 14028 10149 14056
rect 10100 14016 10106 14028
rect 10137 14025 10149 14028
rect 10183 14025 10195 14059
rect 11422 14056 11428 14068
rect 11383 14028 11428 14056
rect 10137 14019 10195 14025
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 12158 14056 12164 14068
rect 12119 14028 12164 14056
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 13446 14056 13452 14068
rect 13407 14028 13452 14056
rect 13446 14016 13452 14028
rect 13504 14056 13510 14068
rect 14001 14059 14059 14065
rect 14001 14056 14013 14059
rect 13504 14028 14013 14056
rect 13504 14016 13510 14028
rect 14001 14025 14013 14028
rect 14047 14056 14059 14059
rect 14093 14059 14151 14065
rect 14093 14056 14105 14059
rect 14047 14028 14105 14056
rect 14047 14025 14059 14028
rect 14001 14019 14059 14025
rect 14093 14025 14105 14028
rect 14139 14025 14151 14059
rect 14093 14019 14151 14025
rect 15197 14059 15255 14065
rect 15197 14025 15209 14059
rect 15243 14056 15255 14059
rect 15470 14056 15476 14068
rect 15243 14028 15476 14056
rect 15243 14025 15255 14028
rect 15197 14019 15255 14025
rect 15470 14016 15476 14028
rect 15528 14016 15534 14068
rect 16022 14016 16028 14068
rect 16080 14056 16086 14068
rect 16080 14028 16896 14056
rect 16080 14016 16086 14028
rect 9692 13988 9720 14016
rect 10505 13991 10563 13997
rect 10505 13988 10517 13991
rect 9692 13960 10517 13988
rect 9214 13920 9220 13932
rect 9175 13892 9220 13920
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 1946 13852 1952 13864
rect 1443 13824 1952 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 7926 13852 7932 13864
rect 7887 13824 7932 13852
rect 7926 13812 7932 13824
rect 7984 13812 7990 13864
rect 8110 13852 8116 13864
rect 8023 13824 8116 13852
rect 8110 13812 8116 13824
rect 8168 13852 8174 13864
rect 9692 13852 9720 13960
rect 10505 13957 10517 13960
rect 10551 13988 10563 13991
rect 10870 13988 10876 14000
rect 10551 13960 10876 13988
rect 10551 13957 10563 13960
rect 10505 13951 10563 13957
rect 10870 13948 10876 13960
rect 10928 13948 10934 14000
rect 13630 13988 13636 14000
rect 13004 13960 13636 13988
rect 8168 13824 8193 13852
rect 9416 13824 9720 13852
rect 11032 13855 11090 13861
rect 8168 13812 8174 13824
rect 7561 13787 7619 13793
rect 7561 13753 7573 13787
rect 7607 13784 7619 13787
rect 8128 13784 8156 13812
rect 8386 13784 8392 13796
rect 7607 13756 8156 13784
rect 8347 13756 8392 13784
rect 7607 13753 7619 13756
rect 7561 13747 7619 13753
rect 8386 13744 8392 13756
rect 8444 13744 8450 13796
rect 9416 13784 9444 13824
rect 11032 13821 11044 13855
rect 11078 13852 11090 13855
rect 11422 13852 11428 13864
rect 11078 13824 11428 13852
rect 11078 13821 11090 13824
rect 11032 13815 11090 13821
rect 11422 13812 11428 13824
rect 11480 13812 11486 13864
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 13004 13861 13032 13960
rect 13630 13948 13636 13960
rect 13688 13948 13694 14000
rect 16209 13991 16267 13997
rect 16209 13988 16221 13991
rect 13786 13960 16221 13988
rect 13078 13880 13084 13932
rect 13136 13920 13142 13932
rect 13786 13920 13814 13960
rect 16209 13957 16221 13960
rect 16255 13988 16267 13991
rect 16868 13988 16896 14028
rect 17310 14016 17316 14068
rect 17368 14056 17374 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 17368 14028 17785 14056
rect 17368 14016 17374 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 18230 14056 18236 14068
rect 18191 14028 18236 14056
rect 17773 14019 17831 14025
rect 18230 14016 18236 14028
rect 18288 14016 18294 14068
rect 20162 14056 20168 14068
rect 18340 14028 19334 14056
rect 20123 14028 20168 14056
rect 17494 13988 17500 14000
rect 16255 13960 16804 13988
rect 16868 13960 17500 13988
rect 16255 13957 16267 13960
rect 16209 13951 16267 13957
rect 13136 13892 13814 13920
rect 13136 13880 13142 13892
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12216 13824 12449 13852
rect 12216 13812 12222 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 12989 13855 13047 13861
rect 12989 13821 13001 13855
rect 13035 13821 13047 13855
rect 14274 13852 14280 13864
rect 14235 13824 14280 13852
rect 12989 13815 13047 13821
rect 14274 13812 14280 13824
rect 14332 13812 14338 13864
rect 15933 13855 15991 13861
rect 15933 13821 15945 13855
rect 15979 13852 15991 13855
rect 16393 13855 16451 13861
rect 16393 13852 16405 13855
rect 15979 13824 16405 13852
rect 15979 13821 15991 13824
rect 15933 13815 15991 13821
rect 16393 13821 16405 13824
rect 16439 13852 16451 13855
rect 16666 13852 16672 13864
rect 16439 13824 16672 13852
rect 16439 13821 16451 13824
rect 16393 13815 16451 13821
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 16776 13852 16804 13960
rect 17494 13948 17500 13960
rect 17552 13988 17558 14000
rect 18340 13988 18368 14028
rect 17552 13960 18368 13988
rect 19306 13988 19334 14028
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 22278 14016 22284 14068
rect 22336 14056 22342 14068
rect 22373 14059 22431 14065
rect 22373 14056 22385 14059
rect 22336 14028 22385 14056
rect 22336 14016 22342 14028
rect 22373 14025 22385 14028
rect 22419 14025 22431 14059
rect 22373 14019 22431 14025
rect 22922 14016 22928 14068
rect 22980 14056 22986 14068
rect 23017 14059 23075 14065
rect 23017 14056 23029 14059
rect 22980 14028 23029 14056
rect 22980 14016 22986 14028
rect 23017 14025 23029 14028
rect 23063 14025 23075 14059
rect 23017 14019 23075 14025
rect 24213 14059 24271 14065
rect 24213 14025 24225 14059
rect 24259 14056 24271 14059
rect 24854 14056 24860 14068
rect 24259 14028 24860 14056
rect 24259 14025 24271 14028
rect 24213 14019 24271 14025
rect 20441 13991 20499 13997
rect 20441 13988 20453 13991
rect 19306 13960 20453 13988
rect 17552 13948 17558 13960
rect 20441 13957 20453 13960
rect 20487 13988 20499 13991
rect 20487 13960 20944 13988
rect 20487 13957 20499 13960
rect 20441 13951 20499 13957
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 18874 13920 18880 13932
rect 17175 13892 18880 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 18874 13880 18880 13892
rect 18932 13880 18938 13932
rect 19444 13892 20576 13920
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 16776 13824 16865 13852
rect 16853 13821 16865 13824
rect 16899 13852 16911 13855
rect 17402 13852 17408 13864
rect 16899 13824 17408 13852
rect 16899 13821 16911 13824
rect 16853 13815 16911 13821
rect 17402 13812 17408 13824
rect 17460 13812 17466 13864
rect 17957 13855 18015 13861
rect 17957 13821 17969 13855
rect 18003 13852 18015 13855
rect 18046 13852 18052 13864
rect 18003 13824 18052 13852
rect 18003 13821 18015 13824
rect 17957 13815 18015 13821
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 19241 13855 19299 13861
rect 19241 13821 19253 13855
rect 19287 13821 19299 13855
rect 19241 13815 19299 13821
rect 9538 13787 9596 13793
rect 9538 13784 9550 13787
rect 9416 13756 9550 13784
rect 9538 13753 9550 13756
rect 9584 13753 9596 13787
rect 11330 13784 11336 13796
rect 9538 13747 9596 13753
rect 9646 13756 11336 13784
rect 9646 13728 9674 13756
rect 11330 13744 11336 13756
rect 11388 13744 11394 13796
rect 13078 13744 13084 13796
rect 13136 13784 13142 13796
rect 13173 13787 13231 13793
rect 13173 13784 13185 13787
rect 13136 13756 13185 13784
rect 13136 13744 13142 13756
rect 13173 13753 13185 13756
rect 13219 13753 13231 13787
rect 13173 13747 13231 13753
rect 14001 13787 14059 13793
rect 14001 13753 14013 13787
rect 14047 13784 14059 13787
rect 14639 13787 14697 13793
rect 14639 13784 14651 13787
rect 14047 13756 14651 13784
rect 14047 13753 14059 13756
rect 14001 13747 14059 13753
rect 14639 13753 14651 13756
rect 14685 13784 14697 13787
rect 15565 13787 15623 13793
rect 15565 13784 15577 13787
rect 14685 13756 15577 13784
rect 14685 13753 14697 13756
rect 14639 13747 14697 13753
rect 15565 13753 15577 13756
rect 15611 13784 15623 13787
rect 15654 13784 15660 13796
rect 15611 13756 15660 13784
rect 15611 13753 15623 13756
rect 15565 13747 15623 13753
rect 15654 13744 15660 13756
rect 15712 13744 15718 13796
rect 19254 13784 19282 13815
rect 19444 13784 19472 13892
rect 19254 13756 19472 13784
rect 19566 13787 19624 13793
rect 19566 13753 19578 13787
rect 19612 13753 19624 13787
rect 19566 13747 19624 13753
rect 7193 13719 7251 13725
rect 7193 13685 7205 13719
rect 7239 13716 7251 13719
rect 8202 13716 8208 13728
rect 7239 13688 8208 13716
rect 7239 13685 7251 13688
rect 7193 13679 7251 13685
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 8757 13719 8815 13725
rect 8757 13685 8769 13719
rect 8803 13716 8815 13719
rect 9030 13716 9036 13728
rect 8803 13688 9036 13716
rect 8803 13685 8815 13688
rect 8757 13679 8815 13685
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 9628 13676 9634 13728
rect 9686 13676 9692 13728
rect 10962 13676 10968 13728
rect 11020 13716 11026 13728
rect 11103 13719 11161 13725
rect 11103 13716 11115 13719
rect 11020 13688 11115 13716
rect 11020 13676 11026 13688
rect 11103 13685 11115 13688
rect 11149 13685 11161 13719
rect 11103 13679 11161 13685
rect 18785 13719 18843 13725
rect 18785 13685 18797 13719
rect 18831 13716 18843 13719
rect 19061 13719 19119 13725
rect 19061 13716 19073 13719
rect 18831 13688 19073 13716
rect 18831 13685 18843 13688
rect 18785 13679 18843 13685
rect 19061 13685 19073 13688
rect 19107 13716 19119 13719
rect 19334 13716 19340 13728
rect 19107 13688 19340 13716
rect 19107 13685 19119 13688
rect 19061 13679 19119 13685
rect 19334 13676 19340 13688
rect 19392 13716 19398 13728
rect 19581 13716 19609 13747
rect 19392 13688 19609 13716
rect 19392 13676 19398 13688
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 20548 13716 20576 13892
rect 20806 13852 20812 13864
rect 20719 13824 20812 13852
rect 20806 13812 20812 13824
rect 20864 13812 20870 13864
rect 20916 13852 20944 13960
rect 20993 13855 21051 13861
rect 20993 13852 21005 13855
rect 20916 13824 21005 13852
rect 20993 13821 21005 13824
rect 21039 13852 21051 13855
rect 21266 13852 21272 13864
rect 21039 13824 21272 13852
rect 21039 13821 21051 13824
rect 20993 13815 21051 13821
rect 21266 13812 21272 13824
rect 21324 13812 21330 13864
rect 21453 13855 21511 13861
rect 21453 13821 21465 13855
rect 21499 13852 21511 13855
rect 22624 13855 22682 13861
rect 21499 13824 21533 13852
rect 21499 13821 21511 13824
rect 21453 13815 21511 13821
rect 22624 13821 22636 13855
rect 22670 13852 22682 13855
rect 22922 13852 22928 13864
rect 22670 13824 22928 13852
rect 22670 13821 22682 13824
rect 22624 13815 22682 13821
rect 20824 13784 20852 13812
rect 21468 13784 21496 13815
rect 22922 13812 22928 13824
rect 22980 13812 22986 13864
rect 23728 13855 23786 13861
rect 23728 13821 23740 13855
rect 23774 13852 23786 13855
rect 24228 13852 24256 14019
rect 24854 14016 24860 14028
rect 24912 14016 24918 14068
rect 23774 13824 24256 13852
rect 23774 13821 23786 13824
rect 23728 13815 23786 13821
rect 20824 13756 21496 13784
rect 21910 13744 21916 13796
rect 21968 13784 21974 13796
rect 22005 13787 22063 13793
rect 22005 13784 22017 13787
rect 21968 13756 22017 13784
rect 21968 13744 21974 13756
rect 22005 13753 22017 13756
rect 22051 13784 22063 13787
rect 23290 13784 23296 13796
rect 22051 13756 23296 13784
rect 22051 13753 22063 13756
rect 22005 13747 22063 13753
rect 23290 13744 23296 13756
rect 23348 13744 23354 13796
rect 24026 13744 24032 13796
rect 24084 13784 24090 13796
rect 24489 13787 24547 13793
rect 24489 13784 24501 13787
rect 24084 13756 24501 13784
rect 24084 13744 24090 13756
rect 24489 13753 24501 13756
rect 24535 13753 24547 13787
rect 24489 13747 24547 13753
rect 21085 13719 21143 13725
rect 21085 13716 21097 13719
rect 20220 13688 21097 13716
rect 20220 13676 20226 13688
rect 21085 13685 21097 13688
rect 21131 13685 21143 13719
rect 21085 13679 21143 13685
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 22695 13719 22753 13725
rect 22695 13716 22707 13719
rect 22152 13688 22707 13716
rect 22152 13676 22158 13688
rect 22695 13685 22707 13688
rect 22741 13685 22753 13719
rect 22695 13679 22753 13685
rect 23658 13676 23664 13728
rect 23716 13716 23722 13728
rect 23799 13719 23857 13725
rect 23799 13716 23811 13719
rect 23716 13688 23811 13716
rect 23716 13676 23722 13688
rect 23799 13685 23811 13688
rect 23845 13685 23857 13719
rect 23799 13679 23857 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 9582 13512 9588 13524
rect 9180 13484 9588 13512
rect 9180 13472 9186 13484
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 10686 13512 10692 13524
rect 10647 13484 10692 13512
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 11057 13515 11115 13521
rect 11057 13512 11069 13515
rect 11020 13484 11069 13512
rect 11020 13472 11026 13484
rect 11057 13481 11069 13484
rect 11103 13481 11115 13515
rect 11057 13475 11115 13481
rect 13081 13515 13139 13521
rect 13081 13481 13093 13515
rect 13127 13512 13139 13515
rect 13170 13512 13176 13524
rect 13127 13484 13176 13512
rect 13127 13481 13139 13484
rect 13081 13475 13139 13481
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 20162 13512 20168 13524
rect 20123 13484 20168 13512
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 20717 13515 20775 13521
rect 20717 13481 20729 13515
rect 20763 13512 20775 13515
rect 20990 13512 20996 13524
rect 20763 13484 20996 13512
rect 20763 13481 20775 13484
rect 20717 13475 20775 13481
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 23658 13472 23664 13524
rect 23716 13512 23722 13524
rect 23753 13515 23811 13521
rect 23753 13512 23765 13515
rect 23716 13484 23765 13512
rect 23716 13472 23722 13484
rect 23753 13481 23765 13484
rect 23799 13481 23811 13515
rect 23753 13475 23811 13481
rect 7745 13447 7803 13453
rect 7745 13413 7757 13447
rect 7791 13444 7803 13447
rect 7926 13444 7932 13456
rect 7791 13416 7932 13444
rect 7791 13413 7803 13416
rect 7745 13407 7803 13413
rect 7926 13404 7932 13416
rect 7984 13444 7990 13456
rect 11330 13444 11336 13456
rect 7984 13416 9674 13444
rect 11291 13416 11336 13444
rect 7984 13404 7990 13416
rect 8018 13376 8024 13388
rect 7979 13348 8024 13376
rect 8018 13336 8024 13348
rect 8076 13336 8082 13388
rect 8110 13336 8116 13388
rect 8168 13376 8174 13388
rect 8481 13379 8539 13385
rect 8481 13376 8493 13379
rect 8168 13348 8493 13376
rect 8168 13336 8174 13348
rect 8481 13345 8493 13348
rect 8527 13345 8539 13379
rect 9646 13376 9674 13416
rect 11330 13404 11336 13416
rect 11388 13404 11394 13456
rect 11425 13447 11483 13453
rect 11425 13413 11437 13447
rect 11471 13444 11483 13447
rect 11514 13444 11520 13456
rect 11471 13416 11520 13444
rect 11471 13413 11483 13416
rect 11425 13407 11483 13413
rect 11514 13404 11520 13416
rect 11572 13444 11578 13456
rect 11790 13444 11796 13456
rect 11572 13416 11796 13444
rect 11572 13404 11578 13416
rect 11790 13404 11796 13416
rect 11848 13404 11854 13456
rect 12529 13447 12587 13453
rect 12529 13413 12541 13447
rect 12575 13444 12587 13447
rect 18049 13447 18107 13453
rect 12575 13416 13676 13444
rect 12575 13413 12587 13416
rect 12529 13407 12587 13413
rect 13648 13388 13676 13416
rect 14108 13416 17356 13444
rect 9950 13376 9956 13388
rect 9646 13348 9956 13376
rect 8481 13339 8539 13345
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10134 13376 10140 13388
rect 10095 13348 10140 13376
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 13173 13379 13231 13385
rect 13173 13376 13185 13379
rect 12860 13348 13185 13376
rect 12860 13336 12866 13348
rect 13173 13345 13185 13348
rect 13219 13345 13231 13379
rect 13630 13376 13636 13388
rect 13591 13348 13636 13376
rect 13173 13339 13231 13345
rect 8754 13308 8760 13320
rect 8715 13280 8760 13308
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 9272 13280 10241 13308
rect 9272 13268 9278 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 11609 13311 11667 13317
rect 11609 13308 11621 13311
rect 10229 13271 10287 13277
rect 11440 13280 11621 13308
rect 9858 13200 9864 13252
rect 9916 13240 9922 13252
rect 11440 13240 11468 13280
rect 11609 13277 11621 13280
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 9916 13212 11468 13240
rect 13188 13240 13216 13339
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 13722 13308 13728 13320
rect 13683 13280 13728 13308
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 14108 13240 14136 13416
rect 17328 13388 17356 13416
rect 18049 13413 18061 13447
rect 18095 13444 18107 13447
rect 19058 13444 19064 13456
rect 18095 13416 19064 13444
rect 18095 13413 18107 13416
rect 18049 13407 18107 13413
rect 19058 13404 19064 13416
rect 19116 13404 19122 13456
rect 19239 13447 19297 13453
rect 19239 13413 19251 13447
rect 19285 13444 19297 13447
rect 19334 13444 19340 13456
rect 19285 13416 19340 13444
rect 19285 13413 19297 13416
rect 19239 13407 19297 13413
rect 19334 13404 19340 13416
rect 19392 13404 19398 13456
rect 20806 13404 20812 13456
rect 20864 13444 20870 13456
rect 21085 13447 21143 13453
rect 21085 13444 21097 13447
rect 20864 13416 21097 13444
rect 20864 13404 20870 13416
rect 21085 13413 21097 13416
rect 21131 13413 21143 13447
rect 21085 13407 21143 13413
rect 22649 13447 22707 13453
rect 22649 13413 22661 13447
rect 22695 13444 22707 13447
rect 22830 13444 22836 13456
rect 22695 13416 22836 13444
rect 22695 13413 22707 13416
rect 22649 13407 22707 13413
rect 22830 13404 22836 13416
rect 22888 13404 22894 13456
rect 22922 13404 22928 13456
rect 22980 13444 22986 13456
rect 22980 13416 23025 13444
rect 22980 13404 22986 13416
rect 16022 13376 16028 13388
rect 15983 13348 16028 13376
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13376 16359 13379
rect 16574 13376 16580 13388
rect 16347 13348 16580 13376
rect 16347 13345 16359 13348
rect 16301 13339 16359 13345
rect 16574 13336 16580 13348
rect 16632 13336 16638 13388
rect 17310 13376 17316 13388
rect 17223 13348 17316 13376
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 17402 13336 17408 13388
rect 17460 13376 17466 13388
rect 17773 13379 17831 13385
rect 17773 13376 17785 13379
rect 17460 13348 17785 13376
rect 17460 13336 17466 13348
rect 17773 13345 17785 13348
rect 17819 13345 17831 13379
rect 17773 13339 17831 13345
rect 24648 13379 24706 13385
rect 24648 13345 24660 13379
rect 24694 13376 24706 13379
rect 24762 13376 24768 13388
rect 24694 13348 24768 13376
rect 24694 13345 24706 13348
rect 24648 13339 24706 13345
rect 24762 13336 24768 13348
rect 24820 13376 24826 13388
rect 26234 13376 26240 13388
rect 24820 13348 26240 13376
rect 24820 13336 24826 13348
rect 26234 13336 26240 13348
rect 26292 13336 26298 13388
rect 15378 13268 15384 13320
rect 15436 13308 15442 13320
rect 15473 13311 15531 13317
rect 15473 13308 15485 13311
rect 15436 13280 15485 13308
rect 15436 13268 15442 13280
rect 15473 13277 15485 13280
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 16485 13311 16543 13317
rect 16485 13277 16497 13311
rect 16531 13308 16543 13311
rect 18506 13308 18512 13320
rect 16531 13280 18512 13308
rect 16531 13277 16543 13280
rect 16485 13271 16543 13277
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 18874 13308 18880 13320
rect 18835 13280 18880 13308
rect 18874 13268 18880 13280
rect 18932 13268 18938 13320
rect 20622 13268 20628 13320
rect 20680 13308 20686 13320
rect 20993 13311 21051 13317
rect 20993 13308 21005 13311
rect 20680 13280 21005 13308
rect 20680 13268 20686 13280
rect 20993 13277 21005 13280
rect 21039 13277 21051 13311
rect 20993 13271 21051 13277
rect 21637 13311 21695 13317
rect 21637 13277 21649 13311
rect 21683 13308 21695 13311
rect 21726 13308 21732 13320
rect 21683 13280 21732 13308
rect 21683 13277 21695 13280
rect 21637 13271 21695 13277
rect 21726 13268 21732 13280
rect 21784 13268 21790 13320
rect 23477 13311 23535 13317
rect 23477 13277 23489 13311
rect 23523 13308 23535 13311
rect 24026 13308 24032 13320
rect 23523 13280 24032 13308
rect 23523 13277 23535 13280
rect 23477 13271 23535 13277
rect 24026 13268 24032 13280
rect 24084 13268 24090 13320
rect 14274 13240 14280 13252
rect 13188 13212 14136 13240
rect 14235 13212 14280 13240
rect 9916 13200 9922 13212
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 14642 13200 14648 13252
rect 14700 13240 14706 13252
rect 24719 13243 24777 13249
rect 24719 13240 24731 13243
rect 14700 13212 24731 13240
rect 14700 13200 14706 13212
rect 24719 13209 24731 13212
rect 24765 13209 24777 13243
rect 24719 13203 24777 13209
rect 9214 13172 9220 13184
rect 9175 13144 9220 13172
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 18417 13175 18475 13181
rect 18417 13141 18429 13175
rect 18463 13172 18475 13175
rect 18690 13172 18696 13184
rect 18463 13144 18696 13172
rect 18463 13141 18475 13144
rect 18417 13135 18475 13141
rect 18690 13132 18696 13144
rect 18748 13132 18754 13184
rect 19797 13175 19855 13181
rect 19797 13141 19809 13175
rect 19843 13172 19855 13175
rect 22646 13172 22652 13184
rect 19843 13144 22652 13172
rect 19843 13141 19855 13144
rect 19797 13135 19855 13141
rect 22646 13132 22652 13144
rect 22704 13132 22710 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 106 12928 112 12980
rect 164 12968 170 12980
rect 1581 12971 1639 12977
rect 1581 12968 1593 12971
rect 164 12940 1593 12968
rect 164 12928 170 12940
rect 1581 12937 1593 12940
rect 1627 12937 1639 12971
rect 8110 12968 8116 12980
rect 8071 12940 8116 12968
rect 1581 12931 1639 12937
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 11790 12968 11796 12980
rect 11751 12940 11796 12968
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 12802 12968 12808 12980
rect 12763 12940 12808 12968
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 12986 12928 12992 12980
rect 13044 12968 13050 12980
rect 13173 12971 13231 12977
rect 13173 12968 13185 12971
rect 13044 12940 13185 12968
rect 13044 12928 13050 12940
rect 13173 12937 13185 12940
rect 13219 12968 13231 12971
rect 13630 12968 13636 12980
rect 13219 12940 13636 12968
rect 13219 12937 13231 12940
rect 13173 12931 13231 12937
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 15930 12968 15936 12980
rect 13786 12940 15936 12968
rect 8018 12860 8024 12912
rect 8076 12900 8082 12912
rect 8481 12903 8539 12909
rect 8481 12900 8493 12903
rect 8076 12872 8493 12900
rect 8076 12860 8082 12872
rect 8481 12869 8493 12872
rect 8527 12900 8539 12903
rect 9214 12900 9220 12912
rect 8527 12872 9220 12900
rect 8527 12869 8539 12872
rect 8481 12863 8539 12869
rect 9214 12860 9220 12872
rect 9272 12900 9278 12912
rect 9272 12872 11284 12900
rect 9272 12860 9278 12872
rect 9508 12773 9536 12872
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 10962 12832 10968 12844
rect 10919 12804 10968 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 10962 12792 10968 12804
rect 11020 12792 11026 12844
rect 11256 12832 11284 12872
rect 11330 12860 11336 12912
rect 11388 12900 11394 12912
rect 12161 12903 12219 12909
rect 12161 12900 12173 12903
rect 11388 12872 12173 12900
rect 11388 12860 11394 12872
rect 12161 12869 12173 12872
rect 12207 12869 12219 12903
rect 12710 12900 12716 12912
rect 12161 12863 12219 12869
rect 12268 12872 12716 12900
rect 12268 12832 12296 12872
rect 12710 12860 12716 12872
rect 12768 12900 12774 12912
rect 13786 12900 13814 12940
rect 15930 12928 15936 12940
rect 15988 12928 15994 12980
rect 17402 12968 17408 12980
rect 17363 12940 17408 12968
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 18969 12971 19027 12977
rect 18969 12937 18981 12971
rect 19015 12968 19027 12971
rect 21082 12968 21088 12980
rect 19015 12940 21088 12968
rect 19015 12937 19027 12940
rect 18969 12931 19027 12937
rect 21082 12928 21088 12940
rect 21140 12968 21146 12980
rect 22373 12971 22431 12977
rect 22373 12968 22385 12971
rect 21140 12940 22385 12968
rect 21140 12928 21146 12940
rect 22373 12937 22385 12940
rect 22419 12968 22431 12971
rect 22922 12968 22928 12980
rect 22419 12940 22928 12968
rect 22419 12937 22431 12940
rect 22373 12931 22431 12937
rect 22922 12928 22928 12940
rect 22980 12928 22986 12980
rect 24762 12968 24768 12980
rect 24723 12940 24768 12968
rect 24762 12928 24768 12940
rect 24820 12928 24826 12980
rect 25409 12971 25467 12977
rect 25409 12937 25421 12971
rect 25455 12968 25467 12971
rect 27614 12968 27620 12980
rect 25455 12940 27620 12968
rect 25455 12937 25467 12940
rect 25409 12931 25467 12937
rect 27614 12928 27620 12940
rect 27672 12928 27678 12980
rect 12768 12872 13814 12900
rect 15473 12903 15531 12909
rect 12768 12860 12774 12872
rect 15473 12869 15485 12903
rect 15519 12900 15531 12903
rect 16022 12900 16028 12912
rect 15519 12872 16028 12900
rect 15519 12869 15531 12872
rect 15473 12863 15531 12869
rect 16022 12860 16028 12872
rect 16080 12900 16086 12912
rect 18046 12900 18052 12912
rect 16080 12872 18052 12900
rect 16080 12860 16086 12872
rect 18046 12860 18052 12872
rect 18104 12860 18110 12912
rect 19334 12860 19340 12912
rect 19392 12900 19398 12912
rect 20162 12900 20168 12912
rect 19392 12872 19437 12900
rect 20123 12872 20168 12900
rect 19392 12860 19398 12872
rect 20162 12860 20168 12872
rect 20220 12860 20226 12912
rect 23658 12860 23664 12912
rect 23716 12900 23722 12912
rect 23716 12872 23796 12900
rect 23716 12860 23722 12872
rect 13633 12835 13691 12841
rect 13633 12832 13645 12835
rect 11256 12804 12296 12832
rect 12636 12804 13645 12832
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 9493 12767 9551 12773
rect 1443 12736 2084 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 2056 12640 2084 12736
rect 9493 12733 9505 12767
rect 9539 12733 9551 12767
rect 9674 12764 9680 12776
rect 9635 12736 9680 12764
rect 9493 12727 9551 12733
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 9030 12656 9036 12708
rect 9088 12696 9094 12708
rect 9125 12699 9183 12705
rect 9125 12696 9137 12699
rect 9088 12668 9137 12696
rect 9088 12656 9094 12668
rect 9125 12665 9137 12668
rect 9171 12696 9183 12699
rect 9692 12696 9720 12724
rect 12636 12708 12664 12804
rect 13633 12801 13645 12804
rect 13679 12832 13691 12835
rect 14918 12832 14924 12844
rect 13679 12804 14924 12832
rect 13679 12801 13691 12804
rect 13633 12795 13691 12801
rect 14918 12792 14924 12804
rect 14976 12792 14982 12844
rect 16666 12792 16672 12844
rect 16724 12832 16730 12844
rect 16724 12804 18822 12832
rect 16724 12792 16730 12804
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 16574 12764 16580 12776
rect 16347 12736 16580 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 16758 12724 16764 12776
rect 16816 12764 16822 12776
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 16816 12736 16865 12764
rect 16816 12724 16822 12736
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12764 18107 12767
rect 18690 12764 18696 12776
rect 18095 12736 18696 12764
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 18794 12764 18822 12804
rect 18874 12792 18880 12844
rect 18932 12832 18938 12844
rect 19705 12835 19763 12841
rect 19705 12832 19717 12835
rect 18932 12804 19717 12832
rect 18932 12792 18938 12804
rect 19705 12801 19717 12804
rect 19751 12832 19763 12835
rect 20254 12832 20260 12844
rect 19751 12804 20260 12832
rect 19751 12801 19763 12804
rect 19705 12795 19763 12801
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 21085 12835 21143 12841
rect 21085 12832 21097 12835
rect 20404 12804 21097 12832
rect 20404 12792 20410 12804
rect 21085 12801 21097 12804
rect 21131 12832 21143 12835
rect 22094 12832 22100 12844
rect 21131 12804 22100 12832
rect 21131 12801 21143 12804
rect 21085 12795 21143 12801
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 22370 12792 22376 12844
rect 22428 12832 22434 12844
rect 23768 12841 23796 12872
rect 23017 12835 23075 12841
rect 23017 12832 23029 12835
rect 22428 12804 23029 12832
rect 22428 12792 22434 12804
rect 19832 12767 19890 12773
rect 19832 12764 19844 12767
rect 18794 12736 19844 12764
rect 19832 12733 19844 12736
rect 19878 12733 19890 12767
rect 19832 12727 19890 12733
rect 10134 12696 10140 12708
rect 9171 12668 10140 12696
rect 9171 12665 9183 12668
rect 9125 12659 9183 12665
rect 10134 12656 10140 12668
rect 10192 12696 10198 12708
rect 10229 12699 10287 12705
rect 10229 12696 10241 12699
rect 10192 12668 10241 12696
rect 10192 12656 10198 12668
rect 10229 12665 10241 12668
rect 10275 12665 10287 12699
rect 10229 12659 10287 12665
rect 10689 12699 10747 12705
rect 10689 12665 10701 12699
rect 10735 12696 10747 12699
rect 10962 12696 10968 12708
rect 10735 12668 10968 12696
rect 10735 12665 10747 12668
rect 10689 12659 10747 12665
rect 10962 12656 10968 12668
rect 11020 12656 11026 12708
rect 11517 12699 11575 12705
rect 11517 12665 11529 12699
rect 11563 12696 11575 12699
rect 12618 12696 12624 12708
rect 11563 12668 12624 12696
rect 11563 12665 11575 12668
rect 11517 12659 11575 12665
rect 12618 12656 12624 12668
rect 12676 12656 12682 12708
rect 13357 12699 13415 12705
rect 13357 12665 13369 12699
rect 13403 12665 13415 12699
rect 13357 12659 13415 12665
rect 2038 12628 2044 12640
rect 1999 12600 2044 12628
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 9306 12628 9312 12640
rect 9267 12600 9312 12628
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 13372 12628 13400 12659
rect 13446 12656 13452 12708
rect 13504 12696 13510 12708
rect 15013 12699 15071 12705
rect 13504 12668 13549 12696
rect 13504 12656 13510 12668
rect 15013 12665 15025 12699
rect 15059 12665 15071 12699
rect 15013 12659 15071 12665
rect 17129 12699 17187 12705
rect 17129 12665 17141 12699
rect 17175 12696 17187 12699
rect 18138 12696 18144 12708
rect 17175 12668 18144 12696
rect 17175 12665 17187 12668
rect 17129 12659 17187 12665
rect 13906 12628 13912 12640
rect 13372 12600 13912 12628
rect 13906 12588 13912 12600
rect 13964 12628 13970 12640
rect 14642 12628 14648 12640
rect 13964 12600 14648 12628
rect 13964 12588 13970 12600
rect 14642 12588 14648 12600
rect 14700 12588 14706 12640
rect 14737 12631 14795 12637
rect 14737 12597 14749 12631
rect 14783 12628 14795 12631
rect 14826 12628 14832 12640
rect 14783 12600 14832 12628
rect 14783 12597 14795 12600
rect 14737 12591 14795 12597
rect 14826 12588 14832 12600
rect 14884 12628 14890 12640
rect 15028 12628 15056 12659
rect 18138 12656 18144 12668
rect 18196 12656 18202 12708
rect 18370 12699 18428 12705
rect 18370 12665 18382 12699
rect 18416 12665 18428 12699
rect 19857 12696 19885 12727
rect 20070 12724 20076 12776
rect 20128 12764 20134 12776
rect 20806 12764 20812 12776
rect 20128 12736 20812 12764
rect 20128 12724 20134 12736
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 22526 12764 22554 12804
rect 23017 12801 23029 12804
rect 23063 12801 23075 12835
rect 23017 12795 23075 12801
rect 23753 12835 23811 12841
rect 23753 12801 23765 12835
rect 23799 12801 23811 12835
rect 24026 12832 24032 12844
rect 23987 12804 24032 12832
rect 23753 12795 23811 12801
rect 24026 12792 24032 12804
rect 24084 12792 24090 12844
rect 22592 12767 22650 12773
rect 22592 12764 22604 12767
rect 22526 12736 22604 12764
rect 22592 12733 22604 12736
rect 22638 12733 22650 12767
rect 22592 12727 22650 12733
rect 24854 12724 24860 12776
rect 24912 12764 24918 12776
rect 25225 12767 25283 12773
rect 25225 12764 25237 12767
rect 24912 12736 25237 12764
rect 24912 12724 24918 12736
rect 25225 12733 25237 12736
rect 25271 12764 25283 12767
rect 25777 12767 25835 12773
rect 25777 12764 25789 12767
rect 25271 12736 25789 12764
rect 25271 12733 25283 12736
rect 25225 12727 25283 12733
rect 25777 12733 25789 12736
rect 25823 12733 25835 12767
rect 25777 12727 25835 12733
rect 20257 12699 20315 12705
rect 20257 12696 20269 12699
rect 19857 12668 20269 12696
rect 18370 12659 18428 12665
rect 20257 12665 20269 12668
rect 20303 12665 20315 12699
rect 20257 12659 20315 12665
rect 17862 12628 17868 12640
rect 14884 12600 15056 12628
rect 17823 12600 17868 12628
rect 14884 12588 14890 12600
rect 17862 12588 17868 12600
rect 17920 12628 17926 12640
rect 18385 12628 18413 12659
rect 20438 12656 20444 12708
rect 20496 12696 20502 12708
rect 21177 12699 21235 12705
rect 21177 12696 21189 12699
rect 20496 12668 21189 12696
rect 20496 12656 20502 12668
rect 21177 12665 21189 12668
rect 21223 12696 21235 12699
rect 21726 12696 21732 12708
rect 21223 12668 21404 12696
rect 21687 12668 21732 12696
rect 21223 12665 21235 12668
rect 21177 12659 21235 12665
rect 17920 12600 18413 12628
rect 19935 12631 19993 12637
rect 17920 12588 17926 12600
rect 19935 12597 19947 12631
rect 19981 12628 19993 12631
rect 20162 12628 20168 12640
rect 19981 12600 20168 12628
rect 19981 12597 19993 12600
rect 19935 12591 19993 12597
rect 20162 12588 20168 12600
rect 20220 12588 20226 12640
rect 21376 12628 21404 12668
rect 21726 12656 21732 12668
rect 21784 12656 21790 12708
rect 22278 12656 22284 12708
rect 22336 12696 22342 12708
rect 23385 12699 23443 12705
rect 23385 12696 23397 12699
rect 22336 12668 23397 12696
rect 22336 12656 22342 12668
rect 23385 12665 23397 12668
rect 23431 12696 23443 12699
rect 23845 12699 23903 12705
rect 23845 12696 23857 12699
rect 23431 12668 23857 12696
rect 23431 12665 23443 12668
rect 23385 12659 23443 12665
rect 23845 12665 23857 12668
rect 23891 12665 23903 12699
rect 23845 12659 23903 12665
rect 22005 12631 22063 12637
rect 22005 12628 22017 12631
rect 21376 12600 22017 12628
rect 22005 12597 22017 12600
rect 22051 12628 22063 12631
rect 22186 12628 22192 12640
rect 22051 12600 22192 12628
rect 22051 12597 22063 12600
rect 22005 12591 22063 12597
rect 22186 12588 22192 12600
rect 22244 12588 22250 12640
rect 22695 12631 22753 12637
rect 22695 12597 22707 12631
rect 22741 12628 22753 12631
rect 22922 12628 22928 12640
rect 22741 12600 22928 12628
rect 22741 12597 22753 12600
rect 22695 12591 22753 12597
rect 22922 12588 22928 12600
rect 22980 12588 22986 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 10870 12424 10876 12436
rect 10831 12396 10876 12424
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 10962 12384 10968 12436
rect 11020 12424 11026 12436
rect 11425 12427 11483 12433
rect 11425 12424 11437 12427
rect 11020 12396 11437 12424
rect 11020 12384 11026 12396
rect 11425 12393 11437 12396
rect 11471 12393 11483 12427
rect 11425 12387 11483 12393
rect 11808 12396 13400 12424
rect 9950 12356 9956 12368
rect 9863 12328 9956 12356
rect 9950 12316 9956 12328
rect 10008 12356 10014 12368
rect 11808 12356 11836 12396
rect 10008 12328 11836 12356
rect 10008 12316 10014 12328
rect 11882 12316 11888 12368
rect 11940 12356 11946 12368
rect 12437 12359 12495 12365
rect 12437 12356 12449 12359
rect 11940 12328 12449 12356
rect 11940 12316 11946 12328
rect 12437 12325 12449 12328
rect 12483 12325 12495 12359
rect 13372 12356 13400 12396
rect 13538 12384 13544 12436
rect 13596 12424 13602 12436
rect 14001 12427 14059 12433
rect 14001 12424 14013 12427
rect 13596 12396 14013 12424
rect 13596 12384 13602 12396
rect 14001 12393 14013 12396
rect 14047 12393 14059 12427
rect 14001 12387 14059 12393
rect 14182 12384 14188 12436
rect 14240 12424 14246 12436
rect 14323 12427 14381 12433
rect 14323 12424 14335 12427
rect 14240 12396 14335 12424
rect 14240 12384 14246 12396
rect 14323 12393 14335 12396
rect 14369 12393 14381 12427
rect 14918 12424 14924 12436
rect 14879 12396 14924 12424
rect 14323 12387 14381 12393
rect 14918 12384 14924 12396
rect 14976 12384 14982 12436
rect 16758 12424 16764 12436
rect 15028 12396 16764 12424
rect 13630 12356 13636 12368
rect 13372 12328 13636 12356
rect 12437 12319 12495 12325
rect 13630 12316 13636 12328
rect 13688 12356 13694 12368
rect 15028 12356 15056 12396
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 17310 12424 17316 12436
rect 17271 12396 17316 12424
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 18601 12427 18659 12433
rect 18601 12393 18613 12427
rect 18647 12424 18659 12427
rect 20070 12424 20076 12436
rect 18647 12396 20076 12424
rect 18647 12393 18659 12396
rect 18601 12387 18659 12393
rect 20070 12384 20076 12396
rect 20128 12384 20134 12436
rect 20346 12424 20352 12436
rect 20307 12396 20352 12424
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 23014 12384 23020 12436
rect 23072 12424 23078 12436
rect 23072 12396 24256 12424
rect 23072 12384 23078 12396
rect 15470 12356 15476 12368
rect 13688 12328 15056 12356
rect 15431 12328 15476 12356
rect 13688 12316 13694 12328
rect 15470 12316 15476 12328
rect 15528 12316 15534 12368
rect 16022 12356 16028 12368
rect 15983 12328 16028 12356
rect 16022 12316 16028 12328
rect 16080 12316 16086 12368
rect 16393 12359 16451 12365
rect 16393 12325 16405 12359
rect 16439 12356 16451 12359
rect 16574 12356 16580 12368
rect 16439 12328 16580 12356
rect 16439 12325 16451 12328
rect 16393 12319 16451 12325
rect 8608 12291 8666 12297
rect 8608 12288 8620 12291
rect 8588 12257 8620 12288
rect 8654 12257 8666 12291
rect 8588 12251 8666 12257
rect 8711 12291 8769 12297
rect 8711 12257 8723 12291
rect 8757 12288 8769 12291
rect 13725 12291 13783 12297
rect 8757 12260 12204 12288
rect 8757 12257 8769 12260
rect 8711 12251 8769 12257
rect 8588 12152 8616 12251
rect 10505 12223 10563 12229
rect 10505 12220 10517 12223
rect 10336 12192 10517 12220
rect 8754 12152 8760 12164
rect 8588 12124 8760 12152
rect 8754 12112 8760 12124
rect 8812 12112 8818 12164
rect 8846 12112 8852 12164
rect 8904 12152 8910 12164
rect 9401 12155 9459 12161
rect 9401 12152 9413 12155
rect 8904 12124 9413 12152
rect 8904 12112 8910 12124
rect 9401 12121 9413 12124
rect 9447 12121 9459 12155
rect 9401 12115 9459 12121
rect 9125 12087 9183 12093
rect 9125 12053 9137 12087
rect 9171 12084 9183 12087
rect 9306 12084 9312 12096
rect 9171 12056 9312 12084
rect 9171 12053 9183 12056
rect 9125 12047 9183 12053
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 10042 12044 10048 12096
rect 10100 12084 10106 12096
rect 10336 12093 10364 12192
rect 10505 12189 10517 12192
rect 10551 12189 10563 12223
rect 12176 12220 12204 12260
rect 13725 12257 13737 12291
rect 13771 12288 13783 12291
rect 13906 12288 13912 12300
rect 13771 12260 13912 12288
rect 13771 12257 13783 12260
rect 13725 12251 13783 12257
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 14231 12291 14289 12297
rect 14231 12257 14243 12291
rect 14277 12257 14289 12291
rect 14231 12251 14289 12257
rect 12342 12220 12348 12232
rect 12176 12192 12348 12220
rect 10505 12183 10563 12189
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 12618 12220 12624 12232
rect 12579 12192 12624 12220
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14246 12220 14274 12251
rect 15378 12220 15384 12232
rect 13872 12192 14274 12220
rect 15339 12192 15384 12220
rect 13872 12180 13878 12192
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 11422 12112 11428 12164
rect 11480 12152 11486 12164
rect 16408 12152 16436 12319
rect 16574 12316 16580 12328
rect 16632 12316 16638 12368
rect 17862 12316 17868 12368
rect 17920 12356 17926 12368
rect 18002 12359 18060 12365
rect 18002 12356 18014 12359
rect 17920 12328 18014 12356
rect 17920 12316 17926 12328
rect 18002 12325 18014 12328
rect 18048 12325 18060 12359
rect 18002 12319 18060 12325
rect 20162 12316 20168 12368
rect 20220 12356 20226 12368
rect 20990 12356 20996 12368
rect 20220 12328 20996 12356
rect 20220 12316 20226 12328
rect 20990 12316 20996 12328
rect 21048 12316 21054 12368
rect 21082 12316 21088 12368
rect 21140 12356 21146 12368
rect 22646 12356 22652 12368
rect 21140 12328 21185 12356
rect 22607 12328 22652 12356
rect 21140 12316 21146 12328
rect 22646 12316 22652 12328
rect 22704 12316 22710 12368
rect 22922 12316 22928 12368
rect 22980 12356 22986 12368
rect 24228 12365 24256 12396
rect 24213 12359 24271 12365
rect 22980 12328 23474 12356
rect 22980 12316 22986 12328
rect 19864 12291 19922 12297
rect 19864 12257 19876 12291
rect 19910 12288 19922 12291
rect 19978 12288 19984 12300
rect 19910 12260 19984 12288
rect 19910 12257 19922 12260
rect 19864 12251 19922 12257
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 17681 12223 17739 12229
rect 17681 12189 17693 12223
rect 17727 12220 17739 12223
rect 18322 12220 18328 12232
rect 17727 12192 18328 12220
rect 17727 12189 17739 12192
rect 17681 12183 17739 12189
rect 18322 12180 18328 12192
rect 18380 12180 18386 12232
rect 21637 12223 21695 12229
rect 21637 12189 21649 12223
rect 21683 12220 21695 12223
rect 21726 12220 21732 12232
rect 21683 12192 21732 12220
rect 21683 12189 21695 12192
rect 21637 12183 21695 12189
rect 21726 12180 21732 12192
rect 21784 12220 21790 12232
rect 22554 12220 22560 12232
rect 21784 12192 22560 12220
rect 21784 12180 21790 12192
rect 22554 12180 22560 12192
rect 22612 12180 22618 12232
rect 22830 12220 22836 12232
rect 22791 12192 22836 12220
rect 22830 12180 22836 12192
rect 22888 12180 22894 12232
rect 23446 12220 23474 12328
rect 24213 12325 24225 12359
rect 24259 12356 24271 12359
rect 24762 12356 24768 12368
rect 24259 12328 24768 12356
rect 24259 12325 24271 12328
rect 24213 12319 24271 12325
rect 24762 12316 24768 12328
rect 24820 12316 24826 12368
rect 24118 12220 24124 12232
rect 23446 12192 24124 12220
rect 24118 12180 24124 12192
rect 24176 12180 24182 12232
rect 24210 12180 24216 12232
rect 24268 12220 24274 12232
rect 24397 12223 24455 12229
rect 24397 12220 24409 12223
rect 24268 12192 24409 12220
rect 24268 12180 24274 12192
rect 24397 12189 24409 12192
rect 24443 12189 24455 12223
rect 24397 12183 24455 12189
rect 11480 12124 16436 12152
rect 11480 12112 11486 12124
rect 16758 12112 16764 12164
rect 16816 12152 16822 12164
rect 19935 12155 19993 12161
rect 19935 12152 19947 12155
rect 16816 12124 19947 12152
rect 16816 12112 16822 12124
rect 19935 12121 19947 12124
rect 19981 12121 19993 12155
rect 19935 12115 19993 12121
rect 10321 12087 10379 12093
rect 10321 12084 10333 12087
rect 10100 12056 10333 12084
rect 10100 12044 10106 12056
rect 10321 12053 10333 12056
rect 10367 12053 10379 12087
rect 13354 12084 13360 12096
rect 13315 12056 13360 12084
rect 10321 12047 10379 12053
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 19610 12084 19616 12096
rect 19571 12056 19616 12084
rect 19610 12044 19616 12056
rect 19668 12044 19674 12096
rect 20622 12084 20628 12096
rect 20583 12056 20628 12084
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 23106 12044 23112 12096
rect 23164 12084 23170 12096
rect 23661 12087 23719 12093
rect 23661 12084 23673 12087
rect 23164 12056 23673 12084
rect 23164 12044 23170 12056
rect 23661 12053 23673 12056
rect 23707 12053 23719 12087
rect 23661 12047 23719 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 10137 11883 10195 11889
rect 10137 11849 10149 11883
rect 10183 11880 10195 11883
rect 10505 11883 10563 11889
rect 10505 11880 10517 11883
rect 10183 11852 10517 11880
rect 10183 11849 10195 11852
rect 10137 11843 10195 11849
rect 10505 11849 10517 11852
rect 10551 11880 10563 11883
rect 10870 11880 10876 11892
rect 10551 11852 10876 11880
rect 10551 11849 10563 11852
rect 10505 11843 10563 11849
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 11514 11880 11520 11892
rect 11427 11852 11520 11880
rect 11514 11840 11520 11852
rect 11572 11880 11578 11892
rect 11882 11880 11888 11892
rect 11572 11852 11888 11880
rect 11572 11840 11578 11852
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 13541 11883 13599 11889
rect 13541 11849 13553 11883
rect 13587 11880 13599 11883
rect 13722 11880 13728 11892
rect 13587 11852 13728 11880
rect 13587 11849 13599 11852
rect 13541 11843 13599 11849
rect 13722 11840 13728 11852
rect 13780 11880 13786 11892
rect 13780 11840 13814 11880
rect 14826 11840 14832 11892
rect 14884 11880 14890 11892
rect 14921 11883 14979 11889
rect 14921 11880 14933 11883
rect 14884 11852 14933 11880
rect 14884 11840 14890 11852
rect 14921 11849 14933 11852
rect 14967 11849 14979 11883
rect 14921 11843 14979 11849
rect 18647 11883 18705 11889
rect 18647 11849 18659 11883
rect 18693 11880 18705 11883
rect 20622 11880 20628 11892
rect 18693 11852 20628 11880
rect 18693 11849 18705 11852
rect 18647 11843 18705 11849
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 20898 11880 20904 11892
rect 20859 11852 20904 11880
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 20990 11840 20996 11892
rect 21048 11880 21054 11892
rect 21269 11883 21327 11889
rect 21269 11880 21281 11883
rect 21048 11852 21281 11880
rect 21048 11840 21054 11852
rect 21269 11849 21281 11852
rect 21315 11849 21327 11883
rect 21269 11843 21327 11849
rect 22646 11840 22652 11892
rect 22704 11880 22710 11892
rect 23017 11883 23075 11889
rect 23017 11880 23029 11883
rect 22704 11852 23029 11880
rect 22704 11840 22710 11852
rect 23017 11849 23029 11852
rect 23063 11849 23075 11883
rect 24762 11880 24768 11892
rect 23017 11843 23075 11849
rect 23446 11852 24440 11880
rect 24723 11852 24768 11880
rect 10888 11812 10916 11840
rect 10888 11784 11002 11812
rect 7926 11744 7932 11756
rect 7668 11716 7932 11744
rect 1486 11636 1492 11688
rect 1544 11676 1550 11688
rect 7668 11685 7696 11716
rect 7926 11704 7932 11716
rect 7984 11744 7990 11756
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 7984 11716 8493 11744
rect 7984 11704 7990 11716
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 9490 11744 9496 11756
rect 9451 11716 9496 11744
rect 8481 11707 8539 11713
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11744 10655 11747
rect 10870 11744 10876 11756
rect 10643 11716 10876 11744
rect 10643 11713 10655 11716
rect 10597 11707 10655 11713
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 7653 11679 7711 11685
rect 7653 11676 7665 11679
rect 1544 11648 7665 11676
rect 1544 11636 1550 11648
rect 7653 11645 7665 11648
rect 7699 11645 7711 11679
rect 7653 11639 7711 11645
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11645 7895 11679
rect 7837 11639 7895 11645
rect 7558 11540 7564 11552
rect 7519 11512 7564 11540
rect 7558 11500 7564 11512
rect 7616 11540 7622 11552
rect 7852 11540 7880 11639
rect 8846 11636 8852 11688
rect 8904 11676 8910 11688
rect 9033 11679 9091 11685
rect 9033 11676 9045 11679
rect 8904 11648 9045 11676
rect 8904 11636 8910 11648
rect 9033 11645 9045 11648
rect 9079 11645 9091 11679
rect 9033 11639 9091 11645
rect 9122 11636 9128 11688
rect 9180 11676 9186 11688
rect 9309 11679 9367 11685
rect 9180 11648 9225 11676
rect 9180 11636 9186 11648
rect 9309 11645 9321 11679
rect 9355 11676 9367 11679
rect 9398 11676 9404 11688
rect 9355 11648 9404 11676
rect 9355 11645 9367 11648
rect 9309 11639 9367 11645
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 8202 11608 8208 11620
rect 8163 11580 8208 11608
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 10974 11617 11002 11784
rect 13786 11744 13814 11840
rect 16022 11772 16028 11824
rect 16080 11812 16086 11824
rect 16393 11815 16451 11821
rect 16393 11812 16405 11815
rect 16080 11784 16405 11812
rect 16080 11772 16086 11784
rect 16393 11781 16405 11784
rect 16439 11781 16451 11815
rect 16393 11775 16451 11781
rect 19334 11772 19340 11824
rect 19392 11812 19398 11824
rect 19610 11812 19616 11824
rect 19392 11784 19437 11812
rect 19523 11784 19616 11812
rect 19392 11772 19398 11784
rect 14001 11747 14059 11753
rect 14001 11744 14013 11747
rect 13786 11716 14013 11744
rect 14001 11713 14013 11716
rect 14047 11713 14059 11747
rect 14001 11707 14059 11713
rect 15657 11747 15715 11753
rect 15657 11713 15669 11747
rect 15703 11744 15715 11747
rect 15841 11747 15899 11753
rect 15841 11744 15853 11747
rect 15703 11716 15853 11744
rect 15703 11713 15715 11716
rect 15657 11707 15715 11713
rect 15841 11713 15853 11716
rect 15887 11744 15899 11747
rect 18046 11744 18052 11756
rect 15887 11716 18052 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 19536 11753 19564 11784
rect 19610 11772 19616 11784
rect 19668 11812 19674 11824
rect 23446 11812 23474 11852
rect 24412 11824 24440 11852
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 19668 11784 23474 11812
rect 19668 11772 19674 11784
rect 23566 11772 23572 11824
rect 23624 11812 23630 11824
rect 24210 11812 24216 11824
rect 23624 11784 24216 11812
rect 23624 11772 23630 11784
rect 24210 11772 24216 11784
rect 24268 11812 24274 11824
rect 24305 11815 24363 11821
rect 24305 11812 24317 11815
rect 24268 11784 24317 11812
rect 24268 11772 24274 11784
rect 24305 11781 24317 11784
rect 24351 11781 24363 11815
rect 24305 11775 24363 11781
rect 24394 11772 24400 11824
rect 24452 11772 24458 11824
rect 19521 11747 19579 11753
rect 19521 11713 19533 11747
rect 19567 11713 19579 11747
rect 19521 11707 19579 11713
rect 21082 11704 21088 11756
rect 21140 11744 21146 11756
rect 22373 11747 22431 11753
rect 22373 11744 22385 11747
rect 21140 11716 22385 11744
rect 21140 11704 21146 11716
rect 22373 11713 22385 11716
rect 22419 11744 22431 11747
rect 23477 11747 23535 11753
rect 22419 11716 22784 11744
rect 22419 11713 22431 11716
rect 22373 11707 22431 11713
rect 12710 11676 12716 11688
rect 12671 11648 12716 11676
rect 12710 11636 12716 11648
rect 12768 11636 12774 11688
rect 12986 11676 12992 11688
rect 12947 11648 12992 11676
rect 12986 11636 12992 11648
rect 13044 11636 13050 11688
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11676 13231 11679
rect 13722 11676 13728 11688
rect 13219 11648 13728 11676
rect 13219 11645 13231 11648
rect 13173 11639 13231 11645
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 18598 11685 18604 11688
rect 18576 11679 18604 11685
rect 18576 11676 18588 11679
rect 18511 11648 18588 11676
rect 18576 11645 18588 11648
rect 18656 11676 18662 11688
rect 18969 11679 19027 11685
rect 18969 11676 18981 11679
rect 18656 11648 18981 11676
rect 18576 11639 18604 11645
rect 18598 11636 18604 11639
rect 18656 11636 18662 11648
rect 18969 11645 18981 11648
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 19334 11636 19340 11688
rect 19392 11676 19398 11688
rect 20438 11676 20444 11688
rect 19392 11648 19885 11676
rect 20399 11648 20444 11676
rect 19392 11636 19398 11648
rect 10959 11611 11017 11617
rect 10959 11577 10971 11611
rect 11005 11577 11017 11611
rect 10959 11571 11017 11577
rect 12253 11611 12311 11617
rect 12253 11577 12265 11611
rect 12299 11608 12311 11611
rect 12526 11608 12532 11620
rect 12299 11580 12532 11608
rect 12299 11577 12311 11580
rect 12253 11571 12311 11577
rect 12526 11568 12532 11580
rect 12584 11608 12590 11620
rect 13004 11608 13032 11636
rect 12584 11580 13032 11608
rect 12584 11568 12590 11580
rect 13538 11568 13544 11620
rect 13596 11608 13602 11620
rect 15933 11611 15991 11617
rect 13596 11580 14274 11608
rect 13596 11568 13602 11580
rect 7616 11512 7880 11540
rect 7616 11500 7622 11512
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 8849 11543 8907 11549
rect 8849 11540 8861 11543
rect 8812 11512 8861 11540
rect 8812 11500 8818 11512
rect 8849 11509 8861 11512
rect 8895 11509 8907 11543
rect 8849 11503 8907 11509
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 14246 11540 14274 11580
rect 15933 11577 15945 11611
rect 15979 11577 15991 11611
rect 18322 11608 18328 11620
rect 18235 11580 18328 11608
rect 15933 11571 15991 11577
rect 14369 11543 14427 11549
rect 14369 11540 14381 11543
rect 13872 11512 13917 11540
rect 14246 11512 14381 11540
rect 13872 11500 13878 11512
rect 14369 11509 14381 11512
rect 14415 11509 14427 11543
rect 14369 11503 14427 11509
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 15197 11543 15255 11549
rect 15197 11540 15209 11543
rect 14884 11512 15209 11540
rect 14884 11500 14890 11512
rect 15197 11509 15209 11512
rect 15243 11540 15255 11543
rect 15470 11540 15476 11552
rect 15243 11512 15476 11540
rect 15243 11509 15255 11512
rect 15197 11503 15255 11509
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 15948 11540 15976 11571
rect 18322 11568 18328 11580
rect 18380 11608 18386 11620
rect 19857 11617 19885 11648
rect 20438 11636 20444 11648
rect 20496 11636 20502 11688
rect 20806 11636 20812 11688
rect 20864 11676 20870 11688
rect 21821 11679 21879 11685
rect 21821 11676 21833 11679
rect 20864 11648 21833 11676
rect 20864 11636 20870 11648
rect 21821 11645 21833 11648
rect 21867 11645 21879 11679
rect 21821 11639 21879 11645
rect 19842 11611 19900 11617
rect 18380 11580 19472 11608
rect 18380 11568 18386 11580
rect 16206 11540 16212 11552
rect 15948 11512 16212 11540
rect 16206 11500 16212 11512
rect 16264 11540 16270 11552
rect 16761 11543 16819 11549
rect 16761 11540 16773 11543
rect 16264 11512 16773 11540
rect 16264 11500 16270 11512
rect 16761 11509 16773 11512
rect 16807 11509 16819 11543
rect 16761 11503 16819 11509
rect 17773 11543 17831 11549
rect 17773 11509 17785 11543
rect 17819 11540 17831 11543
rect 17862 11540 17868 11552
rect 17819 11512 17868 11540
rect 17819 11509 17831 11512
rect 17773 11503 17831 11509
rect 17862 11500 17868 11512
rect 17920 11540 17926 11552
rect 19334 11540 19340 11552
rect 17920 11512 19340 11540
rect 17920 11500 17926 11512
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 19444 11540 19472 11580
rect 19842 11577 19854 11611
rect 19888 11577 19900 11611
rect 19842 11571 19900 11577
rect 21358 11540 21364 11552
rect 19444 11512 21364 11540
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 21836 11540 21864 11639
rect 22094 11608 22100 11620
rect 22055 11580 22100 11608
rect 22094 11568 22100 11580
rect 22152 11568 22158 11620
rect 22189 11611 22247 11617
rect 22189 11577 22201 11611
rect 22235 11608 22247 11611
rect 22278 11608 22284 11620
rect 22235 11580 22284 11608
rect 22235 11577 22247 11580
rect 22189 11571 22247 11577
rect 22204 11540 22232 11571
rect 22278 11568 22284 11580
rect 22336 11568 22342 11620
rect 21836 11512 22232 11540
rect 22756 11540 22784 11716
rect 23477 11713 23489 11747
rect 23523 11744 23535 11747
rect 23753 11747 23811 11753
rect 23753 11744 23765 11747
rect 23523 11716 23765 11744
rect 23523 11713 23535 11716
rect 23477 11707 23535 11713
rect 23753 11713 23765 11716
rect 23799 11744 23811 11747
rect 25225 11747 25283 11753
rect 25225 11744 25237 11747
rect 23799 11716 25237 11744
rect 23799 11713 23811 11716
rect 23753 11707 23811 11713
rect 25225 11713 25237 11716
rect 25271 11713 25283 11747
rect 25225 11707 25283 11713
rect 23106 11568 23112 11620
rect 23164 11608 23170 11620
rect 23845 11611 23903 11617
rect 23845 11608 23857 11611
rect 23164 11580 23857 11608
rect 23164 11568 23170 11580
rect 23845 11577 23857 11580
rect 23891 11577 23903 11611
rect 23845 11571 23903 11577
rect 23474 11540 23480 11552
rect 22756 11512 23480 11540
rect 23474 11500 23480 11512
rect 23532 11500 23538 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 10042 11336 10048 11348
rect 10003 11308 10048 11336
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 10778 11336 10784 11348
rect 10739 11308 10784 11336
rect 10778 11296 10784 11308
rect 10836 11296 10842 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 12805 11339 12863 11345
rect 12805 11336 12817 11339
rect 12400 11308 12817 11336
rect 12400 11296 12406 11308
rect 12805 11305 12817 11308
rect 12851 11305 12863 11339
rect 16206 11336 16212 11348
rect 16167 11308 16212 11336
rect 12805 11299 12863 11305
rect 16206 11296 16212 11308
rect 16264 11296 16270 11348
rect 19334 11296 19340 11348
rect 19392 11336 19398 11348
rect 19429 11339 19487 11345
rect 19429 11336 19441 11339
rect 19392 11308 19441 11336
rect 19392 11296 19398 11308
rect 19429 11305 19441 11308
rect 19475 11305 19487 11339
rect 19429 11299 19487 11305
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 20349 11339 20407 11345
rect 20349 11336 20361 11339
rect 20036 11308 20361 11336
rect 20036 11296 20042 11308
rect 20349 11305 20361 11308
rect 20395 11336 20407 11339
rect 22554 11336 22560 11348
rect 20395 11308 21772 11336
rect 22515 11308 22560 11336
rect 20395 11305 20407 11308
rect 20349 11299 20407 11305
rect 11514 11268 11520 11280
rect 11475 11240 11520 11268
rect 11514 11228 11520 11240
rect 11572 11228 11578 11280
rect 12434 11228 12440 11280
rect 12492 11268 12498 11280
rect 12529 11271 12587 11277
rect 12529 11268 12541 11271
rect 12492 11240 12541 11268
rect 12492 11228 12498 11240
rect 12529 11237 12541 11240
rect 12575 11268 12587 11271
rect 12710 11268 12716 11280
rect 12575 11240 12716 11268
rect 12575 11237 12587 11240
rect 12529 11231 12587 11237
rect 12710 11228 12716 11240
rect 12768 11228 12774 11280
rect 13443 11271 13501 11277
rect 13443 11237 13455 11271
rect 13489 11268 13501 11271
rect 13538 11268 13544 11280
rect 13489 11240 13544 11268
rect 13489 11237 13501 11240
rect 13443 11231 13501 11237
rect 13538 11228 13544 11240
rect 13596 11228 13602 11280
rect 15470 11228 15476 11280
rect 15528 11268 15534 11280
rect 15610 11271 15668 11277
rect 15610 11268 15622 11271
rect 15528 11240 15622 11268
rect 15528 11228 15534 11240
rect 15610 11237 15622 11240
rect 15656 11237 15668 11271
rect 21174 11268 21180 11280
rect 21135 11240 21180 11268
rect 15610 11231 15668 11237
rect 21174 11228 21180 11240
rect 21232 11228 21238 11280
rect 21744 11277 21772 11308
rect 22554 11296 22560 11308
rect 22612 11296 22618 11348
rect 24118 11336 24124 11348
rect 24079 11308 24124 11336
rect 24118 11296 24124 11308
rect 24176 11296 24182 11348
rect 24394 11336 24400 11348
rect 24355 11308 24400 11336
rect 24394 11296 24400 11308
rect 24452 11296 24458 11348
rect 21729 11271 21787 11277
rect 21729 11237 21741 11271
rect 21775 11268 21787 11271
rect 21818 11268 21824 11280
rect 21775 11240 21824 11268
rect 21775 11237 21787 11240
rect 21729 11231 21787 11237
rect 21818 11228 21824 11240
rect 21876 11268 21882 11280
rect 22830 11268 22836 11280
rect 21876 11240 22836 11268
rect 21876 11228 21882 11240
rect 22830 11228 22836 11240
rect 22888 11228 22894 11280
rect 22934 11271 22992 11277
rect 22934 11237 22946 11271
rect 22980 11268 22992 11271
rect 23106 11268 23112 11280
rect 22980 11240 23112 11268
rect 22980 11237 22992 11240
rect 22934 11231 22992 11237
rect 23106 11228 23112 11240
rect 23164 11228 23170 11280
rect 23198 11228 23204 11280
rect 23256 11268 23262 11280
rect 23477 11271 23535 11277
rect 23477 11268 23489 11271
rect 23256 11240 23489 11268
rect 23256 11228 23262 11240
rect 23477 11237 23489 11240
rect 23523 11268 23535 11271
rect 24026 11268 24032 11280
rect 23523 11240 24032 11268
rect 23523 11237 23535 11240
rect 23477 11231 23535 11237
rect 24026 11228 24032 11240
rect 24084 11228 24090 11280
rect 7837 11203 7895 11209
rect 7837 11200 7849 11203
rect 7576 11172 7849 11200
rect 7282 10996 7288 11008
rect 7243 10968 7288 10996
rect 7282 10956 7288 10968
rect 7340 10956 7346 11008
rect 7466 10956 7472 11008
rect 7524 10996 7530 11008
rect 7576 11005 7604 11172
rect 7837 11169 7849 11172
rect 7883 11200 7895 11203
rect 8757 11203 8815 11209
rect 8757 11200 8769 11203
rect 7883 11172 8769 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 8757 11169 8769 11172
rect 8803 11169 8815 11203
rect 8757 11163 8815 11169
rect 8938 11160 8944 11212
rect 8996 11200 9002 11212
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 8996 11172 10057 11200
rect 8996 11160 9002 11172
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10318 11200 10324 11212
rect 10279 11172 10324 11200
rect 10045 11163 10103 11169
rect 7742 11132 7748 11144
rect 7703 11104 7748 11132
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 10060 11132 10088 11163
rect 10318 11160 10324 11172
rect 10376 11160 10382 11212
rect 12069 11203 12127 11209
rect 12069 11169 12081 11203
rect 12115 11200 12127 11203
rect 12115 11172 13629 11200
rect 12115 11169 12127 11172
rect 12069 11163 12127 11169
rect 11146 11132 11152 11144
rect 10060 11104 11152 11132
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11132 11483 11135
rect 11882 11132 11888 11144
rect 11471 11104 11888 11132
rect 11471 11101 11483 11104
rect 11425 11095 11483 11101
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 13078 11132 13084 11144
rect 13039 11104 13084 11132
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 13601 11132 13629 11172
rect 13722 11160 13728 11212
rect 13780 11200 13786 11212
rect 15286 11200 15292 11212
rect 13780 11172 15292 11200
rect 13780 11160 13786 11172
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 17494 11200 17500 11212
rect 17455 11172 17500 11200
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 17954 11200 17960 11212
rect 17915 11172 17960 11200
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 18506 11160 18512 11212
rect 18564 11200 18570 11212
rect 19061 11203 19119 11209
rect 19061 11200 19073 11203
rect 18564 11172 19073 11200
rect 18564 11160 18570 11172
rect 19061 11169 19073 11172
rect 19107 11200 19119 11203
rect 19242 11200 19248 11212
rect 19107 11172 19248 11200
rect 19107 11169 19119 11172
rect 19061 11163 19119 11169
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 24581 11203 24639 11209
rect 24581 11169 24593 11203
rect 24627 11200 24639 11203
rect 24670 11200 24676 11212
rect 24627 11172 24676 11200
rect 24627 11169 24639 11172
rect 24581 11163 24639 11169
rect 24670 11160 24676 11172
rect 24728 11160 24734 11212
rect 24857 11203 24915 11209
rect 24857 11169 24869 11203
rect 24903 11200 24915 11203
rect 25038 11200 25044 11212
rect 24903 11172 25044 11200
rect 24903 11169 24915 11172
rect 24857 11163 24915 11169
rect 25038 11160 25044 11172
rect 25096 11160 25102 11212
rect 15105 11135 15163 11141
rect 15105 11132 15117 11135
rect 13601 11104 15117 11132
rect 15105 11101 15117 11104
rect 15151 11132 15163 11135
rect 15378 11132 15384 11144
rect 15151 11104 15384 11132
rect 15151 11101 15163 11104
rect 15105 11095 15163 11101
rect 15378 11092 15384 11104
rect 15436 11132 15442 11144
rect 16022 11132 16028 11144
rect 15436 11104 16028 11132
rect 15436 11092 15442 11104
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 18230 11132 18236 11144
rect 18191 11104 18236 11132
rect 18230 11092 18236 11104
rect 18288 11092 18294 11144
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 21082 11132 21088 11144
rect 20772 11104 21088 11132
rect 20772 11092 20778 11104
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 22278 11092 22284 11144
rect 22336 11132 22342 11144
rect 22833 11135 22891 11141
rect 22833 11132 22845 11135
rect 22336 11104 22845 11132
rect 22336 11092 22342 11104
rect 22833 11101 22845 11104
rect 22879 11101 22891 11135
rect 22833 11095 22891 11101
rect 14001 11067 14059 11073
rect 14001 11064 14013 11067
rect 13786 11036 14013 11064
rect 7561 10999 7619 11005
rect 7561 10996 7573 10999
rect 7524 10968 7573 10996
rect 7524 10956 7530 10968
rect 7561 10965 7573 10968
rect 7607 10965 7619 10999
rect 7561 10959 7619 10965
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 9217 10999 9275 11005
rect 9217 10996 9229 10999
rect 9180 10968 9229 10996
rect 9180 10956 9186 10968
rect 9217 10965 9229 10968
rect 9263 10996 9275 10999
rect 9950 10996 9956 11008
rect 9263 10968 9956 10996
rect 9263 10965 9275 10968
rect 9217 10959 9275 10965
rect 9950 10956 9956 10968
rect 10008 10956 10014 11008
rect 10870 10956 10876 11008
rect 10928 10996 10934 11008
rect 11149 10999 11207 11005
rect 11149 10996 11161 10999
rect 10928 10968 11161 10996
rect 10928 10956 10934 10968
rect 11149 10965 11161 10968
rect 11195 10965 11207 10999
rect 11149 10959 11207 10965
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 13786 10996 13814 11036
rect 14001 11033 14013 11036
rect 14047 11064 14059 11067
rect 15838 11064 15844 11076
rect 14047 11036 15844 11064
rect 14047 11033 14059 11036
rect 14001 11027 14059 11033
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 14274 10996 14280 11008
rect 13412 10968 13814 10996
rect 14235 10968 14280 10996
rect 13412 10956 13418 10968
rect 14274 10956 14280 10968
rect 14332 10956 14338 11008
rect 15746 10956 15752 11008
rect 15804 10996 15810 11008
rect 16485 10999 16543 11005
rect 16485 10996 16497 10999
rect 15804 10968 16497 10996
rect 15804 10956 15810 10968
rect 16485 10965 16497 10968
rect 16531 10965 16543 10999
rect 19978 10996 19984 11008
rect 19939 10968 19984 10996
rect 16485 10959 16543 10965
rect 19978 10956 19984 10968
rect 20036 10956 20042 11008
rect 22094 10996 22100 11008
rect 22055 10968 22100 10996
rect 22094 10956 22100 10968
rect 22152 10956 22158 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 7009 10795 7067 10801
rect 7009 10792 7021 10795
rect 2832 10764 7021 10792
rect 2832 10752 2838 10764
rect 7009 10761 7021 10764
rect 7055 10761 7067 10795
rect 11514 10792 11520 10804
rect 11475 10764 11520 10792
rect 7009 10755 7067 10761
rect 7024 10588 7052 10755
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 12805 10795 12863 10801
rect 12805 10761 12817 10795
rect 12851 10792 12863 10795
rect 13538 10792 13544 10804
rect 12851 10764 13544 10792
rect 12851 10761 12863 10764
rect 12805 10755 12863 10761
rect 13538 10752 13544 10764
rect 13596 10792 13602 10804
rect 13725 10795 13783 10801
rect 13725 10792 13737 10795
rect 13596 10764 13737 10792
rect 13596 10752 13602 10764
rect 13725 10761 13737 10764
rect 13771 10761 13783 10795
rect 14826 10792 14832 10804
rect 14787 10764 14832 10792
rect 13725 10755 13783 10761
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 17221 10795 17279 10801
rect 17221 10761 17233 10795
rect 17267 10792 17279 10795
rect 17494 10792 17500 10804
rect 17267 10764 17500 10792
rect 17267 10761 17279 10764
rect 17221 10755 17279 10761
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 19978 10752 19984 10804
rect 20036 10792 20042 10804
rect 20625 10795 20683 10801
rect 20625 10792 20637 10795
rect 20036 10764 20637 10792
rect 20036 10752 20042 10764
rect 20625 10761 20637 10764
rect 20671 10792 20683 10795
rect 21174 10792 21180 10804
rect 20671 10764 21180 10792
rect 20671 10761 20683 10764
rect 20625 10755 20683 10761
rect 21174 10752 21180 10764
rect 21232 10752 21238 10804
rect 22186 10752 22192 10804
rect 22244 10792 22250 10804
rect 22741 10795 22799 10801
rect 22741 10792 22753 10795
rect 22244 10764 22753 10792
rect 22244 10752 22250 10764
rect 22741 10761 22753 10764
rect 22787 10792 22799 10795
rect 23106 10792 23112 10804
rect 22787 10764 23112 10792
rect 22787 10761 22799 10764
rect 22741 10755 22799 10761
rect 23106 10752 23112 10764
rect 23164 10752 23170 10804
rect 24670 10792 24676 10804
rect 24631 10764 24676 10792
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 25406 10792 25412 10804
rect 25367 10764 25412 10792
rect 25406 10752 25412 10764
rect 25464 10752 25470 10804
rect 8478 10684 8484 10736
rect 8536 10724 8542 10736
rect 8849 10727 8907 10733
rect 8849 10724 8861 10727
rect 8536 10696 8861 10724
rect 8536 10684 8542 10696
rect 8849 10693 8861 10696
rect 8895 10693 8907 10727
rect 21818 10724 21824 10736
rect 21779 10696 21824 10724
rect 8849 10687 8907 10693
rect 21818 10684 21824 10696
rect 21876 10684 21882 10736
rect 7745 10659 7803 10665
rect 7745 10625 7757 10659
rect 7791 10656 7803 10659
rect 8018 10656 8024 10668
rect 7791 10628 8024 10656
rect 7791 10625 7803 10628
rect 7745 10619 7803 10625
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 8113 10659 8171 10665
rect 8113 10625 8125 10659
rect 8159 10656 8171 10659
rect 8570 10656 8576 10668
rect 8159 10628 8576 10656
rect 8159 10625 8171 10628
rect 8113 10619 8171 10625
rect 8570 10616 8576 10628
rect 8628 10656 8634 10668
rect 8941 10659 8999 10665
rect 8941 10656 8953 10659
rect 8628 10628 8953 10656
rect 8628 10616 8634 10628
rect 8941 10625 8953 10628
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 9677 10659 9735 10665
rect 9677 10656 9689 10659
rect 9355 10628 9689 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 9677 10625 9689 10628
rect 9723 10656 9735 10659
rect 10045 10659 10103 10665
rect 10045 10656 10057 10659
rect 9723 10628 10057 10656
rect 9723 10625 9735 10628
rect 9677 10619 9735 10625
rect 10045 10625 10057 10628
rect 10091 10656 10103 10659
rect 10318 10656 10324 10668
rect 10091 10628 10324 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 10318 10616 10324 10628
rect 10376 10656 10382 10668
rect 10870 10656 10876 10668
rect 10376 10628 10732 10656
rect 10831 10628 10876 10656
rect 10376 10616 10382 10628
rect 7377 10591 7435 10597
rect 7377 10588 7389 10591
rect 7024 10560 7389 10588
rect 7377 10557 7389 10560
rect 7423 10588 7435 10591
rect 7466 10588 7472 10600
rect 7423 10560 7472 10588
rect 7423 10557 7435 10560
rect 7377 10551 7435 10557
rect 7466 10548 7472 10560
rect 7524 10588 7530 10600
rect 10704 10597 10732 10628
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 13035 10659 13093 10665
rect 13035 10625 13047 10659
rect 13081 10656 13093 10659
rect 13909 10659 13967 10665
rect 13081 10628 13814 10656
rect 13081 10625 13093 10628
rect 13035 10619 13093 10625
rect 8720 10591 8778 10597
rect 8720 10588 8732 10591
rect 7524 10560 8732 10588
rect 7524 10548 7530 10560
rect 8720 10557 8732 10560
rect 8766 10557 8778 10591
rect 8720 10551 8778 10557
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10557 10471 10591
rect 10413 10551 10471 10557
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10588 10747 10591
rect 12526 10588 12532 10600
rect 10735 10560 12532 10588
rect 10735 10557 10747 10560
rect 10689 10551 10747 10557
rect 7193 10523 7251 10529
rect 7193 10489 7205 10523
rect 7239 10520 7251 10523
rect 7282 10520 7288 10532
rect 7239 10492 7288 10520
rect 7239 10489 7251 10492
rect 7193 10483 7251 10489
rect 7282 10480 7288 10492
rect 7340 10520 7346 10532
rect 8202 10520 8208 10532
rect 7340 10492 8208 10520
rect 7340 10480 7346 10492
rect 8202 10480 8208 10492
rect 8260 10520 8266 10532
rect 8573 10523 8631 10529
rect 8573 10520 8585 10523
rect 8260 10492 8585 10520
rect 8260 10480 8266 10492
rect 8573 10489 8585 10492
rect 8619 10520 8631 10523
rect 9030 10520 9036 10532
rect 8619 10492 9036 10520
rect 8619 10489 8631 10492
rect 8573 10483 8631 10489
rect 9030 10480 9036 10492
rect 9088 10480 9094 10532
rect 10428 10520 10456 10551
rect 12526 10548 12532 10560
rect 12584 10548 12590 10600
rect 12948 10591 13006 10597
rect 12948 10557 12960 10591
rect 12994 10588 13006 10591
rect 13786 10588 13814 10628
rect 13909 10625 13921 10659
rect 13955 10656 13967 10659
rect 14274 10656 14280 10668
rect 13955 10628 14280 10656
rect 13955 10625 13967 10628
rect 13909 10619 13967 10625
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 15746 10656 15752 10668
rect 14384 10628 15752 10656
rect 14384 10588 14412 10628
rect 15746 10616 15752 10628
rect 15804 10616 15810 10668
rect 16022 10656 16028 10668
rect 15983 10628 16028 10656
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 18046 10656 18052 10668
rect 18007 10628 18052 10656
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 18138 10616 18144 10668
rect 18196 10656 18202 10668
rect 19429 10659 19487 10665
rect 19429 10656 19441 10659
rect 18196 10628 19441 10656
rect 18196 10616 18202 10628
rect 19429 10625 19441 10628
rect 19475 10656 19487 10659
rect 19978 10656 19984 10668
rect 19475 10628 19984 10656
rect 19475 10625 19487 10628
rect 19429 10619 19487 10625
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 20898 10616 20904 10668
rect 20956 10656 20962 10668
rect 22002 10656 22008 10668
rect 20956 10628 22008 10656
rect 20956 10616 20962 10628
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 24688 10656 24716 10752
rect 23952 10628 24716 10656
rect 12994 10560 13492 10588
rect 13786 10560 14412 10588
rect 20349 10591 20407 10597
rect 12994 10557 13006 10560
rect 12948 10551 13006 10557
rect 10778 10520 10784 10532
rect 10428 10492 10784 10520
rect 10778 10480 10784 10492
rect 10836 10520 10842 10532
rect 11330 10520 11336 10532
rect 10836 10492 11336 10520
rect 10836 10480 10842 10492
rect 11330 10480 11336 10492
rect 11388 10520 11394 10532
rect 12618 10520 12624 10532
rect 11388 10492 12624 10520
rect 11388 10480 11394 10492
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 13464 10464 13492 10560
rect 20349 10557 20361 10591
rect 20395 10588 20407 10591
rect 20993 10591 21051 10597
rect 20993 10588 21005 10591
rect 20395 10560 21005 10588
rect 20395 10557 20407 10560
rect 20349 10551 20407 10557
rect 20993 10557 21005 10560
rect 21039 10557 21051 10591
rect 20993 10551 21051 10557
rect 13538 10480 13544 10532
rect 13596 10520 13602 10532
rect 14231 10523 14289 10529
rect 13596 10492 13814 10520
rect 13596 10480 13602 10492
rect 8478 10452 8484 10464
rect 8439 10424 8484 10452
rect 8478 10412 8484 10424
rect 8536 10412 8542 10464
rect 11146 10452 11152 10464
rect 11107 10424 11152 10452
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11882 10452 11888 10464
rect 11843 10424 11888 10452
rect 11882 10412 11888 10424
rect 11940 10412 11946 10464
rect 13446 10452 13452 10464
rect 13407 10424 13452 10452
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 13786 10452 13814 10492
rect 14231 10489 14243 10523
rect 14277 10489 14289 10523
rect 15838 10520 15844 10532
rect 15751 10492 15844 10520
rect 14231 10483 14289 10489
rect 14246 10452 14274 10483
rect 15838 10480 15844 10492
rect 15896 10480 15902 10532
rect 19334 10520 19340 10532
rect 19076 10492 19340 10520
rect 15378 10452 15384 10464
rect 13786 10424 15384 10452
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 15856 10452 15884 10480
rect 16669 10455 16727 10461
rect 16669 10452 16681 10455
rect 15856 10424 16681 10452
rect 16669 10421 16681 10424
rect 16715 10421 16727 10455
rect 16669 10415 16727 10421
rect 17589 10455 17647 10461
rect 17589 10421 17601 10455
rect 17635 10452 17647 10455
rect 17954 10452 17960 10464
rect 17635 10424 17960 10452
rect 17635 10421 17647 10424
rect 17589 10415 17647 10421
rect 17954 10412 17960 10424
rect 18012 10452 18018 10464
rect 18138 10452 18144 10464
rect 18012 10424 18144 10452
rect 18012 10412 18018 10424
rect 18138 10412 18144 10424
rect 18196 10412 18202 10464
rect 18690 10452 18696 10464
rect 18651 10424 18696 10452
rect 18690 10412 18696 10424
rect 18748 10452 18754 10464
rect 19076 10461 19104 10492
rect 19334 10480 19340 10492
rect 19392 10520 19398 10532
rect 19750 10523 19808 10529
rect 19750 10520 19762 10523
rect 19392 10492 19762 10520
rect 19392 10480 19398 10492
rect 19750 10489 19762 10492
rect 19796 10489 19808 10523
rect 19750 10483 19808 10489
rect 19061 10455 19119 10461
rect 19061 10452 19073 10455
rect 18748 10424 19073 10452
rect 18748 10412 18754 10424
rect 19061 10421 19073 10424
rect 19107 10421 19119 10455
rect 21008 10452 21036 10551
rect 22370 10548 22376 10600
rect 22428 10588 22434 10600
rect 22738 10588 22744 10600
rect 22428 10560 22744 10588
rect 22428 10548 22434 10560
rect 22738 10548 22744 10560
rect 22796 10548 22802 10600
rect 23952 10597 23980 10628
rect 23937 10591 23995 10597
rect 23937 10588 23949 10591
rect 23400 10560 23949 10588
rect 21266 10520 21272 10532
rect 21227 10492 21272 10520
rect 21266 10480 21272 10492
rect 21324 10480 21330 10532
rect 21361 10523 21419 10529
rect 21361 10489 21373 10523
rect 21407 10489 21419 10523
rect 21361 10483 21419 10489
rect 21376 10452 21404 10483
rect 21008 10424 21404 10452
rect 19061 10415 19119 10421
rect 22278 10412 22284 10464
rect 22336 10452 22342 10464
rect 22373 10455 22431 10461
rect 22373 10452 22385 10455
rect 22336 10424 22385 10452
rect 22336 10412 22342 10424
rect 22373 10421 22385 10424
rect 22419 10421 22431 10455
rect 22373 10415 22431 10421
rect 23290 10412 23296 10464
rect 23348 10452 23354 10464
rect 23400 10461 23428 10560
rect 23937 10557 23949 10560
rect 23983 10557 23995 10591
rect 24118 10588 24124 10600
rect 24079 10560 24124 10588
rect 23937 10551 23995 10557
rect 24118 10548 24124 10560
rect 24176 10548 24182 10600
rect 25222 10588 25228 10600
rect 25183 10560 25228 10588
rect 25222 10548 25228 10560
rect 25280 10588 25286 10600
rect 25777 10591 25835 10597
rect 25777 10588 25789 10591
rect 25280 10560 25789 10588
rect 25280 10548 25286 10560
rect 25777 10557 25789 10560
rect 25823 10557 25835 10591
rect 25777 10551 25835 10557
rect 23385 10455 23443 10461
rect 23385 10452 23397 10455
rect 23348 10424 23397 10452
rect 23348 10412 23354 10424
rect 23385 10421 23397 10424
rect 23431 10421 23443 10455
rect 23750 10452 23756 10464
rect 23711 10424 23756 10452
rect 23385 10415 23443 10421
rect 23750 10412 23756 10424
rect 23808 10412 23814 10464
rect 25038 10452 25044 10464
rect 24999 10424 25044 10452
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 9309 10251 9367 10257
rect 9309 10248 9321 10251
rect 7800 10220 9321 10248
rect 7800 10208 7806 10220
rect 9309 10217 9321 10220
rect 9355 10248 9367 10251
rect 9401 10251 9459 10257
rect 9401 10248 9413 10251
rect 9355 10220 9413 10248
rect 9355 10217 9367 10220
rect 9309 10211 9367 10217
rect 9401 10217 9413 10220
rect 9447 10217 9459 10251
rect 9401 10211 9459 10217
rect 10321 10251 10379 10257
rect 10321 10217 10333 10251
rect 10367 10248 10379 10251
rect 12894 10248 12900 10260
rect 10367 10220 12900 10248
rect 10367 10217 10379 10220
rect 10321 10211 10379 10217
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 13078 10248 13084 10260
rect 13039 10220 13084 10248
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 15105 10251 15163 10257
rect 15105 10217 15117 10251
rect 15151 10248 15163 10251
rect 15286 10248 15292 10260
rect 15151 10220 15292 10248
rect 15151 10217 15163 10220
rect 15105 10211 15163 10217
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 18230 10208 18236 10260
rect 18288 10248 18294 10260
rect 18969 10251 19027 10257
rect 18969 10248 18981 10251
rect 18288 10220 18981 10248
rect 18288 10208 18294 10220
rect 18969 10217 18981 10220
rect 19015 10217 19027 10251
rect 18969 10211 19027 10217
rect 19242 10208 19248 10260
rect 19300 10248 19306 10260
rect 19337 10251 19395 10257
rect 19337 10248 19349 10251
rect 19300 10220 19349 10248
rect 19300 10208 19306 10220
rect 19337 10217 19349 10220
rect 19383 10217 19395 10251
rect 19978 10248 19984 10260
rect 19939 10220 19984 10248
rect 19337 10211 19395 10217
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 20714 10248 20720 10260
rect 20675 10220 20720 10248
rect 20714 10208 20720 10220
rect 20772 10208 20778 10260
rect 21266 10208 21272 10260
rect 21324 10248 21330 10260
rect 22005 10251 22063 10257
rect 22005 10248 22017 10251
rect 21324 10220 22017 10248
rect 21324 10208 21330 10220
rect 22005 10217 22017 10220
rect 22051 10248 22063 10251
rect 23198 10248 23204 10260
rect 22051 10220 23204 10248
rect 22051 10217 22063 10220
rect 22005 10211 22063 10217
rect 23198 10208 23204 10220
rect 23256 10208 23262 10260
rect 23753 10251 23811 10257
rect 23753 10248 23765 10251
rect 23446 10220 23765 10248
rect 5442 10180 5448 10192
rect 5403 10152 5448 10180
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 11882 10180 11888 10192
rect 7208 10152 11888 10180
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 1486 10112 1492 10124
rect 1443 10084 1492 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 1486 10072 1492 10084
rect 1544 10072 1550 10124
rect 3970 10072 3976 10124
rect 4028 10112 4034 10124
rect 4100 10115 4158 10121
rect 4100 10112 4112 10115
rect 4028 10084 4112 10112
rect 4028 10072 4034 10084
rect 4100 10081 4112 10084
rect 4146 10081 4158 10115
rect 4100 10075 4158 10081
rect 4203 10047 4261 10053
rect 4203 10013 4215 10047
rect 4249 10044 4261 10047
rect 5350 10044 5356 10056
rect 4249 10016 5356 10044
rect 4249 10013 4261 10016
rect 4203 10007 4261 10013
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 5994 10044 6000 10056
rect 5955 10016 6000 10044
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 7208 9976 7236 10152
rect 11882 10140 11888 10152
rect 11940 10140 11946 10192
rect 12805 10183 12863 10189
rect 12805 10149 12817 10183
rect 12851 10180 12863 10183
rect 14274 10180 14280 10192
rect 12851 10152 14280 10180
rect 12851 10149 12863 10152
rect 12805 10143 12863 10149
rect 14274 10140 14280 10152
rect 14332 10140 14338 10192
rect 15212 10152 16160 10180
rect 7742 10112 7748 10124
rect 7703 10084 7748 10112
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 7926 10112 7932 10124
rect 7887 10084 7932 10112
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10081 8355 10115
rect 8297 10075 8355 10081
rect 8312 10044 8340 10075
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9088 10084 9689 10112
rect 9088 10072 9094 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 10686 10112 10692 10124
rect 9677 10075 9735 10081
rect 9857 10084 10692 10112
rect 4126 9948 7236 9976
rect 7300 10016 8340 10044
rect 8757 10047 8815 10053
rect 1535 9911 1593 9917
rect 1535 9877 1547 9911
rect 1581 9908 1593 9911
rect 4126 9908 4154 9948
rect 1581 9880 4154 9908
rect 1581 9877 1593 9880
rect 1535 9871 1593 9877
rect 7098 9868 7104 9920
rect 7156 9908 7162 9920
rect 7300 9917 7328 10016
rect 8757 10013 8769 10047
rect 8803 10044 8815 10047
rect 8846 10044 8852 10056
rect 8803 10016 8852 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 8846 10004 8852 10016
rect 8904 10044 8910 10056
rect 9857 10044 9885 10084
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 12345 10115 12403 10121
rect 12345 10081 12357 10115
rect 12391 10081 12403 10115
rect 12526 10112 12532 10124
rect 12487 10084 12532 10112
rect 12345 10075 12403 10081
rect 10042 10044 10048 10056
rect 8904 10016 9885 10044
rect 10003 10016 10048 10044
rect 8904 10004 8910 10016
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 12066 10004 12072 10056
rect 12124 10044 12130 10056
rect 12360 10044 12388 10075
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 13630 10112 13636 10124
rect 13591 10084 13636 10112
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 13722 10072 13728 10124
rect 13780 10112 13786 10124
rect 14185 10115 14243 10121
rect 14185 10112 14197 10115
rect 13780 10084 14197 10112
rect 13780 10072 13786 10084
rect 14185 10081 14197 10084
rect 14231 10112 14243 10115
rect 15212 10112 15240 10152
rect 15930 10112 15936 10124
rect 14231 10084 15240 10112
rect 15891 10084 15936 10112
rect 14231 10081 14243 10084
rect 14185 10075 14243 10081
rect 15930 10072 15936 10084
rect 15988 10072 15994 10124
rect 16132 10121 16160 10152
rect 20990 10140 20996 10192
rect 21048 10180 21054 10192
rect 21085 10183 21143 10189
rect 21085 10180 21097 10183
rect 21048 10152 21097 10180
rect 21048 10140 21054 10152
rect 21085 10149 21097 10152
rect 21131 10149 21143 10183
rect 23290 10180 23296 10192
rect 21085 10143 21143 10149
rect 22756 10152 23296 10180
rect 16117 10115 16175 10121
rect 16117 10081 16129 10115
rect 16163 10112 16175 10115
rect 16574 10112 16580 10124
rect 16163 10084 16580 10112
rect 16163 10081 16175 10084
rect 16117 10075 16175 10081
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 17494 10072 17500 10124
rect 17552 10112 17558 10124
rect 17957 10115 18015 10121
rect 17957 10112 17969 10115
rect 17552 10084 17969 10112
rect 17552 10072 17558 10084
rect 17957 10081 17969 10084
rect 18003 10081 18015 10115
rect 17957 10075 18015 10081
rect 18138 10072 18144 10124
rect 18196 10112 18202 10124
rect 18417 10115 18475 10121
rect 18417 10112 18429 10115
rect 18196 10084 18429 10112
rect 18196 10072 18202 10084
rect 18417 10081 18429 10084
rect 18463 10081 18475 10115
rect 18417 10075 18475 10081
rect 19150 10072 19156 10124
rect 19208 10112 19214 10124
rect 22756 10121 22784 10152
rect 23290 10140 23296 10152
rect 23348 10140 23354 10192
rect 19521 10115 19579 10121
rect 19521 10112 19533 10115
rect 19208 10084 19533 10112
rect 19208 10072 19214 10084
rect 19521 10081 19533 10084
rect 19567 10081 19579 10115
rect 19521 10075 19579 10081
rect 22741 10115 22799 10121
rect 22741 10081 22753 10115
rect 22787 10081 22799 10115
rect 22922 10112 22928 10124
rect 22883 10084 22928 10112
rect 22741 10075 22799 10081
rect 22922 10072 22928 10084
rect 22980 10072 22986 10124
rect 13648 10044 13676 10072
rect 14090 10044 14096 10056
rect 12124 10016 14096 10044
rect 12124 10004 12130 10016
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 14366 10044 14372 10056
rect 14327 10016 14372 10044
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 16206 10044 16212 10056
rect 16167 10016 16212 10044
rect 16206 10004 16212 10016
rect 16264 10004 16270 10056
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10044 18751 10047
rect 19426 10044 19432 10056
rect 18739 10016 19432 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 20806 10004 20812 10056
rect 20864 10044 20870 10056
rect 20993 10047 21051 10053
rect 20993 10044 21005 10047
rect 20864 10016 21005 10044
rect 20864 10004 20870 10016
rect 20993 10013 21005 10016
rect 21039 10013 21051 10047
rect 23017 10047 23075 10053
rect 23017 10044 23029 10047
rect 20993 10007 21051 10013
rect 21100 10016 23029 10044
rect 8938 9936 8944 9988
rect 8996 9976 9002 9988
rect 11885 9979 11943 9985
rect 11885 9976 11897 9979
rect 8996 9948 11897 9976
rect 8996 9936 9002 9948
rect 11885 9945 11897 9948
rect 11931 9976 11943 9979
rect 12526 9976 12532 9988
rect 11931 9948 12532 9976
rect 11931 9945 11943 9948
rect 11885 9939 11943 9945
rect 12526 9936 12532 9948
rect 12584 9936 12590 9988
rect 20254 9936 20260 9988
rect 20312 9976 20318 9988
rect 21100 9976 21128 10016
rect 23017 10013 23029 10016
rect 23063 10013 23075 10047
rect 23017 10007 23075 10013
rect 21542 9976 21548 9988
rect 20312 9948 21128 9976
rect 21503 9948 21548 9976
rect 20312 9936 20318 9948
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 23446 9920 23474 10220
rect 23753 10217 23765 10220
rect 23799 10248 23811 10251
rect 24118 10248 24124 10260
rect 23799 10220 24124 10248
rect 23799 10217 23811 10220
rect 23753 10211 23811 10217
rect 24118 10208 24124 10220
rect 24176 10208 24182 10260
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 7156 9880 7297 9908
rect 7156 9868 7162 9880
rect 7285 9877 7297 9880
rect 7331 9877 7343 9911
rect 9030 9908 9036 9920
rect 8991 9880 9036 9908
rect 7285 9871 7343 9877
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 9306 9908 9312 9920
rect 9219 9880 9312 9908
rect 9306 9868 9312 9880
rect 9364 9908 9370 9920
rect 9815 9911 9873 9917
rect 9815 9908 9827 9911
rect 9364 9880 9827 9908
rect 9364 9868 9370 9880
rect 9815 9877 9827 9880
rect 9861 9877 9873 9911
rect 9950 9908 9956 9920
rect 9911 9880 9956 9908
rect 9815 9871 9873 9877
rect 9950 9868 9956 9880
rect 10008 9868 10014 9920
rect 10594 9868 10600 9920
rect 10652 9908 10658 9920
rect 10689 9911 10747 9917
rect 10689 9908 10701 9911
rect 10652 9880 10701 9908
rect 10652 9868 10658 9880
rect 10689 9877 10701 9880
rect 10735 9877 10747 9911
rect 11054 9908 11060 9920
rect 11015 9880 11060 9908
rect 10689 9871 10747 9877
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 15562 9908 15568 9920
rect 15523 9880 15568 9908
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 16850 9868 16856 9920
rect 16908 9908 16914 9920
rect 23198 9908 23204 9920
rect 16908 9880 23204 9908
rect 16908 9868 16914 9880
rect 23198 9868 23204 9880
rect 23256 9868 23262 9920
rect 23382 9868 23388 9920
rect 23440 9880 23474 9920
rect 23440 9868 23446 9880
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 3970 9704 3976 9716
rect 3931 9676 3976 9704
rect 3970 9664 3976 9676
rect 4028 9664 4034 9716
rect 5350 9664 5356 9716
rect 5408 9704 5414 9716
rect 6549 9707 6607 9713
rect 6549 9704 6561 9707
rect 5408 9676 6561 9704
rect 5408 9664 5414 9676
rect 6549 9673 6561 9676
rect 6595 9673 6607 9707
rect 7558 9704 7564 9716
rect 7519 9676 7564 9704
rect 6549 9667 6607 9673
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 7926 9664 7932 9716
rect 7984 9704 7990 9716
rect 8297 9707 8355 9713
rect 8297 9704 8309 9707
rect 7984 9676 8309 9704
rect 7984 9664 7990 9676
rect 8297 9673 8309 9676
rect 8343 9673 8355 9707
rect 9674 9704 9680 9716
rect 9635 9676 9680 9704
rect 8297 9667 8355 9673
rect 9674 9664 9680 9676
rect 9732 9664 9738 9716
rect 12161 9707 12219 9713
rect 12161 9673 12173 9707
rect 12207 9704 12219 9707
rect 12434 9704 12440 9716
rect 12207 9676 12440 9704
rect 12207 9673 12219 9676
rect 12161 9667 12219 9673
rect 12434 9664 12440 9676
rect 12492 9664 12498 9716
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 12676 9676 15332 9704
rect 12676 9664 12682 9676
rect 4295 9639 4353 9645
rect 4295 9605 4307 9639
rect 4341 9636 4353 9639
rect 8938 9636 8944 9648
rect 4341 9608 8944 9636
rect 4341 9605 4353 9608
rect 4295 9599 4353 9605
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 9309 9639 9367 9645
rect 9309 9605 9321 9639
rect 9355 9636 9367 9639
rect 9582 9636 9588 9648
rect 9355 9608 9588 9636
rect 9355 9605 9367 9608
rect 9309 9599 9367 9605
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 10594 9636 10600 9648
rect 9876 9608 10600 9636
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 5261 9571 5319 9577
rect 5261 9568 5273 9571
rect 4120 9540 5273 9568
rect 4120 9528 4126 9540
rect 5261 9537 5273 9540
rect 5307 9568 5319 9571
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 5307 9540 6193 9568
rect 5307 9537 5319 9540
rect 5261 9531 5319 9537
rect 6181 9537 6193 9540
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 9398 9568 9404 9580
rect 8260 9540 9404 9568
rect 8260 9528 8266 9540
rect 9398 9528 9404 9540
rect 9456 9568 9462 9580
rect 9876 9568 9904 9608
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 15304 9636 15332 9676
rect 15562 9664 15568 9716
rect 15620 9704 15626 9716
rect 20257 9707 20315 9713
rect 20257 9704 20269 9707
rect 15620 9676 20269 9704
rect 15620 9664 15626 9676
rect 20257 9673 20269 9676
rect 20303 9704 20315 9707
rect 20625 9707 20683 9713
rect 20625 9704 20637 9707
rect 20303 9676 20637 9704
rect 20303 9673 20315 9676
rect 20257 9667 20315 9673
rect 20625 9673 20637 9676
rect 20671 9704 20683 9707
rect 20990 9704 20996 9716
rect 20671 9676 20996 9704
rect 20671 9673 20683 9676
rect 20625 9667 20683 9673
rect 20990 9664 20996 9676
rect 21048 9664 21054 9716
rect 22094 9664 22100 9716
rect 22152 9704 22158 9716
rect 22511 9707 22569 9713
rect 22511 9704 22523 9707
rect 22152 9676 22523 9704
rect 22152 9664 22158 9676
rect 22511 9673 22523 9676
rect 22557 9673 22569 9707
rect 23290 9704 23296 9716
rect 23251 9676 23296 9704
rect 22511 9667 22569 9673
rect 23290 9664 23296 9676
rect 23348 9664 23354 9716
rect 15381 9639 15439 9645
rect 15381 9636 15393 9639
rect 15304 9608 15393 9636
rect 15381 9605 15393 9608
rect 15427 9636 15439 9639
rect 15930 9636 15936 9648
rect 15427 9608 15936 9636
rect 15427 9605 15439 9608
rect 15381 9599 15439 9605
rect 15930 9596 15936 9608
rect 15988 9596 15994 9648
rect 19245 9639 19303 9645
rect 19245 9605 19257 9639
rect 19291 9636 19303 9639
rect 21266 9636 21272 9648
rect 19291 9608 21272 9636
rect 19291 9605 19303 9608
rect 19245 9599 19303 9605
rect 21266 9596 21272 9608
rect 21324 9596 21330 9648
rect 22186 9636 22192 9648
rect 22147 9608 22192 9636
rect 22186 9596 22192 9608
rect 22244 9636 22250 9648
rect 22922 9636 22928 9648
rect 22244 9608 22928 9636
rect 22244 9596 22250 9608
rect 22922 9596 22928 9608
rect 22980 9596 22986 9648
rect 9456 9540 9904 9568
rect 9456 9528 9462 9540
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 10008 9540 10793 9568
rect 10008 9528 10014 9540
rect 10781 9537 10793 9540
rect 10827 9568 10839 9571
rect 11054 9568 11060 9580
rect 10827 9540 11060 9568
rect 10827 9537 10839 9540
rect 10781 9531 10839 9537
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 11422 9568 11428 9580
rect 11383 9540 11428 9568
rect 11422 9528 11428 9540
rect 11480 9528 11486 9580
rect 12526 9568 12532 9580
rect 12487 9540 12532 9568
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9568 15071 9571
rect 15565 9571 15623 9577
rect 15565 9568 15577 9571
rect 15059 9540 15577 9568
rect 15059 9537 15071 9540
rect 15013 9531 15071 9537
rect 15565 9537 15577 9540
rect 15611 9568 15623 9571
rect 15746 9568 15752 9580
rect 15611 9540 15752 9568
rect 15611 9537 15623 9540
rect 15565 9531 15623 9537
rect 15746 9528 15752 9540
rect 15804 9528 15810 9580
rect 16022 9568 16028 9580
rect 15983 9540 16028 9568
rect 16022 9528 16028 9540
rect 16080 9528 16086 9580
rect 18230 9528 18236 9580
rect 18288 9568 18294 9580
rect 18325 9571 18383 9577
rect 18325 9568 18337 9571
rect 18288 9540 18337 9568
rect 18288 9528 18294 9540
rect 18325 9537 18337 9540
rect 18371 9537 18383 9571
rect 18325 9531 18383 9537
rect 19981 9571 20039 9577
rect 19981 9537 19993 9571
rect 20027 9568 20039 9571
rect 20898 9568 20904 9580
rect 20027 9540 20904 9568
rect 20027 9537 20039 9540
rect 19981 9531 20039 9537
rect 20898 9528 20904 9540
rect 20956 9528 20962 9580
rect 21174 9568 21180 9580
rect 21135 9540 21180 9568
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 4246 9509 4252 9512
rect 4224 9503 4252 9509
rect 4224 9500 4236 9503
rect 4159 9472 4236 9500
rect 4224 9469 4236 9472
rect 4304 9500 4310 9512
rect 4617 9503 4675 9509
rect 4617 9500 4629 9503
rect 4304 9472 4629 9500
rect 4224 9463 4252 9469
rect 4246 9460 4252 9463
rect 4304 9460 4310 9472
rect 4617 9469 4629 9472
rect 4663 9469 4675 9503
rect 7377 9503 7435 9509
rect 7377 9500 7389 9503
rect 4617 9463 4675 9469
rect 7116 9472 7389 9500
rect 5077 9435 5135 9441
rect 5077 9401 5089 9435
rect 5123 9432 5135 9435
rect 5350 9432 5356 9444
rect 5123 9404 5356 9432
rect 5123 9401 5135 9404
rect 5077 9395 5135 9401
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 5905 9435 5963 9441
rect 5905 9401 5917 9435
rect 5951 9432 5963 9435
rect 6270 9432 6276 9444
rect 5951 9404 6276 9432
rect 5951 9401 5963 9404
rect 5905 9395 5963 9401
rect 6270 9392 6276 9404
rect 6328 9392 6334 9444
rect 7116 9376 7144 9472
rect 7377 9469 7389 9472
rect 7423 9469 7435 9503
rect 7377 9463 7435 9469
rect 9180 9503 9238 9509
rect 9180 9469 9192 9503
rect 9226 9500 9238 9503
rect 9306 9500 9312 9512
rect 9226 9472 9312 9500
rect 9226 9469 9238 9472
rect 9180 9463 9238 9469
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 10686 9500 10692 9512
rect 10647 9472 10692 9500
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 10962 9500 10968 9512
rect 10923 9472 10968 9500
rect 10962 9460 10968 9472
rect 11020 9460 11026 9512
rect 13998 9500 14004 9512
rect 13959 9472 14004 9500
rect 13998 9460 14004 9472
rect 14056 9500 14062 9512
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 14056 9472 14565 9500
rect 14056 9460 14062 9472
rect 14553 9469 14565 9472
rect 14599 9469 14611 9503
rect 14553 9463 14611 9469
rect 22094 9460 22100 9512
rect 22152 9500 22158 9512
rect 22408 9503 22466 9509
rect 22408 9500 22420 9503
rect 22152 9472 22420 9500
rect 22152 9460 22158 9472
rect 22408 9469 22420 9472
rect 22454 9500 22466 9503
rect 22833 9503 22891 9509
rect 22833 9500 22845 9503
rect 22454 9472 22845 9500
rect 22454 9469 22466 9472
rect 22408 9463 22466 9469
rect 22833 9469 22845 9472
rect 22879 9500 22891 9503
rect 25222 9500 25228 9512
rect 22879 9472 25228 9500
rect 22879 9469 22891 9472
rect 22833 9463 22891 9469
rect 25222 9460 25228 9472
rect 25280 9460 25286 9512
rect 9030 9432 9036 9444
rect 8991 9404 9036 9432
rect 9030 9392 9036 9404
rect 9088 9392 9094 9444
rect 10704 9432 10732 9460
rect 11701 9435 11759 9441
rect 11701 9432 11713 9435
rect 10704 9404 11713 9432
rect 11701 9401 11713 9404
rect 11747 9401 11759 9435
rect 11701 9395 11759 9401
rect 12621 9435 12679 9441
rect 12621 9401 12633 9435
rect 12667 9432 12679 9435
rect 12802 9432 12808 9444
rect 12667 9404 12808 9432
rect 12667 9401 12679 9404
rect 12621 9395 12679 9401
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 13173 9435 13231 9441
rect 13173 9401 13185 9435
rect 13219 9432 13231 9435
rect 13354 9432 13360 9444
rect 13219 9404 13360 9432
rect 13219 9401 13231 9404
rect 13173 9395 13231 9401
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 15562 9392 15568 9444
rect 15620 9432 15626 9444
rect 15657 9435 15715 9441
rect 15657 9432 15669 9435
rect 15620 9404 15669 9432
rect 15620 9392 15626 9404
rect 15657 9401 15669 9404
rect 15703 9401 15715 9435
rect 16574 9432 16580 9444
rect 16487 9404 16580 9432
rect 15657 9395 15715 9401
rect 16574 9392 16580 9404
rect 16632 9432 16638 9444
rect 18138 9432 18144 9444
rect 16632 9404 18144 9432
rect 16632 9392 16638 9404
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 20990 9392 20996 9444
rect 21048 9432 21054 9444
rect 21048 9404 21093 9432
rect 21048 9392 21054 9404
rect 1486 9324 1492 9376
rect 1544 9364 1550 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 1544 9336 1593 9364
rect 1544 9324 1550 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 7098 9364 7104 9376
rect 7059 9336 7104 9364
rect 1581 9327 1639 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 8478 9324 8484 9376
rect 8536 9364 8542 9376
rect 8941 9367 8999 9373
rect 8941 9364 8953 9367
rect 8536 9336 8953 9364
rect 8536 9324 8542 9336
rect 8941 9333 8953 9336
rect 8987 9364 8999 9367
rect 9582 9364 9588 9376
rect 8987 9336 9588 9364
rect 8987 9333 8999 9336
rect 8941 9327 8999 9333
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 10042 9364 10048 9376
rect 10003 9336 10048 9364
rect 10042 9324 10048 9336
rect 10100 9364 10106 9376
rect 10505 9367 10563 9373
rect 10505 9364 10517 9367
rect 10100 9336 10517 9364
rect 10100 9324 10106 9336
rect 10505 9333 10517 9336
rect 10551 9364 10563 9367
rect 10962 9364 10968 9376
rect 10551 9336 10968 9364
rect 10551 9333 10563 9336
rect 10505 9327 10563 9333
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 13633 9367 13691 9373
rect 13633 9364 13645 9367
rect 12952 9336 13645 9364
rect 12952 9324 12958 9336
rect 13633 9333 13645 9336
rect 13679 9364 13691 9367
rect 13722 9364 13728 9376
rect 13679 9336 13728 9364
rect 13679 9333 13691 9336
rect 13633 9327 13691 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 14182 9364 14188 9376
rect 14143 9336 14188 9364
rect 14182 9324 14188 9336
rect 14240 9324 14246 9376
rect 17494 9364 17500 9376
rect 17455 9336 17500 9364
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17770 9364 17776 9376
rect 17731 9336 17776 9364
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 18690 9324 18696 9376
rect 18748 9364 18754 9376
rect 18748 9336 18793 9364
rect 18748 9324 18754 9336
rect 20806 9324 20812 9376
rect 20864 9364 20870 9376
rect 21821 9367 21879 9373
rect 21821 9364 21833 9367
rect 20864 9336 21833 9364
rect 20864 9324 20870 9336
rect 21821 9333 21833 9336
rect 21867 9333 21879 9367
rect 21821 9327 21879 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 7193 9163 7251 9169
rect 7193 9129 7205 9163
rect 7239 9160 7251 9163
rect 7742 9160 7748 9172
rect 7239 9132 7748 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 11054 9160 11060 9172
rect 11015 9132 11060 9160
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11606 9120 11612 9172
rect 11664 9160 11670 9172
rect 12066 9160 12072 9172
rect 11664 9132 12072 9160
rect 11664 9120 11670 9132
rect 12066 9120 12072 9132
rect 12124 9160 12130 9172
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 12124 9132 12357 9160
rect 12124 9120 12130 9132
rect 12345 9129 12357 9132
rect 12391 9129 12403 9163
rect 12345 9123 12403 9129
rect 13630 9120 13636 9172
rect 13688 9160 13694 9172
rect 13814 9160 13820 9172
rect 13688 9132 13820 9160
rect 13688 9120 13694 9132
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 17175 9163 17233 9169
rect 17175 9160 17187 9163
rect 15804 9132 17187 9160
rect 15804 9120 15810 9132
rect 17175 9129 17187 9132
rect 17221 9129 17233 9163
rect 17175 9123 17233 9129
rect 19426 9120 19432 9172
rect 19484 9160 19490 9172
rect 19981 9163 20039 9169
rect 19981 9160 19993 9163
rect 19484 9132 19993 9160
rect 19484 9120 19490 9132
rect 19981 9129 19993 9132
rect 20027 9129 20039 9163
rect 19981 9123 20039 9129
rect 5899 9095 5957 9101
rect 5899 9061 5911 9095
rect 5945 9092 5957 9095
rect 6178 9092 6184 9104
rect 5945 9064 6184 9092
rect 5945 9061 5957 9064
rect 5899 9055 5957 9061
rect 6178 9052 6184 9064
rect 6236 9052 6242 9104
rect 10413 9095 10471 9101
rect 10413 9061 10425 9095
rect 10459 9092 10471 9095
rect 12894 9092 12900 9104
rect 10459 9064 12900 9092
rect 10459 9061 10471 9064
rect 10413 9055 10471 9061
rect 12894 9052 12900 9064
rect 12952 9052 12958 9104
rect 13170 9092 13176 9104
rect 13131 9064 13176 9092
rect 13170 9052 13176 9064
rect 13228 9052 13234 9104
rect 15378 9052 15384 9104
rect 15436 9092 15442 9104
rect 15651 9095 15709 9101
rect 15651 9092 15663 9095
rect 15436 9064 15663 9092
rect 15436 9052 15442 9064
rect 15651 9061 15663 9064
rect 15697 9092 15709 9095
rect 15838 9092 15844 9104
rect 15697 9064 15844 9092
rect 15697 9061 15709 9064
rect 15651 9055 15709 9061
rect 15838 9052 15844 9064
rect 15896 9052 15902 9104
rect 18779 9095 18837 9101
rect 18779 9061 18791 9095
rect 18825 9092 18837 9095
rect 19610 9092 19616 9104
rect 18825 9064 19616 9092
rect 18825 9061 18837 9064
rect 18779 9055 18837 9061
rect 19610 9052 19616 9064
rect 19668 9052 19674 9104
rect 20622 9052 20628 9104
rect 20680 9092 20686 9104
rect 21085 9095 21143 9101
rect 21085 9092 21097 9095
rect 20680 9064 21097 9092
rect 20680 9052 20686 9064
rect 21085 9061 21097 9064
rect 21131 9061 21143 9095
rect 21085 9055 21143 9061
rect 7466 9024 7472 9036
rect 7427 8996 7472 9024
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 9030 8984 9036 9036
rect 9088 9024 9094 9036
rect 9125 9027 9183 9033
rect 9125 9024 9137 9027
rect 9088 8996 9137 9024
rect 9088 8984 9094 8996
rect 9125 8993 9137 8996
rect 9171 9024 9183 9027
rect 9490 9024 9496 9036
rect 9171 8996 9496 9024
rect 9171 8993 9183 8996
rect 9125 8987 9183 8993
rect 9490 8984 9496 8996
rect 9548 9024 9554 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 9548 8996 9689 9024
rect 9548 8984 9554 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 10134 9024 10140 9036
rect 9677 8987 9735 8993
rect 9857 8996 10140 9024
rect 4522 8956 4528 8968
rect 4483 8928 4528 8956
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 5534 8956 5540 8968
rect 5495 8928 5540 8956
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 7282 8956 7288 8968
rect 7243 8928 7288 8956
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 9306 8916 9312 8968
rect 9364 8956 9370 8968
rect 9857 8965 9885 8996
rect 10134 8984 10140 8996
rect 10192 9024 10198 9036
rect 10689 9027 10747 9033
rect 10689 9024 10701 9027
rect 10192 8996 10701 9024
rect 10192 8984 10198 8996
rect 10689 8993 10701 8996
rect 10735 8993 10747 9027
rect 11606 9024 11612 9036
rect 11567 8996 11612 9024
rect 10689 8987 10747 8993
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 11790 9024 11796 9036
rect 11751 8996 11796 9024
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 14366 8984 14372 9036
rect 14424 9024 14430 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 14424 8996 15301 9024
rect 14424 8984 14430 8996
rect 15289 8993 15301 8996
rect 15335 9024 15347 9027
rect 15470 9024 15476 9036
rect 15335 8996 15476 9024
rect 15335 8993 15347 8996
rect 15289 8987 15347 8993
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 17034 9024 17040 9036
rect 16995 8996 17040 9024
rect 17034 8984 17040 8996
rect 17092 8984 17098 9036
rect 9824 8959 9885 8965
rect 9824 8956 9836 8959
rect 9364 8928 9836 8956
rect 9364 8916 9370 8928
rect 9824 8925 9836 8928
rect 9870 8928 9885 8959
rect 10042 8956 10048 8968
rect 10003 8928 10048 8956
rect 9870 8925 9882 8928
rect 9824 8919 9882 8925
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 12066 8956 12072 8968
rect 12027 8928 12072 8956
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 13078 8956 13084 8968
rect 13039 8928 13084 8956
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 13354 8956 13360 8968
rect 13315 8928 13360 8956
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 18417 8959 18475 8965
rect 18417 8925 18429 8959
rect 18463 8956 18475 8959
rect 18598 8956 18604 8968
rect 18463 8928 18604 8956
rect 18463 8925 18475 8928
rect 18417 8919 18475 8925
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 20990 8956 20996 8968
rect 20903 8928 20996 8956
rect 20990 8916 20996 8928
rect 21048 8956 21054 8968
rect 22465 8959 22523 8965
rect 22465 8956 22477 8959
rect 21048 8928 22477 8956
rect 21048 8916 21054 8928
rect 22465 8925 22477 8928
rect 22511 8925 22523 8959
rect 22465 8919 22523 8925
rect 5261 8891 5319 8897
rect 5261 8857 5273 8891
rect 5307 8888 5319 8891
rect 5350 8888 5356 8900
rect 5307 8860 5356 8888
rect 5307 8857 5319 8860
rect 5261 8851 5319 8857
rect 5350 8848 5356 8860
rect 5408 8888 5414 8900
rect 6457 8891 6515 8897
rect 6457 8888 6469 8891
rect 5408 8860 6469 8888
rect 5408 8848 5414 8860
rect 6457 8857 6469 8860
rect 6503 8888 6515 8891
rect 7466 8888 7472 8900
rect 6503 8860 7472 8888
rect 6503 8857 6515 8860
rect 6457 8851 6515 8857
rect 7466 8848 7472 8860
rect 7524 8848 7530 8900
rect 13372 8888 13400 8916
rect 13906 8888 13912 8900
rect 13372 8860 13912 8888
rect 13906 8848 13912 8860
rect 13964 8848 13970 8900
rect 14090 8888 14096 8900
rect 14003 8860 14096 8888
rect 14090 8848 14096 8860
rect 14148 8888 14154 8900
rect 14148 8860 19748 8888
rect 14148 8848 14154 8860
rect 6825 8823 6883 8829
rect 6825 8789 6837 8823
rect 6871 8820 6883 8823
rect 6914 8820 6920 8832
rect 6871 8792 6920 8820
rect 6871 8789 6883 8792
rect 6825 8783 6883 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 8570 8820 8576 8832
rect 8531 8792 8576 8820
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 9490 8820 9496 8832
rect 9451 8792 9496 8820
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 9953 8823 10011 8829
rect 9953 8820 9965 8823
rect 9640 8792 9965 8820
rect 9640 8780 9646 8792
rect 9953 8789 9965 8792
rect 9999 8820 10011 8823
rect 10778 8820 10784 8832
rect 9999 8792 10784 8820
rect 9999 8789 10011 8792
rect 9953 8783 10011 8789
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 12802 8820 12808 8832
rect 12763 8792 12808 8820
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 16209 8823 16267 8829
rect 16209 8789 16221 8823
rect 16255 8820 16267 8823
rect 16298 8820 16304 8832
rect 16255 8792 16304 8820
rect 16255 8789 16267 8792
rect 16209 8783 16267 8789
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 18049 8823 18107 8829
rect 18049 8789 18061 8823
rect 18095 8820 18107 8823
rect 18138 8820 18144 8832
rect 18095 8792 18144 8820
rect 18095 8789 18107 8792
rect 18049 8783 18107 8789
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 19334 8820 19340 8832
rect 19295 8792 19340 8820
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 19610 8820 19616 8832
rect 19571 8792 19616 8820
rect 19610 8780 19616 8792
rect 19668 8780 19674 8832
rect 19720 8820 19748 8860
rect 21174 8848 21180 8900
rect 21232 8888 21238 8900
rect 21545 8891 21603 8897
rect 21545 8888 21557 8891
rect 21232 8860 21557 8888
rect 21232 8848 21238 8860
rect 21545 8857 21557 8860
rect 21591 8888 21603 8891
rect 21913 8891 21971 8897
rect 21913 8888 21925 8891
rect 21591 8860 21925 8888
rect 21591 8857 21603 8860
rect 21545 8851 21603 8857
rect 21913 8857 21925 8860
rect 21959 8857 21971 8891
rect 21913 8851 21971 8857
rect 23382 8820 23388 8832
rect 19720 8792 23388 8820
rect 23382 8780 23388 8792
rect 23440 8780 23446 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 8018 8616 8024 8628
rect 7979 8588 8024 8616
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 10689 8619 10747 8625
rect 10689 8616 10701 8619
rect 9548 8588 10701 8616
rect 9548 8576 9554 8588
rect 10689 8585 10701 8588
rect 10735 8585 10747 8619
rect 10689 8579 10747 8585
rect 11241 8619 11299 8625
rect 11241 8585 11253 8619
rect 11287 8616 11299 8619
rect 11606 8616 11612 8628
rect 11287 8588 11612 8616
rect 11287 8585 11299 8588
rect 11241 8579 11299 8585
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 12802 8576 12808 8628
rect 12860 8616 12866 8628
rect 13357 8619 13415 8625
rect 13357 8616 13369 8619
rect 12860 8588 13369 8616
rect 12860 8576 12866 8588
rect 13357 8585 13369 8588
rect 13403 8585 13415 8619
rect 13357 8579 13415 8585
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 15841 8619 15899 8625
rect 15841 8616 15853 8619
rect 15620 8588 15853 8616
rect 15620 8576 15626 8588
rect 15841 8585 15853 8588
rect 15887 8585 15899 8619
rect 15841 8579 15899 8585
rect 18463 8619 18521 8625
rect 18463 8585 18475 8619
rect 18509 8616 18521 8619
rect 20806 8616 20812 8628
rect 18509 8588 20812 8616
rect 18509 8585 18521 8588
rect 18463 8579 18521 8585
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 20990 8616 20996 8628
rect 20951 8588 20996 8616
rect 20990 8576 20996 8588
rect 21048 8576 21054 8628
rect 24762 8616 24768 8628
rect 24723 8588 24768 8616
rect 24762 8576 24768 8588
rect 24820 8576 24826 8628
rect 842 8508 848 8560
rect 900 8548 906 8560
rect 7098 8548 7104 8560
rect 900 8520 7104 8548
rect 900 8508 906 8520
rect 7098 8508 7104 8520
rect 7156 8508 7162 8560
rect 8481 8551 8539 8557
rect 8481 8517 8493 8551
rect 8527 8548 8539 8551
rect 9030 8548 9036 8560
rect 8527 8520 9036 8548
rect 8527 8517 8539 8520
rect 8481 8511 8539 8517
rect 9030 8508 9036 8520
rect 9088 8548 9094 8560
rect 17589 8551 17647 8557
rect 9088 8520 10088 8548
rect 9088 8508 9094 8520
rect 4522 8440 4528 8492
rect 4580 8480 4586 8492
rect 5258 8480 5264 8492
rect 4580 8452 5264 8480
rect 4580 8440 4586 8452
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 5994 8480 6000 8492
rect 5951 8452 6000 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 7006 8480 7012 8492
rect 6328 8452 7012 8480
rect 6328 8440 6334 8452
rect 7006 8440 7012 8452
rect 7064 8480 7070 8492
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 7064 8452 7205 8480
rect 7064 8440 7070 8452
rect 7193 8449 7205 8452
rect 7239 8449 7251 8483
rect 9950 8480 9956 8492
rect 7193 8443 7251 8449
rect 9048 8452 9956 8480
rect 8570 8412 8576 8424
rect 8531 8384 8576 8412
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 9048 8421 9076 8452
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 9033 8415 9091 8421
rect 9033 8412 9045 8415
rect 8904 8384 9045 8412
rect 8904 8372 8910 8384
rect 9033 8381 9045 8384
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 9401 8415 9459 8421
rect 9401 8381 9413 8415
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 9861 8415 9919 8421
rect 9861 8381 9873 8415
rect 9907 8412 9919 8415
rect 10060 8412 10088 8520
rect 17589 8517 17601 8551
rect 17635 8548 17647 8551
rect 17635 8520 20024 8548
rect 17635 8517 17647 8520
rect 17589 8511 17647 8517
rect 12066 8440 12072 8492
rect 12124 8480 12130 8492
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 12124 8452 12449 8480
rect 12124 8440 12130 8452
rect 12437 8449 12449 8452
rect 12483 8480 12495 8483
rect 14001 8483 14059 8489
rect 14001 8480 14013 8483
rect 12483 8452 14013 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 14001 8449 14013 8452
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 14090 8440 14096 8492
rect 14148 8480 14154 8492
rect 17034 8480 17040 8492
rect 14148 8452 17040 8480
rect 14148 8440 14154 8452
rect 17034 8440 17040 8452
rect 17092 8480 17098 8492
rect 17129 8483 17187 8489
rect 17129 8480 17141 8483
rect 17092 8452 17141 8480
rect 17092 8440 17098 8452
rect 17129 8449 17141 8452
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 9907 8384 10088 8412
rect 11333 8415 11391 8421
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 11333 8381 11345 8415
rect 11379 8412 11391 8415
rect 13078 8412 13084 8424
rect 11379 8384 13084 8412
rect 11379 8381 11391 8384
rect 11333 8375 11391 8381
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8344 5135 8347
rect 5353 8347 5411 8353
rect 5353 8344 5365 8347
rect 5123 8316 5365 8344
rect 5123 8313 5135 8316
rect 5077 8307 5135 8313
rect 5353 8313 5365 8316
rect 5399 8313 5411 8347
rect 6914 8344 6920 8356
rect 5353 8307 5411 8313
rect 6012 8316 6684 8344
rect 6875 8316 6920 8344
rect 5368 8276 5396 8307
rect 6012 8276 6040 8316
rect 6178 8276 6184 8288
rect 5368 8248 6040 8276
rect 6139 8248 6184 8276
rect 6178 8236 6184 8248
rect 6236 8236 6242 8288
rect 6656 8285 6684 8316
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7009 8347 7067 8353
rect 7009 8313 7021 8347
rect 7055 8344 7067 8347
rect 7282 8344 7288 8356
rect 7055 8316 7288 8344
rect 7055 8313 7067 8316
rect 7009 8307 7067 8313
rect 6641 8279 6699 8285
rect 6641 8245 6653 8279
rect 6687 8276 6699 8279
rect 7024 8276 7052 8307
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 8018 8304 8024 8356
rect 8076 8344 8082 8356
rect 8478 8344 8484 8356
rect 8076 8316 8484 8344
rect 8076 8304 8082 8316
rect 8478 8304 8484 8316
rect 8536 8344 8542 8356
rect 9416 8344 9444 8375
rect 13078 8372 13084 8384
rect 13136 8412 13142 8424
rect 13633 8415 13691 8421
rect 13633 8412 13645 8415
rect 13136 8384 13645 8412
rect 13136 8372 13142 8384
rect 13633 8381 13645 8384
rect 13679 8381 13691 8415
rect 13633 8375 13691 8381
rect 14826 8372 14832 8424
rect 14884 8412 14890 8424
rect 16758 8421 16764 8424
rect 14921 8415 14979 8421
rect 14921 8412 14933 8415
rect 14884 8384 14933 8412
rect 14884 8372 14890 8384
rect 14921 8381 14933 8384
rect 14967 8381 14979 8415
rect 16736 8415 16764 8421
rect 16736 8412 16748 8415
rect 16671 8384 16748 8412
rect 14921 8375 14979 8381
rect 16736 8381 16748 8384
rect 16816 8412 16822 8424
rect 17604 8412 17632 8511
rect 19996 8492 20024 8520
rect 19337 8483 19395 8489
rect 19337 8449 19349 8483
rect 19383 8480 19395 8483
rect 19426 8480 19432 8492
rect 19383 8452 19432 8480
rect 19383 8449 19395 8452
rect 19337 8443 19395 8449
rect 19426 8440 19432 8452
rect 19484 8440 19490 8492
rect 19978 8440 19984 8492
rect 20036 8480 20042 8492
rect 21453 8483 21511 8489
rect 21453 8480 21465 8483
rect 20036 8452 21465 8480
rect 20036 8440 20042 8452
rect 21453 8449 21465 8452
rect 21499 8449 21511 8483
rect 21453 8443 21511 8449
rect 16816 8384 17632 8412
rect 18392 8415 18450 8421
rect 16736 8375 16764 8381
rect 16758 8372 16764 8375
rect 16816 8372 16822 8384
rect 18392 8381 18404 8415
rect 18438 8412 18450 8415
rect 18782 8412 18788 8424
rect 18438 8384 18788 8412
rect 18438 8381 18450 8384
rect 18392 8375 18450 8381
rect 18782 8372 18788 8384
rect 18840 8372 18846 8424
rect 23842 8372 23848 8424
rect 23900 8412 23906 8424
rect 24581 8415 24639 8421
rect 24581 8412 24593 8415
rect 23900 8384 24593 8412
rect 23900 8372 23906 8384
rect 24581 8381 24593 8384
rect 24627 8412 24639 8415
rect 25133 8415 25191 8421
rect 25133 8412 25145 8415
rect 24627 8384 25145 8412
rect 24627 8381 24639 8384
rect 24581 8375 24639 8381
rect 25133 8381 25145 8384
rect 25179 8381 25191 8415
rect 25133 8375 25191 8381
rect 12758 8347 12816 8353
rect 12758 8344 12770 8347
rect 8536 8316 9444 8344
rect 12176 8316 12770 8344
rect 8536 8304 8542 8316
rect 8662 8276 8668 8288
rect 6687 8248 7052 8276
rect 8623 8248 8668 8276
rect 6687 8245 6699 8248
rect 6641 8239 6699 8245
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 10413 8279 10471 8285
rect 10413 8245 10425 8279
rect 10459 8276 10471 8279
rect 10778 8276 10784 8288
rect 10459 8248 10784 8276
rect 10459 8245 10471 8248
rect 10413 8239 10471 8245
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 11238 8236 11244 8288
rect 11296 8276 11302 8288
rect 11790 8276 11796 8288
rect 11296 8248 11796 8276
rect 11296 8236 11302 8248
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 12066 8236 12072 8288
rect 12124 8276 12130 8288
rect 12176 8285 12204 8316
rect 12758 8313 12770 8316
rect 12804 8313 12816 8347
rect 12758 8307 12816 8313
rect 15283 8347 15341 8353
rect 15283 8313 15295 8347
rect 15329 8313 15341 8347
rect 17770 8344 17776 8356
rect 15283 8307 15341 8313
rect 16132 8316 17776 8344
rect 12161 8279 12219 8285
rect 12161 8276 12173 8279
rect 12124 8248 12173 8276
rect 12124 8236 12130 8248
rect 12161 8245 12173 8248
rect 12207 8245 12219 8279
rect 12161 8239 12219 8245
rect 14829 8279 14887 8285
rect 14829 8245 14841 8279
rect 14875 8276 14887 8279
rect 15298 8276 15326 8307
rect 15838 8276 15844 8288
rect 14875 8248 15844 8276
rect 14875 8245 14887 8248
rect 14829 8239 14887 8245
rect 15838 8236 15844 8248
rect 15896 8276 15902 8288
rect 16132 8285 16160 8316
rect 17770 8304 17776 8316
rect 17828 8344 17834 8356
rect 18690 8344 18696 8356
rect 17828 8316 18696 8344
rect 17828 8304 17834 8316
rect 18690 8304 18696 8316
rect 18748 8344 18754 8356
rect 19153 8347 19211 8353
rect 19153 8344 19165 8347
rect 18748 8316 19165 8344
rect 18748 8304 18754 8316
rect 19153 8313 19165 8316
rect 19199 8344 19211 8347
rect 19610 8344 19616 8356
rect 19199 8316 19616 8344
rect 19199 8313 19211 8316
rect 19153 8307 19211 8313
rect 19610 8304 19616 8316
rect 19668 8353 19674 8356
rect 19668 8347 19716 8353
rect 19668 8313 19670 8347
rect 19704 8313 19716 8347
rect 21174 8344 21180 8356
rect 21135 8316 21180 8344
rect 19668 8307 19716 8313
rect 19668 8304 19674 8307
rect 21174 8304 21180 8316
rect 21232 8304 21238 8356
rect 21266 8304 21272 8356
rect 21324 8344 21330 8356
rect 21324 8316 21369 8344
rect 21324 8304 21330 8316
rect 16117 8279 16175 8285
rect 16117 8276 16129 8279
rect 15896 8248 16129 8276
rect 15896 8236 15902 8248
rect 16117 8245 16129 8248
rect 16163 8245 16175 8279
rect 16117 8239 16175 8245
rect 16390 8236 16396 8288
rect 16448 8276 16454 8288
rect 16807 8279 16865 8285
rect 16807 8276 16819 8279
rect 16448 8248 16819 8276
rect 16448 8236 16454 8248
rect 16807 8245 16819 8248
rect 16853 8245 16865 8279
rect 16807 8239 16865 8245
rect 20257 8279 20315 8285
rect 20257 8245 20269 8279
rect 20303 8276 20315 8279
rect 20622 8276 20628 8288
rect 20303 8248 20628 8276
rect 20303 8245 20315 8248
rect 20257 8239 20315 8245
rect 20622 8236 20628 8248
rect 20680 8236 20686 8288
rect 21284 8276 21312 8304
rect 22097 8279 22155 8285
rect 22097 8276 22109 8279
rect 21284 8248 22109 8276
rect 22097 8245 22109 8248
rect 22143 8245 22155 8279
rect 22097 8239 22155 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 5258 8072 5264 8084
rect 5219 8044 5264 8072
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5583 8075 5641 8081
rect 5583 8041 5595 8075
rect 5629 8072 5641 8075
rect 6914 8072 6920 8084
rect 5629 8044 6920 8072
rect 5629 8041 5641 8044
rect 5583 8035 5641 8041
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 7466 8072 7472 8084
rect 7427 8044 7472 8072
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 10134 8032 10140 8084
rect 10192 8072 10198 8084
rect 10229 8075 10287 8081
rect 10229 8072 10241 8075
rect 10192 8044 10241 8072
rect 10192 8032 10198 8044
rect 10229 8041 10241 8044
rect 10275 8041 10287 8075
rect 10229 8035 10287 8041
rect 13170 8032 13176 8084
rect 13228 8072 13234 8084
rect 13265 8075 13323 8081
rect 13265 8072 13277 8075
rect 13228 8044 13277 8072
rect 13228 8032 13234 8044
rect 13265 8041 13277 8044
rect 13311 8072 13323 8075
rect 13541 8075 13599 8081
rect 13541 8072 13553 8075
rect 13311 8044 13553 8072
rect 13311 8041 13323 8044
rect 13265 8035 13323 8041
rect 13541 8041 13553 8044
rect 13587 8041 13599 8075
rect 15470 8072 15476 8084
rect 15431 8044 15476 8072
rect 13541 8035 13599 8041
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 18782 8032 18788 8084
rect 18840 8072 18846 8084
rect 22370 8072 22376 8084
rect 18840 8044 22376 8072
rect 18840 8032 18846 8044
rect 22370 8032 22376 8044
rect 22428 8032 22434 8084
rect 6270 8004 6276 8016
rect 6231 7976 6276 8004
rect 6270 7964 6276 7976
rect 6328 7964 6334 8016
rect 6638 8004 6644 8016
rect 6599 7976 6644 8004
rect 6638 7964 6644 7976
rect 6696 7964 6702 8016
rect 9953 8007 10011 8013
rect 9953 8004 9965 8007
rect 8680 7976 9965 8004
rect 5512 7939 5570 7945
rect 5512 7905 5524 7939
rect 5558 7936 5570 7939
rect 6086 7936 6092 7948
rect 5558 7908 6092 7936
rect 5558 7905 5570 7908
rect 5512 7899 5570 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 8570 7896 8576 7948
rect 8628 7936 8634 7948
rect 8680 7945 8708 7976
rect 9953 7973 9965 7976
rect 9999 8004 10011 8007
rect 10042 8004 10048 8016
rect 9999 7976 10048 8004
rect 9999 7973 10011 7976
rect 9953 7967 10011 7973
rect 10042 7964 10048 7976
rect 10100 8004 10106 8016
rect 10100 7976 10824 8004
rect 10100 7964 10106 7976
rect 8665 7939 8723 7945
rect 8665 7936 8677 7939
rect 8628 7908 8677 7936
rect 8628 7896 8634 7908
rect 8665 7905 8677 7908
rect 8711 7905 8723 7939
rect 8665 7899 8723 7905
rect 10134 7896 10140 7948
rect 10192 7936 10198 7948
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 10192 7908 10517 7936
rect 10192 7896 10198 7908
rect 10505 7905 10517 7908
rect 10551 7936 10563 7939
rect 10686 7936 10692 7948
rect 10551 7908 10692 7936
rect 10551 7905 10563 7908
rect 10505 7899 10563 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 10796 7945 10824 7976
rect 12066 7964 12072 8016
rect 12124 8004 12130 8016
rect 12666 8007 12724 8013
rect 12666 8004 12678 8007
rect 12124 7976 12678 8004
rect 12124 7964 12130 7976
rect 12666 7973 12678 7976
rect 12712 7973 12724 8007
rect 12666 7967 12724 7973
rect 15838 7964 15844 8016
rect 15896 8004 15902 8016
rect 16530 8007 16588 8013
rect 16530 8004 16542 8007
rect 15896 7976 16542 8004
rect 15896 7964 15902 7976
rect 16530 7973 16542 7976
rect 16576 7973 16588 8007
rect 16530 7967 16588 7973
rect 19334 7964 19340 8016
rect 19392 8004 19398 8016
rect 19429 8007 19487 8013
rect 19429 8004 19441 8007
rect 19392 7976 19441 8004
rect 19392 7964 19398 7976
rect 19429 7973 19441 7976
rect 19475 7973 19487 8007
rect 19978 8004 19984 8016
rect 19939 7976 19984 8004
rect 19429 7967 19487 7973
rect 19978 7964 19984 7976
rect 20036 7964 20042 8016
rect 20622 7964 20628 8016
rect 20680 8004 20686 8016
rect 21085 8007 21143 8013
rect 21085 8004 21097 8007
rect 20680 7976 21097 8004
rect 20680 7964 20686 7976
rect 21085 7973 21097 7976
rect 21131 8004 21143 8007
rect 21358 8004 21364 8016
rect 21131 7976 21364 8004
rect 21131 7973 21143 7976
rect 21085 7967 21143 7973
rect 21358 7964 21364 7976
rect 21416 7964 21422 8016
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7936 10839 7939
rect 10870 7936 10876 7948
rect 10827 7908 10876 7936
rect 10827 7905 10839 7908
rect 10781 7899 10839 7905
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 14090 7936 14096 7948
rect 14051 7908 14096 7936
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 16206 7936 16212 7948
rect 16167 7908 16212 7936
rect 16206 7896 16212 7908
rect 16264 7896 16270 7948
rect 16942 7896 16948 7948
rect 17000 7936 17006 7948
rect 17770 7936 17776 7948
rect 17000 7908 17776 7936
rect 17000 7896 17006 7908
rect 17770 7896 17776 7908
rect 17828 7936 17834 7948
rect 17992 7939 18050 7945
rect 17992 7936 18004 7939
rect 17828 7908 18004 7936
rect 17828 7896 17834 7908
rect 17992 7905 18004 7908
rect 18038 7905 18050 7939
rect 22462 7936 22468 7948
rect 22423 7908 22468 7936
rect 17992 7899 18050 7905
rect 22462 7896 22468 7908
rect 22520 7896 22526 7948
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 6549 7871 6607 7877
rect 6549 7868 6561 7871
rect 6052 7840 6561 7868
rect 6052 7828 6058 7840
rect 6549 7837 6561 7840
rect 6595 7837 6607 7871
rect 7190 7868 7196 7880
rect 7151 7840 7196 7868
rect 6549 7831 6607 7837
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 11238 7868 11244 7880
rect 11199 7840 11244 7868
rect 11238 7828 11244 7840
rect 11296 7828 11302 7880
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7868 11943 7871
rect 12342 7868 12348 7880
rect 11931 7840 12348 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 19153 7871 19211 7877
rect 19153 7837 19165 7871
rect 19199 7868 19211 7871
rect 19337 7871 19395 7877
rect 19337 7868 19349 7871
rect 19199 7840 19349 7868
rect 19199 7837 19211 7840
rect 19153 7831 19211 7837
rect 19337 7837 19349 7840
rect 19383 7868 19395 7871
rect 19978 7868 19984 7880
rect 19383 7840 19984 7868
rect 19383 7837 19395 7840
rect 19337 7831 19395 7837
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 20990 7868 20996 7880
rect 20951 7840 20996 7868
rect 20990 7828 20996 7840
rect 21048 7828 21054 7880
rect 21269 7871 21327 7877
rect 21269 7837 21281 7871
rect 21315 7837 21327 7871
rect 21269 7831 21327 7837
rect 5534 7760 5540 7812
rect 5592 7800 5598 7812
rect 5905 7803 5963 7809
rect 5905 7800 5917 7803
rect 5592 7772 5917 7800
rect 5592 7760 5598 7772
rect 5905 7769 5917 7772
rect 5951 7800 5963 7803
rect 8662 7800 8668 7812
rect 5951 7772 8668 7800
rect 5951 7769 5963 7772
rect 5905 7763 5963 7769
rect 8662 7760 8668 7772
rect 8720 7760 8726 7812
rect 10594 7800 10600 7812
rect 10555 7772 10600 7800
rect 10594 7760 10600 7772
rect 10652 7760 10658 7812
rect 17402 7760 17408 7812
rect 17460 7800 17466 7812
rect 21284 7800 21312 7831
rect 17460 7772 21312 7800
rect 17460 7760 17466 7772
rect 8202 7692 8208 7744
rect 8260 7732 8266 7744
rect 8297 7735 8355 7741
rect 8297 7732 8309 7735
rect 8260 7704 8309 7732
rect 8260 7692 8266 7704
rect 8297 7701 8309 7704
rect 8343 7701 8355 7735
rect 8297 7695 8355 7701
rect 8846 7692 8852 7744
rect 8904 7732 8910 7744
rect 9033 7735 9091 7741
rect 9033 7732 9045 7735
rect 8904 7704 9045 7732
rect 8904 7692 8910 7704
rect 9033 7701 9045 7704
rect 9079 7701 9091 7735
rect 9033 7695 9091 7701
rect 12253 7735 12311 7741
rect 12253 7701 12265 7735
rect 12299 7732 12311 7735
rect 12434 7732 12440 7744
rect 12299 7704 12440 7732
rect 12299 7701 12311 7704
rect 12253 7695 12311 7701
rect 12434 7692 12440 7704
rect 12492 7692 12498 7744
rect 14231 7735 14289 7741
rect 14231 7701 14243 7735
rect 14277 7732 14289 7735
rect 14734 7732 14740 7744
rect 14277 7704 14740 7732
rect 14277 7701 14289 7704
rect 14231 7695 14289 7701
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 14921 7735 14979 7741
rect 14921 7732 14933 7735
rect 14884 7704 14933 7732
rect 14884 7692 14890 7704
rect 14921 7701 14933 7704
rect 14967 7701 14979 7735
rect 16022 7732 16028 7744
rect 15983 7704 16028 7732
rect 14921 7695 14979 7701
rect 16022 7692 16028 7704
rect 16080 7692 16086 7744
rect 17126 7732 17132 7744
rect 17087 7704 17132 7732
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 17494 7692 17500 7744
rect 17552 7732 17558 7744
rect 18095 7735 18153 7741
rect 18095 7732 18107 7735
rect 17552 7704 18107 7732
rect 17552 7692 17558 7704
rect 18095 7701 18107 7704
rect 18141 7701 18153 7735
rect 18095 7695 18153 7701
rect 18509 7735 18567 7741
rect 18509 7701 18521 7735
rect 18555 7732 18567 7735
rect 18598 7732 18604 7744
rect 18555 7704 18604 7732
rect 18555 7701 18567 7704
rect 18509 7695 18567 7701
rect 18598 7692 18604 7704
rect 18656 7692 18662 7744
rect 21266 7692 21272 7744
rect 21324 7732 21330 7744
rect 22005 7735 22063 7741
rect 22005 7732 22017 7735
rect 21324 7704 22017 7732
rect 21324 7692 21330 7704
rect 22005 7701 22017 7704
rect 22051 7732 22063 7735
rect 22603 7735 22661 7741
rect 22603 7732 22615 7735
rect 22051 7704 22615 7732
rect 22051 7701 22063 7704
rect 22005 7695 22063 7701
rect 22603 7701 22615 7704
rect 22649 7701 22661 7735
rect 22603 7695 22661 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 6086 7488 6092 7540
rect 6144 7528 6150 7540
rect 6181 7531 6239 7537
rect 6181 7528 6193 7531
rect 6144 7500 6193 7528
rect 6144 7488 6150 7500
rect 6181 7497 6193 7500
rect 6227 7528 6239 7531
rect 6270 7528 6276 7540
rect 6227 7500 6276 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 8113 7531 8171 7537
rect 8113 7497 8125 7531
rect 8159 7528 8171 7531
rect 8570 7528 8576 7540
rect 8159 7500 8576 7528
rect 8159 7497 8171 7500
rect 8113 7491 8171 7497
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 13722 7528 13728 7540
rect 13683 7500 13728 7528
rect 13722 7488 13728 7500
rect 13780 7528 13786 7540
rect 15657 7531 15715 7537
rect 13780 7500 14780 7528
rect 13780 7488 13786 7500
rect 1578 7460 1584 7472
rect 1539 7432 1584 7460
rect 1578 7420 1584 7432
rect 1636 7420 1642 7472
rect 14090 7460 14096 7472
rect 14051 7432 14096 7460
rect 14090 7420 14096 7432
rect 14148 7420 14154 7472
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 5951 7364 6561 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 6549 7361 6561 7364
rect 6595 7392 6607 7395
rect 6638 7392 6644 7404
rect 6595 7364 6644 7392
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 6638 7352 6644 7364
rect 6696 7352 6702 7404
rect 6917 7395 6975 7401
rect 6917 7361 6929 7395
rect 6963 7392 6975 7395
rect 7006 7392 7012 7404
rect 6963 7364 7012 7392
rect 6963 7361 6975 7364
rect 6917 7355 6975 7361
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 7190 7392 7196 7404
rect 7151 7364 7196 7392
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 12158 7392 12164 7404
rect 11072 7364 12164 7392
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7324 1458 7336
rect 1949 7327 2007 7333
rect 1949 7324 1961 7327
rect 1452 7296 1961 7324
rect 1452 7284 1458 7296
rect 1949 7293 1961 7296
rect 1995 7293 2007 7327
rect 1949 7287 2007 7293
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7324 5135 7327
rect 5813 7327 5871 7333
rect 5813 7324 5825 7327
rect 5123 7296 5825 7324
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 5813 7293 5825 7296
rect 5859 7324 5871 7327
rect 9033 7327 9091 7333
rect 5859 7296 6684 7324
rect 5859 7293 5871 7296
rect 5813 7287 5871 7293
rect 6656 7188 6684 7296
rect 9033 7293 9045 7327
rect 9079 7293 9091 7327
rect 9033 7287 9091 7293
rect 7009 7259 7067 7265
rect 7009 7225 7021 7259
rect 7055 7256 7067 7259
rect 7558 7256 7564 7268
rect 7055 7228 7564 7256
rect 7055 7225 7067 7228
rect 7009 7219 7067 7225
rect 7024 7188 7052 7219
rect 7558 7216 7564 7228
rect 7616 7216 7622 7268
rect 8846 7216 8852 7268
rect 8904 7256 8910 7268
rect 8941 7259 8999 7265
rect 8941 7256 8953 7259
rect 8904 7228 8953 7256
rect 8904 7216 8910 7228
rect 8941 7225 8953 7228
rect 8987 7225 8999 7259
rect 8941 7219 8999 7225
rect 9048 7256 9076 7287
rect 10962 7284 10968 7336
rect 11020 7324 11026 7336
rect 11072 7333 11100 7364
rect 12158 7352 12164 7364
rect 12216 7392 12222 7404
rect 12216 7364 13032 7392
rect 12216 7352 12222 7364
rect 11057 7327 11115 7333
rect 11057 7324 11069 7327
rect 11020 7296 11069 7324
rect 11020 7284 11026 7296
rect 11057 7293 11069 7296
rect 11103 7293 11115 7327
rect 11057 7287 11115 7293
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 11333 7327 11391 7333
rect 11333 7324 11345 7327
rect 11296 7296 11345 7324
rect 11296 7284 11302 7296
rect 11333 7293 11345 7296
rect 11379 7324 11391 7327
rect 12434 7324 12440 7336
rect 11379 7296 11744 7324
rect 12395 7296 12440 7324
rect 11379 7293 11391 7296
rect 11333 7287 11391 7293
rect 10505 7259 10563 7265
rect 10505 7256 10517 7259
rect 9048 7228 10517 7256
rect 8386 7188 8392 7200
rect 6656 7160 7052 7188
rect 8347 7160 8392 7188
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 8754 7188 8760 7200
rect 8715 7160 8760 7188
rect 8754 7148 8760 7160
rect 8812 7188 8818 7200
rect 9048 7188 9076 7228
rect 10505 7225 10517 7228
rect 10551 7256 10563 7259
rect 10594 7256 10600 7268
rect 10551 7228 10600 7256
rect 10551 7225 10563 7228
rect 10505 7219 10563 7225
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 11514 7256 11520 7268
rect 11475 7228 11520 7256
rect 11514 7216 11520 7228
rect 11572 7216 11578 7268
rect 11716 7256 11744 7296
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 12544 7296 12909 7324
rect 12544 7256 12572 7296
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 13004 7324 13032 7364
rect 14550 7324 14556 7336
rect 13004 7296 14556 7324
rect 12897 7287 12955 7293
rect 14550 7284 14556 7296
rect 14608 7284 14614 7336
rect 14752 7333 14780 7500
rect 15657 7497 15669 7531
rect 15703 7528 15715 7531
rect 16298 7528 16304 7540
rect 15703 7500 16304 7528
rect 15703 7497 15715 7500
rect 15657 7491 15715 7497
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 19153 7531 19211 7537
rect 19153 7497 19165 7531
rect 19199 7528 19211 7531
rect 19334 7528 19340 7540
rect 19199 7500 19340 7528
rect 19199 7497 19211 7500
rect 19153 7491 19211 7497
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 22462 7528 22468 7540
rect 22423 7500 22468 7528
rect 22462 7488 22468 7500
rect 22520 7488 22526 7540
rect 16758 7460 16764 7472
rect 16719 7432 16764 7460
rect 16758 7420 16764 7432
rect 16816 7420 16822 7472
rect 20257 7463 20315 7469
rect 20257 7429 20269 7463
rect 20303 7460 20315 7463
rect 21174 7460 21180 7472
rect 20303 7432 21180 7460
rect 20303 7429 20315 7432
rect 20257 7423 20315 7429
rect 21174 7420 21180 7432
rect 21232 7420 21238 7472
rect 14826 7352 14832 7404
rect 14884 7392 14890 7404
rect 14884 7364 14929 7392
rect 14884 7352 14890 7364
rect 16022 7352 16028 7404
rect 16080 7392 16086 7404
rect 16209 7395 16267 7401
rect 16209 7392 16221 7395
rect 16080 7364 16221 7392
rect 16080 7352 16086 7364
rect 16209 7361 16221 7364
rect 16255 7392 16267 7395
rect 17402 7392 17408 7404
rect 16255 7364 17408 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 18598 7392 18604 7404
rect 18559 7364 18604 7392
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 19705 7395 19763 7401
rect 19705 7361 19717 7395
rect 19751 7392 19763 7395
rect 20346 7392 20352 7404
rect 19751 7364 20352 7392
rect 19751 7361 19763 7364
rect 19705 7355 19763 7361
rect 20346 7352 20352 7364
rect 20404 7352 20410 7404
rect 21266 7392 21272 7404
rect 21227 7364 21272 7392
rect 21266 7352 21272 7364
rect 21324 7352 21330 7404
rect 21542 7392 21548 7404
rect 21503 7364 21548 7392
rect 21542 7352 21548 7364
rect 21600 7352 21606 7404
rect 14737 7327 14795 7333
rect 14737 7293 14749 7327
rect 14783 7293 14795 7327
rect 14737 7287 14795 7293
rect 17310 7284 17316 7336
rect 17368 7324 17374 7336
rect 17957 7327 18015 7333
rect 17957 7324 17969 7327
rect 17368 7296 17969 7324
rect 17368 7284 17374 7296
rect 11716 7228 12572 7256
rect 11716 7200 11744 7228
rect 16298 7216 16304 7268
rect 16356 7256 16362 7268
rect 16356 7228 16401 7256
rect 16356 7216 16362 7228
rect 8812 7160 9076 7188
rect 10229 7191 10287 7197
rect 8812 7148 8818 7160
rect 10229 7157 10241 7191
rect 10275 7188 10287 7191
rect 10686 7188 10692 7200
rect 10275 7160 10692 7188
rect 10275 7157 10287 7160
rect 10229 7151 10287 7157
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 11793 7191 11851 7197
rect 11793 7188 11805 7191
rect 11756 7160 11805 7188
rect 11756 7148 11762 7160
rect 11793 7157 11805 7160
rect 11839 7157 11851 7191
rect 12158 7188 12164 7200
rect 12119 7160 12164 7188
rect 11793 7151 11851 7157
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 12342 7148 12348 7200
rect 12400 7188 12406 7200
rect 12529 7191 12587 7197
rect 12529 7188 12541 7191
rect 12400 7160 12541 7188
rect 12400 7148 12406 7160
rect 12529 7157 12541 7160
rect 12575 7157 12587 7191
rect 12529 7151 12587 7157
rect 15838 7148 15844 7200
rect 15896 7188 15902 7200
rect 15933 7191 15991 7197
rect 15933 7188 15945 7191
rect 15896 7160 15945 7188
rect 15896 7148 15902 7160
rect 15933 7157 15945 7160
rect 15979 7157 15991 7191
rect 15933 7151 15991 7157
rect 16758 7148 16764 7200
rect 16816 7188 16822 7200
rect 17420 7197 17448 7296
rect 17957 7293 17969 7296
rect 18003 7293 18015 7327
rect 17957 7287 18015 7293
rect 18138 7284 18144 7336
rect 18196 7324 18202 7336
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 18196 7296 18521 7324
rect 18196 7284 18202 7296
rect 18509 7293 18521 7296
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 19797 7259 19855 7265
rect 19797 7225 19809 7259
rect 19843 7225 19855 7259
rect 19797 7219 19855 7225
rect 20993 7259 21051 7265
rect 20993 7225 21005 7259
rect 21039 7256 21051 7259
rect 21358 7256 21364 7268
rect 21039 7228 21364 7256
rect 21039 7225 21051 7228
rect 20993 7219 21051 7225
rect 17405 7191 17463 7197
rect 17405 7188 17417 7191
rect 16816 7160 17417 7188
rect 16816 7148 16822 7160
rect 17405 7157 17417 7160
rect 17451 7157 17463 7191
rect 17770 7188 17776 7200
rect 17731 7160 17776 7188
rect 17405 7151 17463 7157
rect 17770 7148 17776 7160
rect 17828 7148 17834 7200
rect 19426 7188 19432 7200
rect 19387 7160 19432 7188
rect 19426 7148 19432 7160
rect 19484 7188 19490 7200
rect 19812 7188 19840 7219
rect 21358 7216 21364 7228
rect 21416 7216 21422 7268
rect 19484 7160 19840 7188
rect 19484 7148 19490 7160
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 5994 6944 6000 6996
rect 6052 6984 6058 6996
rect 6089 6987 6147 6993
rect 6089 6984 6101 6987
rect 6052 6956 6101 6984
rect 6052 6944 6058 6956
rect 6089 6953 6101 6956
rect 6135 6953 6147 6987
rect 7558 6984 7564 6996
rect 7471 6956 7564 6984
rect 6089 6947 6147 6953
rect 7558 6944 7564 6956
rect 7616 6984 7622 6996
rect 8386 6984 8392 6996
rect 7616 6956 8392 6984
rect 7616 6944 7622 6956
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 9214 6984 9220 6996
rect 8536 6956 9220 6984
rect 8536 6944 8542 6956
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 10873 6987 10931 6993
rect 10873 6953 10885 6987
rect 10919 6984 10931 6987
rect 10962 6984 10968 6996
rect 10919 6956 10968 6984
rect 10919 6953 10931 6956
rect 10873 6947 10931 6953
rect 6962 6919 7020 6925
rect 6962 6885 6974 6919
rect 7008 6885 7020 6919
rect 6962 6879 7020 6885
rect 5534 6848 5540 6860
rect 5495 6820 5540 6848
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 6086 6808 6092 6860
rect 6144 6848 6150 6860
rect 6977 6848 7005 6879
rect 7282 6876 7288 6928
rect 7340 6916 7346 6928
rect 10888 6916 10916 6947
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 16206 6984 16212 6996
rect 16167 6956 16212 6984
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 17310 6944 17316 6996
rect 17368 6984 17374 6996
rect 20993 6987 21051 6993
rect 20993 6984 21005 6987
rect 17368 6956 21005 6984
rect 17368 6944 17374 6956
rect 20993 6953 21005 6956
rect 21039 6953 21051 6987
rect 20993 6947 21051 6953
rect 21358 6944 21364 6996
rect 21416 6984 21422 6996
rect 21913 6987 21971 6993
rect 21913 6984 21925 6987
rect 21416 6956 21925 6984
rect 21416 6944 21422 6956
rect 21913 6953 21925 6956
rect 21959 6953 21971 6987
rect 21913 6947 21971 6953
rect 24765 6987 24823 6993
rect 24765 6953 24777 6987
rect 24811 6984 24823 6987
rect 27614 6984 27620 6996
rect 24811 6956 27620 6984
rect 24811 6953 24823 6956
rect 24765 6947 24823 6953
rect 27614 6944 27620 6956
rect 27672 6944 27678 6996
rect 12437 6919 12495 6925
rect 12437 6916 12449 6919
rect 7340 6888 10916 6916
rect 11716 6888 12449 6916
rect 7340 6876 7346 6888
rect 11716 6860 11744 6888
rect 12437 6885 12449 6888
rect 12483 6916 12495 6919
rect 16758 6916 16764 6928
rect 12483 6888 13216 6916
rect 12483 6885 12495 6888
rect 12437 6879 12495 6885
rect 11330 6848 11336 6860
rect 6144 6820 7005 6848
rect 11291 6820 11336 6848
rect 6144 6808 6150 6820
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 11698 6848 11704 6860
rect 11659 6820 11704 6848
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 12066 6808 12072 6860
rect 12124 6848 12130 6860
rect 13188 6857 13216 6888
rect 13372 6888 16764 6916
rect 12713 6851 12771 6857
rect 12713 6848 12725 6851
rect 12124 6820 12725 6848
rect 12124 6808 12130 6820
rect 12713 6817 12725 6820
rect 12759 6817 12771 6851
rect 12713 6811 12771 6817
rect 13173 6851 13231 6857
rect 13173 6817 13185 6851
rect 13219 6817 13231 6851
rect 13173 6811 13231 6817
rect 6362 6740 6368 6792
rect 6420 6780 6426 6792
rect 6641 6783 6699 6789
rect 6641 6780 6653 6783
rect 6420 6752 6653 6780
rect 6420 6740 6426 6752
rect 6641 6749 6653 6752
rect 6687 6780 6699 6783
rect 8478 6780 8484 6792
rect 6687 6752 8484 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 11882 6780 11888 6792
rect 11843 6752 11888 6780
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 12728 6780 12756 6811
rect 13372 6780 13400 6888
rect 16758 6876 16764 6888
rect 16816 6876 16822 6928
rect 16853 6919 16911 6925
rect 16853 6885 16865 6919
rect 16899 6916 16911 6919
rect 17126 6916 17132 6928
rect 16899 6888 17132 6916
rect 16899 6885 16911 6888
rect 16853 6879 16911 6885
rect 17126 6876 17132 6888
rect 17184 6916 17190 6928
rect 19426 6916 19432 6928
rect 17184 6888 19432 6916
rect 17184 6876 17190 6888
rect 19426 6876 19432 6888
rect 19484 6876 19490 6928
rect 19978 6916 19984 6928
rect 19891 6888 19984 6916
rect 19978 6876 19984 6888
rect 20036 6916 20042 6928
rect 21542 6916 21548 6928
rect 20036 6888 21548 6916
rect 20036 6876 20042 6888
rect 21542 6876 21548 6888
rect 21600 6876 21606 6928
rect 23658 6876 23664 6928
rect 23716 6916 23722 6928
rect 23716 6888 24624 6916
rect 23716 6876 23722 6888
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6848 15623 6851
rect 16022 6848 16028 6860
rect 15611 6820 16028 6848
rect 15611 6817 15623 6820
rect 15565 6811 15623 6817
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 17402 6808 17408 6860
rect 17460 6848 17466 6860
rect 18138 6848 18144 6860
rect 17460 6820 17505 6848
rect 18099 6820 18144 6848
rect 17460 6808 17466 6820
rect 18138 6808 18144 6820
rect 18196 6808 18202 6860
rect 18268 6851 18326 6857
rect 18268 6848 18280 6851
rect 18248 6817 18280 6848
rect 18314 6817 18326 6851
rect 20898 6848 20904 6860
rect 20859 6820 20904 6848
rect 18248 6811 18326 6817
rect 12728 6752 13400 6780
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 15286 6780 15292 6792
rect 13495 6752 15292 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6780 16819 6783
rect 17494 6780 17500 6792
rect 16807 6752 17500 6780
rect 16807 6749 16819 6752
rect 16761 6743 16819 6749
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 18248 6780 18276 6811
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 21361 6851 21419 6857
rect 21361 6817 21373 6851
rect 21407 6817 21419 6851
rect 21361 6811 21419 6817
rect 18966 6780 18972 6792
rect 18017 6752 18972 6780
rect 10134 6712 10140 6724
rect 6840 6684 10140 6712
rect 6840 6656 6868 6684
rect 10134 6672 10140 6684
rect 10192 6712 10198 6724
rect 10413 6715 10471 6721
rect 10413 6712 10425 6715
rect 10192 6684 10425 6712
rect 10192 6672 10198 6684
rect 10413 6681 10425 6684
rect 10459 6681 10471 6715
rect 10413 6675 10471 6681
rect 14369 6715 14427 6721
rect 14369 6681 14381 6715
rect 14415 6712 14427 6715
rect 14550 6712 14556 6724
rect 14415 6684 14556 6712
rect 14415 6681 14427 6684
rect 14369 6675 14427 6681
rect 14550 6672 14556 6684
rect 14608 6712 14614 6724
rect 15378 6712 15384 6724
rect 14608 6684 15384 6712
rect 14608 6672 14614 6684
rect 15378 6672 15384 6684
rect 15436 6672 15442 6724
rect 15470 6672 15476 6724
rect 15528 6712 15534 6724
rect 18017 6712 18045 6752
rect 18966 6740 18972 6752
rect 19024 6740 19030 6792
rect 19337 6783 19395 6789
rect 19337 6749 19349 6783
rect 19383 6749 19395 6783
rect 19337 6743 19395 6749
rect 15528 6684 18045 6712
rect 18371 6715 18429 6721
rect 15528 6672 15534 6684
rect 18371 6681 18383 6715
rect 18417 6712 18429 6715
rect 19061 6715 19119 6721
rect 19061 6712 19073 6715
rect 18417 6684 19073 6712
rect 18417 6681 18429 6684
rect 18371 6675 18429 6681
rect 19061 6681 19073 6684
rect 19107 6712 19119 6715
rect 19352 6712 19380 6743
rect 20806 6740 20812 6792
rect 20864 6780 20870 6792
rect 21376 6780 21404 6811
rect 22370 6808 22376 6860
rect 22428 6848 22434 6860
rect 22500 6851 22558 6857
rect 22500 6848 22512 6851
rect 22428 6820 22512 6848
rect 22428 6808 22434 6820
rect 22500 6817 22512 6820
rect 22546 6817 22558 6851
rect 22500 6811 22558 6817
rect 23544 6851 23602 6857
rect 23544 6817 23556 6851
rect 23590 6848 23602 6851
rect 24026 6848 24032 6860
rect 23590 6820 24032 6848
rect 23590 6817 23602 6820
rect 23544 6811 23602 6817
rect 24026 6808 24032 6820
rect 24084 6808 24090 6860
rect 24596 6857 24624 6888
rect 24581 6851 24639 6857
rect 24581 6817 24593 6851
rect 24627 6848 24639 6851
rect 25498 6848 25504 6860
rect 24627 6820 25504 6848
rect 24627 6817 24639 6820
rect 24581 6811 24639 6817
rect 25498 6808 25504 6820
rect 25556 6808 25562 6860
rect 22646 6780 22652 6792
rect 20864 6752 21404 6780
rect 22607 6752 22652 6780
rect 20864 6740 20870 6752
rect 22646 6740 22652 6752
rect 22704 6740 22710 6792
rect 19107 6684 19380 6712
rect 20717 6715 20775 6721
rect 19107 6681 19119 6684
rect 19061 6675 19119 6681
rect 20717 6681 20729 6715
rect 20763 6712 20775 6715
rect 20990 6712 20996 6724
rect 20763 6684 20996 6712
rect 20763 6681 20775 6684
rect 20717 6675 20775 6681
rect 20990 6672 20996 6684
rect 21048 6712 21054 6724
rect 21048 6684 22048 6712
rect 21048 6672 21054 6684
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5442 6644 5448 6656
rect 5307 6616 5448 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 5721 6647 5779 6653
rect 5721 6613 5733 6647
rect 5767 6644 5779 6647
rect 5994 6644 6000 6656
rect 5767 6616 6000 6644
rect 5767 6613 5779 6616
rect 5721 6607 5779 6613
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 6549 6647 6607 6653
rect 6549 6613 6561 6647
rect 6595 6644 6607 6647
rect 6822 6644 6828 6656
rect 6595 6616 6828 6644
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 8846 6644 8852 6656
rect 8807 6616 8852 6644
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 15749 6647 15807 6653
rect 15749 6613 15761 6647
rect 15795 6644 15807 6647
rect 17402 6644 17408 6656
rect 15795 6616 17408 6644
rect 15795 6613 15807 6616
rect 15749 6607 15807 6613
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 18782 6644 18788 6656
rect 18743 6616 18788 6644
rect 18782 6604 18788 6616
rect 18840 6604 18846 6656
rect 20346 6644 20352 6656
rect 20307 6616 20352 6644
rect 20346 6604 20352 6616
rect 20404 6604 20410 6656
rect 22020 6644 22048 6684
rect 22094 6672 22100 6724
rect 22152 6712 22158 6724
rect 23615 6715 23673 6721
rect 23615 6712 23627 6715
rect 22152 6684 23627 6712
rect 22152 6672 22158 6684
rect 23615 6681 23627 6684
rect 23661 6681 23673 6715
rect 23615 6675 23673 6681
rect 23750 6644 23756 6656
rect 22020 6616 23756 6644
rect 23750 6604 23756 6616
rect 23808 6604 23814 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 14 6400 20 6452
rect 72 6440 78 6452
rect 16022 6440 16028 6452
rect 72 6412 4154 6440
rect 15983 6412 16028 6440
rect 72 6400 78 6412
rect 4126 6304 4154 6412
rect 16022 6400 16028 6412
rect 16080 6440 16086 6452
rect 16715 6443 16773 6449
rect 16715 6440 16727 6443
rect 16080 6412 16727 6440
rect 16080 6400 16086 6412
rect 16715 6409 16727 6412
rect 16761 6409 16773 6443
rect 17126 6440 17132 6452
rect 17087 6412 17132 6440
rect 16715 6403 16773 6409
rect 17126 6400 17132 6412
rect 17184 6400 17190 6452
rect 17494 6440 17500 6452
rect 17455 6412 17500 6440
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 18966 6400 18972 6452
rect 19024 6440 19030 6452
rect 19061 6443 19119 6449
rect 19061 6440 19073 6443
rect 19024 6412 19073 6440
rect 19024 6400 19030 6412
rect 19061 6409 19073 6412
rect 19107 6409 19119 6443
rect 19426 6440 19432 6452
rect 19387 6412 19432 6440
rect 19061 6403 19119 6409
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 20898 6440 20904 6452
rect 20859 6412 20904 6440
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 22370 6400 22376 6452
rect 22428 6440 22434 6452
rect 22465 6443 22523 6449
rect 22465 6440 22477 6443
rect 22428 6412 22477 6440
rect 22428 6400 22434 6412
rect 22465 6409 22477 6412
rect 22511 6409 22523 6443
rect 25498 6440 25504 6452
rect 25459 6412 25504 6440
rect 22465 6403 22523 6409
rect 25498 6400 25504 6412
rect 25556 6400 25562 6452
rect 5997 6375 6055 6381
rect 5997 6341 6009 6375
rect 6043 6372 6055 6375
rect 11146 6372 11152 6384
rect 6043 6344 11152 6372
rect 6043 6341 6055 6344
rect 5997 6335 6055 6341
rect 6546 6304 6552 6316
rect 4126 6276 6552 6304
rect 5184 6245 5212 6276
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 8754 6304 8760 6316
rect 6687 6276 8760 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 6932 6248 6960 6276
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 8846 6264 8852 6316
rect 8904 6304 8910 6316
rect 9950 6304 9956 6316
rect 8904 6276 9956 6304
rect 8904 6264 8910 6276
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6236 5135 6239
rect 5169 6239 5227 6245
rect 5169 6236 5181 6239
rect 5123 6208 5181 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 5169 6205 5181 6208
rect 5215 6205 5227 6239
rect 5169 6199 5227 6205
rect 5258 6196 5264 6248
rect 5316 6236 5322 6248
rect 5442 6236 5448 6248
rect 5316 6208 5361 6236
rect 5403 6208 5448 6236
rect 5316 6196 5322 6208
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 6822 6236 6828 6248
rect 6783 6208 6828 6236
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7098 6236 7104 6248
rect 6972 6208 7017 6236
rect 7059 6208 7104 6236
rect 6972 6196 6978 6208
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 8297 6239 8355 6245
rect 8297 6205 8309 6239
rect 8343 6236 8355 6239
rect 8570 6236 8576 6248
rect 8343 6208 8576 6236
rect 8343 6205 8355 6208
rect 8297 6199 8355 6205
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 9140 6245 9168 6276
rect 9950 6264 9956 6276
rect 10008 6264 10014 6316
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9769 6239 9827 6245
rect 9272 6208 9317 6236
rect 9272 6196 9278 6208
rect 9769 6205 9781 6239
rect 9815 6205 9827 6239
rect 10612 6236 10640 6344
rect 11146 6332 11152 6344
rect 11204 6372 11210 6384
rect 17586 6372 17592 6384
rect 11204 6344 17592 6372
rect 11204 6332 11210 6344
rect 17586 6332 17592 6344
rect 17644 6332 17650 6384
rect 18782 6332 18788 6384
rect 18840 6372 18846 6384
rect 22094 6372 22100 6384
rect 18840 6344 22100 6372
rect 18840 6332 18846 6344
rect 10689 6307 10747 6313
rect 10689 6273 10701 6307
rect 10735 6304 10747 6307
rect 10735 6276 11284 6304
rect 10735 6273 10747 6276
rect 10689 6267 10747 6273
rect 10778 6236 10784 6248
rect 10612 6208 10784 6236
rect 9769 6199 9827 6205
rect 7558 6168 7564 6180
rect 7519 6140 7564 6168
rect 7558 6128 7564 6140
rect 7616 6128 7622 6180
rect 6086 6060 6092 6112
rect 6144 6100 6150 6112
rect 6181 6103 6239 6109
rect 6181 6100 6193 6103
rect 6144 6072 6193 6100
rect 6144 6060 6150 6072
rect 6181 6069 6193 6072
rect 6227 6069 6239 6103
rect 7926 6100 7932 6112
rect 7887 6072 7932 6100
rect 6181 6063 6239 6069
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 8478 6100 8484 6112
rect 8439 6072 8484 6100
rect 8478 6060 8484 6072
rect 8536 6060 8542 6112
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 9784 6100 9812 6199
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 11256 6245 11284 6276
rect 11514 6264 11520 6316
rect 11572 6304 11578 6316
rect 13262 6304 13268 6316
rect 11572 6276 13268 6304
rect 11572 6264 11578 6276
rect 13262 6264 13268 6276
rect 13320 6264 13326 6316
rect 14734 6264 14740 6316
rect 14792 6304 14798 6316
rect 15105 6307 15163 6313
rect 15105 6304 15117 6307
rect 14792 6276 15117 6304
rect 14792 6264 14798 6276
rect 15105 6273 15117 6276
rect 15151 6273 15163 6307
rect 15470 6304 15476 6316
rect 15431 6276 15476 6304
rect 15105 6267 15163 6273
rect 15470 6264 15476 6276
rect 15528 6264 15534 6316
rect 19812 6313 19840 6344
rect 22094 6332 22100 6344
rect 22152 6332 22158 6384
rect 19797 6307 19855 6313
rect 19797 6273 19809 6307
rect 19843 6273 19855 6307
rect 19797 6267 19855 6273
rect 21361 6307 21419 6313
rect 21361 6273 21373 6307
rect 21407 6304 21419 6307
rect 22646 6304 22652 6316
rect 21407 6276 22652 6304
rect 21407 6273 21419 6276
rect 21361 6267 21419 6273
rect 22646 6264 22652 6276
rect 22704 6304 22710 6316
rect 22833 6307 22891 6313
rect 22833 6304 22845 6307
rect 22704 6276 22845 6304
rect 22704 6264 22710 6276
rect 22833 6273 22845 6276
rect 22879 6273 22891 6307
rect 22833 6267 22891 6273
rect 24210 6264 24216 6316
rect 24268 6304 24274 6316
rect 24811 6307 24869 6313
rect 24811 6304 24823 6307
rect 24268 6276 24823 6304
rect 24268 6264 24274 6276
rect 24811 6273 24823 6276
rect 24857 6273 24869 6307
rect 24811 6267 24869 6273
rect 11241 6239 11299 6245
rect 11241 6205 11253 6239
rect 11287 6236 11299 6239
rect 11698 6236 11704 6248
rect 11287 6208 11704 6236
rect 11287 6205 11299 6208
rect 11241 6199 11299 6205
rect 11698 6196 11704 6208
rect 11756 6236 11762 6248
rect 11793 6239 11851 6245
rect 11793 6236 11805 6239
rect 11756 6208 11805 6236
rect 11756 6196 11762 6208
rect 11793 6205 11805 6208
rect 11839 6236 11851 6239
rect 12713 6239 12771 6245
rect 12713 6236 12725 6239
rect 11839 6208 12725 6236
rect 11839 6205 11851 6208
rect 11793 6199 11851 6205
rect 12713 6205 12725 6208
rect 12759 6205 12771 6239
rect 16612 6239 16670 6245
rect 16612 6236 16624 6239
rect 12713 6199 12771 6205
rect 16408 6208 16624 6236
rect 11514 6168 11520 6180
rect 11475 6140 11520 6168
rect 11514 6128 11520 6140
rect 11572 6128 11578 6180
rect 13586 6171 13644 6177
rect 13586 6168 13598 6171
rect 13188 6140 13598 6168
rect 13188 6112 13216 6140
rect 13586 6137 13598 6140
rect 13632 6168 13644 6171
rect 15102 6168 15108 6180
rect 13632 6140 15108 6168
rect 13632 6137 13644 6140
rect 13586 6131 13644 6137
rect 15102 6128 15108 6140
rect 15160 6128 15166 6180
rect 15197 6171 15255 6177
rect 15197 6137 15209 6171
rect 15243 6137 15255 6171
rect 15197 6131 15255 6137
rect 10137 6103 10195 6109
rect 10137 6100 10149 6103
rect 9640 6072 10149 6100
rect 9640 6060 9646 6072
rect 10137 6069 10149 6072
rect 10183 6069 10195 6103
rect 10137 6063 10195 6069
rect 12066 6060 12072 6112
rect 12124 6100 12130 6112
rect 12161 6103 12219 6109
rect 12161 6100 12173 6103
rect 12124 6072 12173 6100
rect 12124 6060 12130 6072
rect 12161 6069 12173 6072
rect 12207 6069 12219 6103
rect 13170 6100 13176 6112
rect 13131 6072 13176 6100
rect 12161 6063 12219 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 14185 6103 14243 6109
rect 14185 6069 14197 6103
rect 14231 6100 14243 6103
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 14231 6072 14841 6100
rect 14231 6069 14243 6072
rect 14185 6063 14243 6069
rect 14829 6069 14841 6072
rect 14875 6100 14887 6103
rect 15212 6100 15240 6131
rect 14875 6072 15240 6100
rect 14875 6069 14887 6072
rect 14829 6063 14887 6069
rect 16114 6060 16120 6112
rect 16172 6100 16178 6112
rect 16408 6109 16436 6208
rect 16612 6205 16624 6208
rect 16658 6205 16670 6239
rect 16612 6199 16670 6205
rect 16850 6196 16856 6248
rect 16908 6236 16914 6248
rect 17773 6239 17831 6245
rect 17773 6236 17785 6239
rect 16908 6208 17785 6236
rect 16908 6196 16914 6208
rect 17773 6205 17785 6208
rect 17819 6236 17831 6239
rect 18141 6239 18199 6245
rect 18141 6236 18153 6239
rect 17819 6208 18153 6236
rect 17819 6205 17831 6208
rect 17773 6199 17831 6205
rect 18141 6205 18153 6208
rect 18187 6205 18199 6239
rect 18141 6199 18199 6205
rect 22462 6196 22468 6248
rect 22520 6236 22526 6248
rect 23728 6239 23786 6245
rect 23728 6236 23740 6239
rect 22520 6208 23740 6236
rect 22520 6196 22526 6208
rect 23728 6205 23740 6208
rect 23774 6236 23786 6239
rect 24489 6239 24547 6245
rect 24489 6236 24501 6239
rect 23774 6208 24501 6236
rect 23774 6205 23786 6208
rect 23728 6199 23786 6205
rect 24489 6205 24501 6208
rect 24535 6205 24547 6239
rect 24489 6199 24547 6205
rect 24708 6239 24766 6245
rect 24708 6205 24720 6239
rect 24754 6205 24766 6239
rect 24708 6199 24766 6205
rect 16758 6128 16764 6180
rect 16816 6168 16822 6180
rect 18049 6171 18107 6177
rect 18049 6168 18061 6171
rect 16816 6140 18061 6168
rect 16816 6128 16822 6140
rect 18049 6137 18061 6140
rect 18095 6137 18107 6171
rect 18049 6131 18107 6137
rect 19889 6171 19947 6177
rect 19889 6137 19901 6171
rect 19935 6168 19947 6171
rect 20254 6168 20260 6180
rect 19935 6140 20260 6168
rect 19935 6137 19947 6140
rect 19889 6131 19947 6137
rect 20254 6128 20260 6140
rect 20312 6128 20318 6180
rect 20438 6168 20444 6180
rect 20351 6140 20444 6168
rect 20438 6128 20444 6140
rect 20496 6168 20502 6180
rect 20496 6140 21036 6168
rect 20496 6128 20502 6140
rect 16393 6103 16451 6109
rect 16393 6100 16405 6103
rect 16172 6072 16405 6100
rect 16172 6060 16178 6072
rect 16393 6069 16405 6072
rect 16439 6069 16451 6103
rect 21008 6100 21036 6140
rect 21358 6128 21364 6180
rect 21416 6168 21422 6180
rect 21453 6171 21511 6177
rect 21453 6168 21465 6171
rect 21416 6140 21465 6168
rect 21416 6128 21422 6140
rect 21453 6137 21465 6140
rect 21499 6137 21511 6171
rect 21453 6131 21511 6137
rect 21634 6128 21640 6180
rect 21692 6168 21698 6180
rect 22005 6171 22063 6177
rect 22005 6168 22017 6171
rect 21692 6140 22017 6168
rect 21692 6128 21698 6140
rect 22005 6137 22017 6140
rect 22051 6137 22063 6171
rect 22005 6131 22063 6137
rect 22094 6128 22100 6180
rect 22152 6168 22158 6180
rect 24723 6168 24751 6199
rect 25133 6171 25191 6177
rect 25133 6168 25145 6171
rect 22152 6140 25145 6168
rect 22152 6128 22158 6140
rect 25133 6137 25145 6140
rect 25179 6137 25191 6171
rect 25133 6131 25191 6137
rect 21652 6100 21680 6128
rect 21008 6072 21680 6100
rect 16393 6063 16451 6069
rect 22554 6060 22560 6112
rect 22612 6100 22618 6112
rect 23799 6103 23857 6109
rect 23799 6100 23811 6103
rect 22612 6072 23811 6100
rect 22612 6060 22618 6072
rect 23799 6069 23811 6072
rect 23845 6069 23857 6103
rect 23799 6063 23857 6069
rect 24026 6060 24032 6112
rect 24084 6100 24090 6112
rect 24121 6103 24179 6109
rect 24121 6100 24133 6103
rect 24084 6072 24133 6100
rect 24084 6060 24090 6072
rect 24121 6069 24133 6072
rect 24167 6069 24179 6103
rect 24121 6063 24179 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 5534 5896 5540 5908
rect 5495 5868 5540 5896
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 6362 5896 6368 5908
rect 6323 5868 6368 5896
rect 6362 5856 6368 5868
rect 6420 5856 6426 5908
rect 8481 5899 8539 5905
rect 8481 5865 8493 5899
rect 8527 5896 8539 5899
rect 12434 5896 12440 5908
rect 8527 5868 12440 5896
rect 8527 5865 8539 5868
rect 8481 5859 8539 5865
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 13262 5896 13268 5908
rect 13223 5868 13268 5896
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 14274 5896 14280 5908
rect 13740 5868 14280 5896
rect 7098 5788 7104 5840
rect 7156 5828 7162 5840
rect 7561 5831 7619 5837
rect 7561 5828 7573 5831
rect 7156 5800 7573 5828
rect 7156 5788 7162 5800
rect 7561 5797 7573 5800
rect 7607 5828 7619 5831
rect 8202 5828 8208 5840
rect 7607 5800 8208 5828
rect 7607 5797 7619 5800
rect 7561 5791 7619 5797
rect 8202 5788 8208 5800
rect 8260 5828 8266 5840
rect 9306 5828 9312 5840
rect 8260 5800 9312 5828
rect 8260 5788 8266 5800
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 10413 5831 10471 5837
rect 10413 5797 10425 5831
rect 10459 5828 10471 5831
rect 12066 5828 12072 5840
rect 10459 5800 12072 5828
rect 10459 5797 10471 5800
rect 10413 5791 10471 5797
rect 12066 5788 12072 5800
rect 12124 5788 12130 5840
rect 12250 5837 12256 5840
rect 12247 5791 12256 5837
rect 12308 5828 12314 5840
rect 13170 5828 13176 5840
rect 12308 5800 13176 5828
rect 12250 5788 12256 5791
rect 12308 5788 12314 5800
rect 13170 5788 13176 5800
rect 13228 5788 13234 5840
rect 13740 5837 13768 5868
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 15013 5899 15071 5905
rect 15013 5896 15025 5899
rect 14792 5868 15025 5896
rect 14792 5856 14798 5868
rect 15013 5865 15025 5868
rect 15059 5865 15071 5899
rect 19518 5896 19524 5908
rect 15013 5859 15071 5865
rect 18984 5868 19524 5896
rect 13725 5831 13783 5837
rect 13725 5797 13737 5831
rect 13771 5797 13783 5831
rect 13725 5791 13783 5797
rect 13814 5788 13820 5840
rect 13872 5828 13878 5840
rect 13872 5800 13917 5828
rect 13872 5788 13878 5800
rect 15102 5788 15108 5840
rect 15160 5828 15166 5840
rect 15610 5831 15668 5837
rect 15610 5828 15622 5831
rect 15160 5800 15622 5828
rect 15160 5788 15166 5800
rect 15610 5797 15622 5800
rect 15656 5828 15668 5831
rect 15838 5828 15844 5840
rect 15656 5800 15844 5828
rect 15656 5797 15668 5800
rect 15610 5791 15668 5797
rect 15838 5788 15844 5800
rect 15896 5788 15902 5840
rect 17126 5788 17132 5840
rect 17184 5828 17190 5840
rect 17542 5831 17600 5837
rect 17542 5828 17554 5831
rect 17184 5800 17554 5828
rect 17184 5788 17190 5800
rect 17542 5797 17554 5800
rect 17588 5797 17600 5831
rect 17542 5791 17600 5797
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5760 6515 5763
rect 6546 5760 6552 5772
rect 6503 5732 6552 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 6730 5760 6736 5772
rect 6691 5732 6736 5760
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 7193 5763 7251 5769
rect 7193 5729 7205 5763
rect 7239 5760 7251 5763
rect 7282 5760 7288 5772
rect 7239 5732 7288 5760
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 7926 5720 7932 5772
rect 7984 5760 7990 5772
rect 8021 5763 8079 5769
rect 8021 5760 8033 5763
rect 7984 5732 8033 5760
rect 7984 5720 7990 5732
rect 8021 5729 8033 5732
rect 8067 5729 8079 5763
rect 8294 5760 8300 5772
rect 8255 5732 8300 5760
rect 8021 5723 8079 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9640 5732 9689 5760
rect 9640 5720 9646 5732
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 9953 5763 10011 5769
rect 9953 5729 9965 5763
rect 9999 5729 10011 5763
rect 10778 5760 10784 5772
rect 10739 5732 10784 5760
rect 9953 5723 10011 5729
rect 8110 5692 8116 5704
rect 8071 5664 8116 5692
rect 8110 5652 8116 5664
rect 8168 5692 8174 5704
rect 9033 5695 9091 5701
rect 9033 5692 9045 5695
rect 8168 5664 9045 5692
rect 8168 5652 8174 5664
rect 9033 5661 9045 5664
rect 9079 5692 9091 5695
rect 9214 5692 9220 5704
rect 9079 5664 9220 5692
rect 9079 5661 9091 5664
rect 9033 5655 9091 5661
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9968 5692 9996 5723
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5760 11299 5763
rect 11330 5760 11336 5772
rect 11287 5732 11336 5760
rect 11287 5729 11299 5732
rect 11241 5723 11299 5729
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 11882 5760 11888 5772
rect 11843 5732 11888 5760
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 15286 5760 15292 5772
rect 15247 5732 15292 5760
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 18984 5769 19012 5868
rect 19518 5856 19524 5868
rect 19576 5896 19582 5908
rect 22557 5899 22615 5905
rect 22557 5896 22569 5899
rect 19576 5868 22569 5896
rect 19576 5856 19582 5868
rect 22557 5865 22569 5868
rect 22603 5865 22615 5899
rect 24118 5896 24124 5908
rect 24079 5868 24124 5896
rect 22557 5859 22615 5865
rect 24118 5856 24124 5868
rect 24176 5856 24182 5908
rect 19331 5831 19389 5837
rect 19331 5797 19343 5831
rect 19377 5828 19389 5831
rect 19426 5828 19432 5840
rect 19377 5800 19432 5828
rect 19377 5797 19389 5800
rect 19331 5791 19389 5797
rect 19426 5788 19432 5800
rect 19484 5788 19490 5840
rect 21082 5828 21088 5840
rect 21043 5800 21088 5828
rect 21082 5788 21088 5800
rect 21140 5788 21146 5840
rect 21634 5828 21640 5840
rect 21595 5800 21640 5828
rect 21634 5788 21640 5800
rect 21692 5788 21698 5840
rect 18969 5763 19027 5769
rect 18969 5729 18981 5763
rect 19015 5729 19027 5763
rect 18969 5723 19027 5729
rect 22186 5720 22192 5772
rect 22244 5760 22250 5772
rect 22465 5763 22523 5769
rect 22465 5760 22477 5763
rect 22244 5732 22477 5760
rect 22244 5720 22250 5732
rect 22465 5729 22477 5732
rect 22511 5729 22523 5763
rect 22922 5760 22928 5772
rect 22883 5732 22928 5760
rect 22465 5723 22523 5729
rect 22922 5720 22928 5732
rect 22980 5720 22986 5772
rect 23382 5720 23388 5772
rect 23440 5760 23446 5772
rect 24029 5763 24087 5769
rect 24029 5760 24041 5763
rect 23440 5732 24041 5760
rect 23440 5720 23446 5732
rect 24029 5729 24041 5732
rect 24075 5729 24087 5763
rect 24029 5723 24087 5729
rect 24489 5763 24547 5769
rect 24489 5729 24501 5763
rect 24535 5729 24547 5763
rect 24489 5723 24547 5729
rect 9416 5664 9996 5692
rect 5258 5624 5264 5636
rect 5171 5596 5264 5624
rect 5258 5584 5264 5596
rect 5316 5624 5322 5636
rect 6178 5624 6184 5636
rect 5316 5596 6184 5624
rect 5316 5584 5322 5596
rect 6178 5584 6184 5596
rect 6236 5624 6242 5636
rect 6549 5627 6607 5633
rect 6549 5624 6561 5627
rect 6236 5596 6561 5624
rect 6236 5584 6242 5596
rect 6549 5593 6561 5596
rect 6595 5624 6607 5627
rect 7374 5624 7380 5636
rect 6595 5596 7380 5624
rect 6595 5593 6607 5596
rect 6549 5587 6607 5593
rect 7374 5584 7380 5596
rect 7432 5584 7438 5636
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 9416 5633 9444 5664
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14001 5695 14059 5701
rect 14001 5692 14013 5695
rect 13964 5664 14013 5692
rect 13964 5652 13970 5664
rect 14001 5661 14013 5664
rect 14047 5692 14059 5695
rect 14458 5692 14464 5704
rect 14047 5664 14464 5692
rect 14047 5661 14059 5664
rect 14001 5655 14059 5661
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 17218 5692 17224 5704
rect 17179 5664 17224 5692
rect 17218 5652 17224 5664
rect 17276 5652 17282 5704
rect 20714 5652 20720 5704
rect 20772 5692 20778 5704
rect 20993 5695 21051 5701
rect 20993 5692 21005 5695
rect 20772 5664 21005 5692
rect 20772 5652 20778 5664
rect 20993 5661 21005 5664
rect 21039 5692 21051 5695
rect 22554 5692 22560 5704
rect 21039 5664 22560 5692
rect 21039 5661 21051 5664
rect 20993 5655 21051 5661
rect 22554 5652 22560 5664
rect 22612 5652 22618 5704
rect 22940 5692 22968 5720
rect 24210 5692 24216 5704
rect 22940 5664 24216 5692
rect 24210 5652 24216 5664
rect 24268 5692 24274 5704
rect 24504 5692 24532 5723
rect 24268 5664 24532 5692
rect 24268 5652 24274 5664
rect 9401 5627 9459 5633
rect 9401 5624 9413 5627
rect 8444 5596 9413 5624
rect 8444 5584 8450 5596
rect 9401 5593 9413 5596
rect 9447 5593 9459 5627
rect 9766 5624 9772 5636
rect 9727 5596 9772 5624
rect 9401 5587 9459 5593
rect 9766 5584 9772 5596
rect 9824 5584 9830 5636
rect 18141 5627 18199 5633
rect 18141 5593 18153 5627
rect 18187 5624 18199 5627
rect 18874 5624 18880 5636
rect 18187 5596 18880 5624
rect 18187 5593 18199 5596
rect 18141 5587 18199 5593
rect 18874 5584 18880 5596
rect 18932 5624 18938 5636
rect 20254 5624 20260 5636
rect 18932 5596 20260 5624
rect 18932 5584 18938 5596
rect 20254 5584 20260 5596
rect 20312 5624 20318 5636
rect 21542 5624 21548 5636
rect 20312 5596 21548 5624
rect 20312 5584 20318 5596
rect 21542 5584 21548 5596
rect 21600 5584 21606 5636
rect 7926 5556 7932 5568
rect 7887 5528 7932 5556
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 11793 5559 11851 5565
rect 11793 5525 11805 5559
rect 11839 5556 11851 5559
rect 12066 5556 12072 5568
rect 11839 5528 12072 5556
rect 11839 5525 11851 5528
rect 11793 5519 11851 5525
rect 12066 5516 12072 5528
rect 12124 5516 12130 5568
rect 12802 5556 12808 5568
rect 12763 5528 12808 5556
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 14274 5516 14280 5568
rect 14332 5556 14338 5568
rect 14737 5559 14795 5565
rect 14737 5556 14749 5559
rect 14332 5528 14749 5556
rect 14332 5516 14338 5528
rect 14737 5525 14749 5528
rect 14783 5556 14795 5559
rect 15470 5556 15476 5568
rect 14783 5528 15476 5556
rect 14783 5525 14795 5528
rect 14737 5519 14795 5525
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 16206 5556 16212 5568
rect 16167 5528 16212 5556
rect 16206 5516 16212 5528
rect 16264 5516 16270 5568
rect 18690 5556 18696 5568
rect 18651 5528 18696 5556
rect 18690 5516 18696 5528
rect 18748 5516 18754 5568
rect 19886 5556 19892 5568
rect 19847 5528 19892 5556
rect 19886 5516 19892 5528
rect 19944 5516 19950 5568
rect 20717 5559 20775 5565
rect 20717 5525 20729 5559
rect 20763 5556 20775 5559
rect 20806 5556 20812 5568
rect 20763 5528 20812 5556
rect 20763 5525 20775 5528
rect 20717 5519 20775 5525
rect 20806 5516 20812 5528
rect 20864 5516 20870 5568
rect 21358 5516 21364 5568
rect 21416 5556 21422 5568
rect 21913 5559 21971 5565
rect 21913 5556 21925 5559
rect 21416 5528 21925 5556
rect 21416 5516 21422 5528
rect 21913 5525 21925 5528
rect 21959 5525 21971 5559
rect 21913 5519 21971 5525
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 6178 5352 6184 5364
rect 6139 5324 6184 5352
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 6730 5312 6736 5364
rect 6788 5352 6794 5364
rect 7009 5355 7067 5361
rect 7009 5352 7021 5355
rect 6788 5324 7021 5352
rect 6788 5312 6794 5324
rect 7009 5321 7021 5324
rect 7055 5352 7067 5355
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7055 5324 7389 5352
rect 7055 5321 7067 5324
rect 7009 5315 7067 5321
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 9030 5352 9036 5364
rect 8991 5324 9036 5352
rect 7377 5315 7435 5321
rect 7392 5148 7420 5315
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 13814 5312 13820 5364
rect 13872 5352 13878 5364
rect 14369 5355 14427 5361
rect 14369 5352 14381 5355
rect 13872 5324 14381 5352
rect 13872 5312 13878 5324
rect 14369 5321 14381 5324
rect 14415 5352 14427 5355
rect 16206 5352 16212 5364
rect 14415 5324 16212 5352
rect 14415 5321 14427 5324
rect 14369 5315 14427 5321
rect 16206 5312 16212 5324
rect 16264 5312 16270 5364
rect 19886 5312 19892 5364
rect 19944 5352 19950 5364
rect 20165 5355 20223 5361
rect 20165 5352 20177 5355
rect 19944 5324 20177 5352
rect 19944 5312 19950 5324
rect 20165 5321 20177 5324
rect 20211 5352 20223 5355
rect 20530 5352 20536 5364
rect 20211 5324 20536 5352
rect 20211 5321 20223 5324
rect 20165 5315 20223 5321
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 23382 5352 23388 5364
rect 23343 5324 23388 5352
rect 23382 5312 23388 5324
rect 23440 5312 23446 5364
rect 24210 5312 24216 5364
rect 24268 5352 24274 5364
rect 24489 5355 24547 5361
rect 24489 5352 24501 5355
rect 24268 5324 24501 5352
rect 24268 5312 24274 5324
rect 24489 5321 24501 5324
rect 24535 5321 24547 5355
rect 24489 5315 24547 5321
rect 9214 5284 9220 5296
rect 9175 5256 9220 5284
rect 9214 5244 9220 5256
rect 9272 5284 9278 5296
rect 15470 5284 15476 5296
rect 9272 5256 9674 5284
rect 15431 5256 15476 5284
rect 9272 5244 9278 5256
rect 9646 5216 9674 5256
rect 15470 5244 15476 5256
rect 15528 5244 15534 5296
rect 15838 5284 15844 5296
rect 15799 5256 15844 5284
rect 15838 5244 15844 5256
rect 15896 5244 15902 5296
rect 18690 5284 18696 5296
rect 18603 5256 18696 5284
rect 10689 5219 10747 5225
rect 10689 5216 10701 5219
rect 9646 5188 10701 5216
rect 10689 5185 10701 5188
rect 10735 5185 10747 5219
rect 10689 5179 10747 5185
rect 11514 5176 11520 5228
rect 11572 5216 11578 5228
rect 13078 5216 13084 5228
rect 11572 5188 13084 5216
rect 11572 5176 11578 5188
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 16666 5176 16672 5228
rect 16724 5216 16730 5228
rect 18616 5225 18644 5256
rect 18690 5244 18696 5256
rect 18748 5284 18754 5296
rect 18748 5256 21036 5284
rect 18748 5244 18754 5256
rect 16761 5219 16819 5225
rect 16761 5216 16773 5219
rect 16724 5188 16773 5216
rect 16724 5176 16730 5188
rect 16761 5185 16773 5188
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 18601 5219 18659 5225
rect 18601 5185 18613 5219
rect 18647 5185 18659 5219
rect 20438 5216 20444 5228
rect 20399 5188 20444 5216
rect 18601 5179 18659 5185
rect 20438 5176 20444 5188
rect 20496 5176 20502 5228
rect 20622 5176 20628 5228
rect 20680 5216 20686 5228
rect 20717 5219 20775 5225
rect 20717 5216 20729 5219
rect 20680 5188 20729 5216
rect 20680 5176 20686 5188
rect 20717 5185 20729 5188
rect 20763 5185 20775 5219
rect 21008 5216 21036 5256
rect 22465 5219 22523 5225
rect 22465 5216 22477 5219
rect 21008 5188 22477 5216
rect 20717 5179 20775 5185
rect 22465 5185 22477 5188
rect 22511 5185 22523 5219
rect 22465 5179 22523 5185
rect 23842 5176 23848 5228
rect 23900 5216 23906 5228
rect 23900 5188 24751 5216
rect 23900 5176 23906 5188
rect 7653 5151 7711 5157
rect 7653 5148 7665 5151
rect 7392 5120 7665 5148
rect 7653 5117 7665 5120
rect 7699 5148 7711 5151
rect 8294 5148 8300 5160
rect 7699 5120 8300 5148
rect 7699 5117 7711 5120
rect 7653 5111 7711 5117
rect 8294 5108 8300 5120
rect 8352 5148 8358 5160
rect 8573 5151 8631 5157
rect 8573 5148 8585 5151
rect 8352 5120 8585 5148
rect 8352 5108 8358 5120
rect 8573 5117 8585 5120
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 5442 5040 5448 5092
rect 5500 5080 5506 5092
rect 7561 5083 7619 5089
rect 7561 5080 7573 5083
rect 5500 5052 7573 5080
rect 5500 5040 5506 5052
rect 7561 5049 7573 5052
rect 7607 5080 7619 5083
rect 8386 5080 8392 5092
rect 7607 5052 8392 5080
rect 7607 5049 7619 5052
rect 7561 5043 7619 5049
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 8588 5080 8616 5111
rect 9030 5108 9036 5160
rect 9088 5148 9094 5160
rect 9125 5151 9183 5157
rect 9125 5148 9137 5151
rect 9088 5120 9137 5148
rect 9088 5108 9094 5120
rect 9125 5117 9137 5120
rect 9171 5117 9183 5151
rect 9125 5111 9183 5117
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5117 9459 5151
rect 9401 5111 9459 5117
rect 9416 5080 9444 5111
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 10229 5151 10287 5157
rect 10229 5148 10241 5151
rect 9824 5120 10241 5148
rect 9824 5108 9830 5120
rect 10229 5117 10241 5120
rect 10275 5148 10287 5151
rect 10597 5151 10655 5157
rect 10597 5148 10609 5151
rect 10275 5120 10609 5148
rect 10275 5117 10287 5120
rect 10229 5111 10287 5117
rect 10597 5117 10609 5120
rect 10643 5148 10655 5151
rect 11330 5148 11336 5160
rect 10643 5120 11336 5148
rect 10643 5117 10655 5120
rect 10597 5111 10655 5117
rect 11330 5108 11336 5120
rect 11388 5108 11394 5160
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5148 14059 5151
rect 14645 5151 14703 5157
rect 14645 5148 14657 5151
rect 14047 5120 14657 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 14645 5117 14657 5120
rect 14691 5117 14703 5151
rect 14645 5111 14703 5117
rect 8588 5052 9444 5080
rect 9861 5083 9919 5089
rect 9861 5049 9873 5083
rect 9907 5080 9919 5083
rect 11606 5080 11612 5092
rect 9907 5052 11612 5080
rect 9907 5049 9919 5052
rect 9861 5043 9919 5049
rect 11606 5040 11612 5052
rect 11664 5040 11670 5092
rect 13170 5080 13176 5092
rect 12912 5052 13176 5080
rect 6546 5012 6552 5024
rect 6459 4984 6552 5012
rect 6546 4972 6552 4984
rect 6604 5012 6610 5024
rect 7742 5012 7748 5024
rect 6604 4984 7748 5012
rect 6604 4972 6610 4984
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 12912 5021 12940 5052
rect 13170 5040 13176 5052
rect 13228 5080 13234 5092
rect 13402 5083 13460 5089
rect 13402 5080 13414 5083
rect 13228 5052 13414 5080
rect 13228 5040 13234 5052
rect 13402 5049 13414 5052
rect 13448 5049 13460 5083
rect 13402 5043 13460 5049
rect 11885 5015 11943 5021
rect 11885 5012 11897 5015
rect 11848 4984 11897 5012
rect 11848 4972 11854 4984
rect 11885 4981 11897 4984
rect 11931 5012 11943 5015
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 11931 4984 12909 5012
rect 11931 4981 11943 4984
rect 11885 4975 11943 4981
rect 12897 4981 12909 4984
rect 12943 4981 12955 5015
rect 14660 5012 14688 5111
rect 18690 5108 18696 5160
rect 18748 5148 18754 5160
rect 19521 5151 19579 5157
rect 18748 5120 19006 5148
rect 18748 5108 18754 5120
rect 14918 5080 14924 5092
rect 14879 5052 14924 5080
rect 14918 5040 14924 5052
rect 14976 5040 14982 5092
rect 15013 5083 15071 5089
rect 15013 5049 15025 5083
rect 15059 5049 15071 5083
rect 16482 5080 16488 5092
rect 16443 5052 16488 5080
rect 15013 5043 15071 5049
rect 15028 5012 15056 5043
rect 16482 5040 16488 5052
rect 16540 5040 16546 5092
rect 16577 5083 16635 5089
rect 16577 5049 16589 5083
rect 16623 5080 16635 5083
rect 16758 5080 16764 5092
rect 16623 5052 16764 5080
rect 16623 5049 16635 5052
rect 16577 5043 16635 5049
rect 14660 4984 15056 5012
rect 16301 5015 16359 5021
rect 12897 4975 12955 4981
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 16592 5012 16620 5043
rect 16758 5040 16764 5052
rect 16816 5040 16822 5092
rect 17218 5040 17224 5092
rect 17276 5080 17282 5092
rect 17865 5083 17923 5089
rect 17865 5080 17877 5083
rect 17276 5052 17877 5080
rect 17276 5040 17282 5052
rect 17865 5049 17877 5052
rect 17911 5080 17923 5083
rect 18782 5080 18788 5092
rect 17911 5052 18788 5080
rect 17911 5049 17923 5052
rect 17865 5043 17923 5049
rect 18782 5040 18788 5052
rect 18840 5040 18846 5092
rect 18978 5089 19006 5120
rect 19521 5117 19533 5151
rect 19567 5148 19579 5151
rect 21910 5148 21916 5160
rect 19567 5120 19885 5148
rect 21871 5120 21916 5148
rect 19567 5117 19579 5120
rect 19521 5111 19579 5117
rect 18963 5083 19021 5089
rect 18963 5049 18975 5083
rect 19009 5080 19021 5083
rect 19150 5080 19156 5092
rect 19009 5052 19156 5080
rect 19009 5049 19021 5052
rect 18963 5043 19021 5049
rect 19150 5040 19156 5052
rect 19208 5080 19214 5092
rect 19857 5080 19885 5120
rect 21910 5108 21916 5120
rect 21968 5108 21974 5160
rect 22370 5148 22376 5160
rect 22331 5120 22376 5148
rect 22370 5108 22376 5120
rect 22428 5108 22434 5160
rect 23728 5151 23786 5157
rect 23728 5117 23740 5151
rect 23774 5148 23786 5151
rect 23934 5148 23940 5160
rect 23774 5120 23940 5148
rect 23774 5117 23786 5120
rect 23728 5111 23786 5117
rect 23934 5108 23940 5120
rect 23992 5148 23998 5160
rect 24723 5157 24751 5188
rect 24121 5151 24179 5157
rect 24121 5148 24133 5151
rect 23992 5120 24133 5148
rect 23992 5108 23998 5120
rect 24121 5117 24133 5120
rect 24167 5117 24179 5151
rect 24121 5111 24179 5117
rect 24708 5151 24766 5157
rect 24708 5117 24720 5151
rect 24754 5148 24766 5151
rect 25133 5151 25191 5157
rect 25133 5148 25145 5151
rect 24754 5120 25145 5148
rect 24754 5117 24766 5120
rect 24708 5111 24766 5117
rect 25133 5117 25145 5120
rect 25179 5117 25191 5151
rect 25133 5111 25191 5117
rect 19208 5052 19472 5080
rect 19857 5052 20484 5080
rect 19208 5040 19214 5052
rect 19444 5024 19472 5052
rect 16347 4984 16620 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 17126 4972 17132 5024
rect 17184 5012 17190 5024
rect 17405 5015 17463 5021
rect 17405 5012 17417 5015
rect 17184 4984 17417 5012
rect 17184 4972 17190 4984
rect 17405 4981 17417 4984
rect 17451 5012 17463 5015
rect 18417 5015 18475 5021
rect 18417 5012 18429 5015
rect 17451 4984 18429 5012
rect 17451 4981 17463 4984
rect 17405 4975 17463 4981
rect 18417 4981 18429 4984
rect 18463 5012 18475 5015
rect 18690 5012 18696 5024
rect 18463 4984 18696 5012
rect 18463 4981 18475 4984
rect 18417 4975 18475 4981
rect 18690 4972 18696 4984
rect 18748 4972 18754 5024
rect 19426 4972 19432 5024
rect 19484 5012 19490 5024
rect 19797 5015 19855 5021
rect 19797 5012 19809 5015
rect 19484 4984 19809 5012
rect 19484 4972 19490 4984
rect 19797 4981 19809 4984
rect 19843 4981 19855 5015
rect 20456 5012 20484 5052
rect 20530 5040 20536 5092
rect 20588 5080 20594 5092
rect 20588 5052 20633 5080
rect 20588 5040 20594 5052
rect 21266 5040 21272 5092
rect 21324 5080 21330 5092
rect 24811 5083 24869 5089
rect 24811 5080 24823 5083
rect 21324 5052 24823 5080
rect 21324 5040 21330 5052
rect 24811 5049 24823 5052
rect 24857 5049 24869 5083
rect 24811 5043 24869 5049
rect 21082 5012 21088 5024
rect 20456 4984 21088 5012
rect 19797 4975 19855 4981
rect 21082 4972 21088 4984
rect 21140 5012 21146 5024
rect 21361 5015 21419 5021
rect 21361 5012 21373 5015
rect 21140 4984 21373 5012
rect 21140 4972 21146 4984
rect 21361 4981 21373 4984
rect 21407 4981 21419 5015
rect 21726 5012 21732 5024
rect 21687 4984 21732 5012
rect 21361 4975 21419 4981
rect 21726 4972 21732 4984
rect 21784 5012 21790 5024
rect 22370 5012 22376 5024
rect 21784 4984 22376 5012
rect 21784 4972 21790 4984
rect 22370 4972 22376 4984
rect 22428 5012 22434 5024
rect 22922 5012 22928 5024
rect 22428 4984 22928 5012
rect 22428 4972 22434 4984
rect 22922 4972 22928 4984
rect 22980 4972 22986 5024
rect 23474 4972 23480 5024
rect 23532 5012 23538 5024
rect 23799 5015 23857 5021
rect 23799 5012 23811 5015
rect 23532 4984 23811 5012
rect 23532 4972 23538 4984
rect 23799 4981 23811 4984
rect 23845 4981 23857 5015
rect 23799 4975 23857 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 7929 4811 7987 4817
rect 7929 4777 7941 4811
rect 7975 4808 7987 4811
rect 8110 4808 8116 4820
rect 7975 4780 8116 4808
rect 7975 4777 7987 4780
rect 7929 4771 7987 4777
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 8481 4811 8539 4817
rect 8481 4777 8493 4811
rect 8527 4808 8539 4811
rect 11238 4808 11244 4820
rect 8527 4780 11244 4808
rect 8527 4777 8539 4780
rect 8481 4771 8539 4777
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 11882 4808 11888 4820
rect 11843 4780 11888 4808
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 13078 4808 13084 4820
rect 13039 4780 13084 4808
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 15473 4811 15531 4817
rect 15473 4808 15485 4811
rect 15344 4780 15485 4808
rect 15344 4768 15350 4780
rect 15473 4777 15485 4780
rect 15519 4777 15531 4811
rect 16482 4808 16488 4820
rect 16443 4780 16488 4808
rect 15473 4771 15531 4777
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 18506 4768 18512 4820
rect 18564 4808 18570 4820
rect 18874 4808 18880 4820
rect 18564 4780 18880 4808
rect 18564 4768 18570 4780
rect 7147 4743 7205 4749
rect 7147 4709 7159 4743
rect 7193 4740 7205 4743
rect 10410 4740 10416 4752
rect 7193 4712 10416 4740
rect 7193 4709 7205 4712
rect 7147 4703 7205 4709
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 12161 4743 12219 4749
rect 12161 4709 12173 4743
rect 12207 4740 12219 4743
rect 12250 4740 12256 4752
rect 12207 4712 12256 4740
rect 12207 4709 12219 4712
rect 12161 4703 12219 4709
rect 12250 4700 12256 4712
rect 12308 4700 12314 4752
rect 12802 4700 12808 4752
rect 12860 4740 12866 4752
rect 13446 4740 13452 4752
rect 12860 4712 13452 4740
rect 12860 4700 12866 4712
rect 13446 4700 13452 4712
rect 13504 4740 13510 4752
rect 13725 4743 13783 4749
rect 13725 4740 13737 4743
rect 13504 4712 13737 4740
rect 13504 4700 13510 4712
rect 13725 4709 13737 4712
rect 13771 4709 13783 4743
rect 14274 4740 14280 4752
rect 14235 4712 14280 4740
rect 13725 4703 13783 4709
rect 14274 4700 14280 4712
rect 14332 4700 14338 4752
rect 15838 4700 15844 4752
rect 15896 4740 15902 4752
rect 17126 4749 17132 4752
rect 17082 4743 17132 4749
rect 17082 4740 17094 4743
rect 15896 4712 17094 4740
rect 15896 4700 15902 4712
rect 17082 4709 17094 4712
rect 17128 4709 17132 4743
rect 17082 4703 17132 4709
rect 17126 4700 17132 4703
rect 17184 4700 17190 4752
rect 18708 4749 18736 4780
rect 18874 4768 18880 4780
rect 18932 4768 18938 4820
rect 19518 4808 19524 4820
rect 19479 4780 19524 4808
rect 19518 4768 19524 4780
rect 19576 4768 19582 4820
rect 20349 4811 20407 4817
rect 20349 4777 20361 4811
rect 20395 4808 20407 4811
rect 20438 4808 20444 4820
rect 20395 4780 20444 4808
rect 20395 4777 20407 4780
rect 20349 4771 20407 4777
rect 20438 4768 20444 4780
rect 20496 4768 20502 4820
rect 20714 4808 20720 4820
rect 20675 4780 20720 4808
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 20993 4811 21051 4817
rect 20993 4777 21005 4811
rect 21039 4777 21051 4811
rect 21910 4808 21916 4820
rect 21871 4780 21916 4808
rect 20993 4771 21051 4777
rect 18693 4743 18751 4749
rect 18693 4709 18705 4743
rect 18739 4709 18751 4743
rect 18693 4703 18751 4709
rect 18782 4700 18788 4752
rect 18840 4740 18846 4752
rect 21008 4740 21036 4771
rect 21910 4768 21916 4780
rect 21968 4768 21974 4820
rect 22186 4768 22192 4820
rect 22244 4808 22250 4820
rect 22281 4811 22339 4817
rect 22281 4808 22293 4811
rect 22244 4780 22293 4808
rect 22244 4768 22250 4780
rect 22281 4777 22293 4780
rect 22327 4777 22339 4811
rect 22554 4808 22560 4820
rect 22515 4780 22560 4808
rect 22281 4771 22339 4777
rect 22554 4768 22560 4780
rect 22612 4768 22618 4820
rect 23290 4740 23296 4752
rect 18840 4712 21036 4740
rect 21284 4712 23296 4740
rect 18840 4700 18846 4712
rect 6546 4632 6552 4684
rect 6604 4672 6610 4684
rect 7044 4675 7102 4681
rect 7044 4672 7056 4675
rect 6604 4644 7056 4672
rect 6604 4632 6610 4644
rect 7044 4641 7056 4644
rect 7090 4641 7102 4675
rect 7044 4635 7102 4641
rect 7926 4632 7932 4684
rect 7984 4672 7990 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7984 4644 8033 4672
rect 7984 4632 7990 4644
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 8294 4672 8300 4684
rect 8255 4644 8300 4672
rect 8021 4635 8079 4641
rect 8294 4632 8300 4644
rect 8352 4672 8358 4684
rect 9125 4675 9183 4681
rect 9125 4672 9137 4675
rect 8352 4644 9137 4672
rect 8352 4632 8358 4644
rect 9125 4641 9137 4644
rect 9171 4641 9183 4675
rect 9674 4672 9680 4684
rect 9635 4644 9680 4672
rect 9125 4635 9183 4641
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 10134 4672 10140 4684
rect 10095 4644 10140 4672
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 10502 4672 10508 4684
rect 10463 4644 10508 4672
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 11057 4675 11115 4681
rect 11057 4641 11069 4675
rect 11103 4672 11115 4675
rect 11422 4672 11428 4684
rect 11103 4644 11428 4672
rect 11103 4641 11115 4644
rect 11057 4635 11115 4641
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 11072 4604 11100 4635
rect 11422 4632 11428 4644
rect 11480 4632 11486 4684
rect 14918 4672 14924 4684
rect 14879 4644 14924 4672
rect 14918 4632 14924 4644
rect 14976 4632 14982 4684
rect 15286 4632 15292 4684
rect 15344 4672 15350 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 15344 4644 15669 4672
rect 15344 4632 15350 4644
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 16761 4675 16819 4681
rect 16761 4641 16773 4675
rect 16807 4672 16819 4675
rect 17310 4672 17316 4684
rect 16807 4644 17316 4672
rect 16807 4641 16819 4644
rect 16761 4635 16819 4641
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 20898 4672 20904 4684
rect 20859 4644 20904 4672
rect 20898 4632 20904 4644
rect 20956 4672 20962 4684
rect 21284 4672 21312 4712
rect 23290 4700 23296 4712
rect 23348 4700 23354 4752
rect 20956 4644 21312 4672
rect 21361 4675 21419 4681
rect 20956 4632 20962 4644
rect 21361 4641 21373 4675
rect 21407 4641 21419 4675
rect 21361 4635 21419 4641
rect 9640 4576 11100 4604
rect 11149 4607 11207 4613
rect 9640 4564 9646 4576
rect 11149 4573 11161 4607
rect 11195 4604 11207 4607
rect 11238 4604 11244 4616
rect 11195 4576 11244 4604
rect 11195 4573 11207 4576
rect 11149 4567 11207 4573
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 12066 4604 12072 4616
rect 12027 4576 12072 4604
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 12713 4607 12771 4613
rect 12713 4573 12725 4607
rect 12759 4604 12771 4607
rect 12802 4604 12808 4616
rect 12759 4576 12808 4604
rect 12759 4573 12771 4576
rect 12713 4567 12771 4573
rect 12802 4564 12808 4576
rect 12860 4564 12866 4616
rect 13633 4607 13691 4613
rect 13633 4573 13645 4607
rect 13679 4604 13691 4607
rect 14642 4604 14648 4616
rect 13679 4576 14648 4604
rect 13679 4573 13691 4576
rect 13633 4567 13691 4573
rect 14642 4564 14648 4576
rect 14700 4564 14706 4616
rect 18601 4607 18659 4613
rect 18601 4573 18613 4607
rect 18647 4604 18659 4607
rect 18690 4604 18696 4616
rect 18647 4576 18696 4604
rect 18647 4573 18659 4576
rect 18601 4567 18659 4573
rect 18690 4564 18696 4576
rect 18748 4564 18754 4616
rect 18874 4604 18880 4616
rect 18835 4576 18880 4604
rect 18874 4564 18880 4576
rect 18932 4564 18938 4616
rect 18966 4564 18972 4616
rect 19024 4604 19030 4616
rect 20806 4604 20812 4616
rect 19024 4576 20812 4604
rect 19024 4564 19030 4576
rect 20806 4564 20812 4576
rect 20864 4604 20870 4616
rect 21376 4604 21404 4635
rect 21450 4632 21456 4684
rect 21508 4672 21514 4684
rect 22465 4675 22523 4681
rect 22465 4672 22477 4675
rect 21508 4644 22477 4672
rect 21508 4632 21514 4644
rect 22465 4641 22477 4644
rect 22511 4672 22523 4675
rect 22830 4672 22836 4684
rect 22511 4644 22836 4672
rect 22511 4641 22523 4644
rect 22465 4635 22523 4641
rect 22830 4632 22836 4644
rect 22888 4632 22894 4684
rect 22922 4632 22928 4684
rect 22980 4672 22986 4684
rect 24026 4672 24032 4684
rect 22980 4644 23025 4672
rect 23987 4644 24032 4672
rect 22980 4632 22986 4644
rect 24026 4632 24032 4644
rect 24084 4632 24090 4684
rect 25108 4675 25166 4681
rect 25108 4641 25120 4675
rect 25154 4672 25166 4675
rect 25498 4672 25504 4684
rect 25154 4644 25504 4672
rect 25154 4641 25166 4644
rect 25108 4635 25166 4641
rect 25498 4632 25504 4644
rect 25556 4632 25562 4684
rect 21726 4604 21732 4616
rect 20864 4576 21732 4604
rect 20864 4564 20870 4576
rect 21726 4564 21732 4576
rect 21784 4564 21790 4616
rect 24118 4564 24124 4616
rect 24176 4604 24182 4616
rect 24854 4604 24860 4616
rect 24176 4576 24860 4604
rect 24176 4564 24182 4576
rect 24854 4564 24860 4576
rect 24912 4564 24918 4616
rect 7466 4496 7472 4548
rect 7524 4536 7530 4548
rect 8113 4539 8171 4545
rect 8113 4536 8125 4539
rect 7524 4508 8125 4536
rect 7524 4496 7530 4508
rect 8113 4505 8125 4508
rect 8159 4536 8171 4539
rect 9766 4536 9772 4548
rect 8159 4508 9772 4536
rect 8159 4505 8171 4508
rect 8113 4499 8171 4505
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 15841 4539 15899 4545
rect 15841 4505 15853 4539
rect 15887 4536 15899 4539
rect 15887 4508 18644 4536
rect 15887 4505 15899 4508
rect 15841 4499 15899 4505
rect 18616 4480 18644 4508
rect 20990 4496 20996 4548
rect 21048 4536 21054 4548
rect 25179 4539 25237 4545
rect 25179 4536 25191 4539
rect 21048 4508 25191 4536
rect 21048 4496 21054 4508
rect 25179 4505 25191 4508
rect 25225 4505 25237 4539
rect 25179 4499 25237 4505
rect 9306 4428 9312 4480
rect 9364 4468 9370 4480
rect 9674 4468 9680 4480
rect 9364 4440 9680 4468
rect 9364 4428 9370 4440
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 11514 4468 11520 4480
rect 11475 4440 11520 4468
rect 11514 4428 11520 4440
rect 11572 4428 11578 4480
rect 14550 4468 14556 4480
rect 14511 4440 14556 4468
rect 14550 4428 14556 4440
rect 14608 4468 14614 4480
rect 15930 4468 15936 4480
rect 14608 4440 15936 4468
rect 14608 4428 14614 4440
rect 15930 4428 15936 4440
rect 15988 4428 15994 4480
rect 17681 4471 17739 4477
rect 17681 4437 17693 4471
rect 17727 4468 17739 4471
rect 17770 4468 17776 4480
rect 17727 4440 17776 4468
rect 17727 4437 17739 4440
rect 17681 4431 17739 4437
rect 17770 4428 17776 4440
rect 17828 4428 17834 4480
rect 18598 4428 18604 4480
rect 18656 4428 18662 4480
rect 22370 4428 22376 4480
rect 22428 4468 22434 4480
rect 24167 4471 24225 4477
rect 24167 4468 24179 4471
rect 22428 4440 24179 4468
rect 22428 4428 22434 4440
rect 24167 4437 24179 4440
rect 24213 4437 24225 4471
rect 24167 4431 24225 4437
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 7055 4267 7113 4273
rect 7055 4233 7067 4267
rect 7101 4264 7113 4267
rect 12066 4264 12072 4276
rect 7101 4236 12072 4264
rect 7101 4233 7113 4236
rect 7055 4227 7113 4233
rect 12066 4224 12072 4236
rect 12124 4224 12130 4276
rect 13446 4264 13452 4276
rect 13407 4236 13452 4264
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 15473 4267 15531 4273
rect 15473 4233 15485 4267
rect 15519 4264 15531 4267
rect 15746 4264 15752 4276
rect 15519 4236 15752 4264
rect 15519 4233 15531 4236
rect 15473 4227 15531 4233
rect 15746 4224 15752 4236
rect 15804 4264 15810 4276
rect 16390 4264 16396 4276
rect 15804 4236 16396 4264
rect 15804 4224 15810 4236
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 17034 4264 17040 4276
rect 16684 4236 17040 4264
rect 16684 4208 16712 4236
rect 17034 4224 17040 4236
rect 17092 4224 17098 4276
rect 17221 4267 17279 4273
rect 17221 4233 17233 4267
rect 17267 4264 17279 4267
rect 17310 4264 17316 4276
rect 17267 4236 17316 4264
rect 17267 4233 17279 4236
rect 17221 4227 17279 4233
rect 17310 4224 17316 4236
rect 17368 4224 17374 4276
rect 18506 4264 18512 4276
rect 18467 4236 18512 4264
rect 18506 4224 18512 4236
rect 18564 4224 18570 4276
rect 18782 4224 18788 4276
rect 18840 4264 18846 4276
rect 19242 4264 19248 4276
rect 18840 4236 19248 4264
rect 18840 4224 18846 4236
rect 19242 4224 19248 4236
rect 19300 4224 19306 4276
rect 20625 4267 20683 4273
rect 20625 4233 20637 4267
rect 20671 4264 20683 4267
rect 20898 4264 20904 4276
rect 20671 4236 20904 4264
rect 20671 4233 20683 4236
rect 20625 4227 20683 4233
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 21726 4264 21732 4276
rect 21687 4236 21732 4264
rect 21726 4224 21732 4236
rect 21784 4264 21790 4276
rect 22741 4267 22799 4273
rect 22741 4264 22753 4267
rect 21784 4236 22753 4264
rect 21784 4224 21790 4236
rect 22741 4233 22753 4236
rect 22787 4233 22799 4267
rect 22741 4227 22799 4233
rect 22830 4224 22836 4276
rect 22888 4264 22894 4276
rect 23109 4267 23167 4273
rect 23109 4264 23121 4267
rect 22888 4236 23121 4264
rect 22888 4224 22894 4236
rect 23109 4233 23121 4236
rect 23155 4233 23167 4267
rect 24026 4264 24032 4276
rect 23987 4236 24032 4264
rect 23109 4227 23167 4233
rect 24026 4224 24032 4236
rect 24084 4224 24090 4276
rect 25130 4264 25136 4276
rect 25091 4236 25136 4264
rect 25130 4224 25136 4236
rect 25188 4224 25194 4276
rect 7466 4196 7472 4208
rect 7427 4168 7472 4196
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 7742 4196 7748 4208
rect 7655 4168 7748 4196
rect 7742 4156 7748 4168
rect 7800 4196 7806 4208
rect 7837 4199 7895 4205
rect 7837 4196 7849 4199
rect 7800 4168 7849 4196
rect 7800 4156 7806 4168
rect 7837 4165 7849 4168
rect 7883 4196 7895 4199
rect 9030 4196 9036 4208
rect 7883 4168 9036 4196
rect 7883 4165 7895 4168
rect 7837 4159 7895 4165
rect 9030 4156 9036 4168
rect 9088 4156 9094 4208
rect 14645 4199 14703 4205
rect 14645 4165 14657 4199
rect 14691 4196 14703 4199
rect 16666 4196 16672 4208
rect 14691 4168 16672 4196
rect 14691 4165 14703 4168
rect 14645 4159 14703 4165
rect 16666 4156 16672 4168
rect 16724 4156 16730 4208
rect 19518 4156 19524 4208
rect 19576 4196 19582 4208
rect 24719 4199 24777 4205
rect 24719 4196 24731 4199
rect 19576 4168 24731 4196
rect 19576 4156 19582 4168
rect 24719 4165 24731 4168
rect 24765 4165 24777 4199
rect 24719 4159 24777 4165
rect 6273 4131 6331 4137
rect 6273 4097 6285 4131
rect 6319 4128 6331 4131
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6319 4100 6837 4128
rect 6319 4097 6331 4100
rect 6273 4091 6331 4097
rect 6825 4097 6837 4100
rect 6871 4128 6883 4131
rect 6914 4128 6920 4140
rect 6871 4100 6920 4128
rect 6871 4097 6883 4100
rect 6825 4091 6883 4097
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7760 4060 7788 4156
rect 7926 4088 7932 4140
rect 7984 4128 7990 4140
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 7984 4100 8677 4128
rect 7984 4088 7990 4100
rect 8665 4097 8677 4100
rect 8711 4128 8723 4131
rect 9582 4128 9588 4140
rect 8711 4100 9588 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 9674 4088 9680 4140
rect 9732 4128 9738 4140
rect 12161 4131 12219 4137
rect 12161 4128 12173 4131
rect 9732 4100 12173 4128
rect 9732 4088 9738 4100
rect 12161 4097 12173 4100
rect 12207 4128 12219 4131
rect 12526 4128 12532 4140
rect 12207 4100 12532 4128
rect 12207 4097 12219 4100
rect 12161 4091 12219 4097
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 12802 4128 12808 4140
rect 12763 4100 12808 4128
rect 12802 4088 12808 4100
rect 12860 4128 12866 4140
rect 13906 4128 13912 4140
rect 12860 4100 13912 4128
rect 12860 4088 12866 4100
rect 13906 4088 13912 4100
rect 13964 4088 13970 4140
rect 14093 4131 14151 4137
rect 14093 4097 14105 4131
rect 14139 4128 14151 4131
rect 14550 4128 14556 4140
rect 14139 4100 14556 4128
rect 14139 4097 14151 4100
rect 14093 4091 14151 4097
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 15838 4088 15844 4140
rect 15896 4128 15902 4140
rect 16758 4128 16764 4140
rect 15896 4100 16764 4128
rect 15896 4088 15902 4100
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 17865 4131 17923 4137
rect 17865 4097 17877 4131
rect 17911 4128 17923 4131
rect 18690 4128 18696 4140
rect 17911 4100 18696 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 18969 4131 19027 4137
rect 18969 4097 18981 4131
rect 19015 4128 19027 4131
rect 19058 4128 19064 4140
rect 19015 4100 19064 4128
rect 19015 4097 19027 4100
rect 18969 4091 19027 4097
rect 19058 4088 19064 4100
rect 19116 4088 19122 4140
rect 19242 4088 19248 4140
rect 19300 4128 19306 4140
rect 20165 4131 20223 4137
rect 20165 4128 20177 4131
rect 19300 4100 20177 4128
rect 19300 4088 19306 4100
rect 20165 4097 20177 4100
rect 20211 4128 20223 4131
rect 20211 4100 21036 4128
rect 20211 4097 20223 4100
rect 20165 4091 20223 4097
rect 8573 4063 8631 4069
rect 8573 4060 8585 4063
rect 7760 4032 8585 4060
rect 8573 4029 8585 4032
rect 8619 4060 8631 4063
rect 8619 4032 9444 4060
rect 8619 4029 8631 4032
rect 8573 4023 8631 4029
rect 3510 3952 3516 4004
rect 3568 3992 3574 4004
rect 6546 3992 6552 4004
rect 3568 3964 6552 3992
rect 3568 3952 3574 3964
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 6822 3952 6828 4004
rect 6880 3992 6886 4004
rect 8941 3995 8999 4001
rect 8941 3992 8953 3995
rect 6880 3964 8953 3992
rect 6880 3952 6886 3964
rect 8941 3961 8953 3964
rect 8987 3992 8999 3995
rect 9122 3992 9128 4004
rect 8987 3964 9128 3992
rect 8987 3961 8999 3964
rect 8941 3955 8999 3961
rect 9122 3952 9128 3964
rect 9180 3952 9186 4004
rect 9416 3933 9444 4032
rect 9490 4020 9496 4072
rect 9548 4060 9554 4072
rect 10134 4060 10140 4072
rect 9548 4032 9593 4060
rect 10095 4032 10140 4060
rect 9548 4020 9554 4032
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 10502 4060 10508 4072
rect 10415 4032 10508 4060
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 10870 4060 10876 4072
rect 10831 4032 10876 4060
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 16390 4020 16396 4072
rect 16448 4060 16454 4072
rect 21008 4069 21036 4100
rect 21450 4088 21456 4140
rect 21508 4128 21514 4140
rect 22554 4128 22560 4140
rect 21508 4100 22560 4128
rect 21508 4088 21514 4100
rect 22554 4088 22560 4100
rect 22612 4088 22618 4140
rect 25498 4128 25504 4140
rect 25411 4100 25504 4128
rect 25498 4088 25504 4100
rect 25556 4128 25562 4140
rect 27062 4128 27068 4140
rect 25556 4100 27068 4128
rect 25556 4088 25562 4100
rect 27062 4088 27068 4100
rect 27120 4088 27126 4140
rect 20717 4063 20775 4069
rect 20717 4060 20729 4063
rect 16448 4032 20729 4060
rect 16448 4020 16454 4032
rect 20717 4029 20729 4032
rect 20763 4029 20775 4063
rect 20717 4023 20775 4029
rect 20993 4063 21051 4069
rect 20993 4029 21005 4063
rect 21039 4029 21051 4063
rect 20993 4023 21051 4029
rect 22005 4063 22063 4069
rect 22005 4029 22017 4063
rect 22051 4060 22063 4063
rect 22316 4063 22374 4069
rect 22316 4060 22328 4063
rect 22051 4032 22328 4060
rect 22051 4029 22063 4032
rect 22005 4023 22063 4029
rect 22316 4029 22328 4032
rect 22362 4029 22374 4063
rect 22316 4023 22374 4029
rect 24648 4063 24706 4069
rect 24648 4029 24660 4063
rect 24694 4060 24706 4063
rect 25130 4060 25136 4072
rect 24694 4032 25136 4060
rect 24694 4029 24706 4032
rect 24648 4023 24706 4029
rect 25130 4020 25136 4032
rect 25188 4020 25194 4072
rect 25660 4063 25718 4069
rect 25660 4029 25672 4063
rect 25706 4060 25718 4063
rect 25866 4060 25872 4072
rect 25706 4032 25872 4060
rect 25706 4029 25718 4032
rect 25660 4023 25718 4029
rect 25866 4020 25872 4032
rect 25924 4060 25930 4072
rect 26053 4063 26111 4069
rect 26053 4060 26065 4063
rect 25924 4032 26065 4060
rect 25924 4020 25930 4032
rect 26053 4029 26065 4032
rect 26099 4029 26111 4063
rect 26053 4023 26111 4029
rect 9401 3927 9459 3933
rect 9401 3893 9413 3927
rect 9447 3924 9459 3927
rect 9858 3924 9864 3936
rect 9447 3896 9864 3924
rect 9447 3893 9459 3896
rect 9401 3887 9459 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 10520 3924 10548 4020
rect 10965 3995 11023 4001
rect 10965 3961 10977 3995
rect 11011 3992 11023 3995
rect 12342 3992 12348 4004
rect 11011 3964 12348 3992
rect 11011 3961 11023 3964
rect 10965 3955 11023 3961
rect 12342 3952 12348 3964
rect 12400 3952 12406 4004
rect 12529 3995 12587 4001
rect 12529 3961 12541 3995
rect 12575 3961 12587 3995
rect 12529 3955 12587 3961
rect 10686 3924 10692 3936
rect 10520 3896 10692 3924
rect 10686 3884 10692 3896
rect 10744 3924 10750 3936
rect 11241 3927 11299 3933
rect 11241 3924 11253 3927
rect 10744 3896 11253 3924
rect 10744 3884 10750 3896
rect 11241 3893 11253 3896
rect 11287 3893 11299 3927
rect 11241 3887 11299 3893
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11609 3927 11667 3933
rect 11609 3924 11621 3927
rect 11480 3896 11621 3924
rect 11480 3884 11486 3896
rect 11609 3893 11621 3896
rect 11655 3893 11667 3927
rect 11609 3887 11667 3893
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12544 3924 12572 3955
rect 12618 3952 12624 4004
rect 12676 3992 12682 4004
rect 13909 3995 13967 4001
rect 12676 3964 12721 3992
rect 12676 3952 12682 3964
rect 13909 3961 13921 3995
rect 13955 3992 13967 3995
rect 14185 3995 14243 4001
rect 14185 3992 14197 3995
rect 13955 3964 14197 3992
rect 13955 3961 13967 3964
rect 13909 3955 13967 3961
rect 14185 3961 14197 3964
rect 14231 3992 14243 3995
rect 14366 3992 14372 4004
rect 14231 3964 14372 3992
rect 14231 3961 14243 3964
rect 14185 3955 14243 3961
rect 14366 3952 14372 3964
rect 14424 3952 14430 4004
rect 15105 3995 15163 4001
rect 15105 3961 15117 3995
rect 15151 3992 15163 3995
rect 15654 3992 15660 4004
rect 15151 3964 15660 3992
rect 15151 3961 15163 3964
rect 15105 3955 15163 3961
rect 15654 3952 15660 3964
rect 15712 3952 15718 4004
rect 15746 3952 15752 4004
rect 15804 3992 15810 4004
rect 15804 3964 15849 3992
rect 15804 3952 15810 3964
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 16301 3995 16359 4001
rect 16301 3992 16313 3995
rect 15988 3964 16313 3992
rect 15988 3952 15994 3964
rect 16301 3961 16313 3964
rect 16347 3961 16359 3995
rect 16301 3955 16359 3961
rect 18414 3952 18420 4004
rect 18472 3992 18478 4004
rect 18874 3992 18880 4004
rect 18472 3964 18880 3992
rect 18472 3952 18478 3964
rect 18874 3952 18880 3964
rect 18932 3952 18938 4004
rect 19150 3952 19156 4004
rect 19208 3992 19214 4004
rect 19290 3995 19348 4001
rect 19290 3992 19302 3995
rect 19208 3964 19302 3992
rect 19208 3952 19214 3964
rect 19290 3961 19302 3964
rect 19336 3961 19348 3995
rect 19290 3955 19348 3961
rect 12492 3896 12572 3924
rect 12492 3884 12498 3896
rect 17954 3884 17960 3936
rect 18012 3924 18018 3936
rect 18785 3927 18843 3933
rect 18785 3924 18797 3927
rect 18012 3896 18797 3924
rect 18012 3884 18018 3896
rect 18785 3893 18797 3896
rect 18831 3893 18843 3927
rect 18785 3887 18843 3893
rect 19889 3927 19947 3933
rect 19889 3893 19901 3927
rect 19935 3924 19947 3927
rect 19978 3924 19984 3936
rect 19935 3896 19984 3924
rect 19935 3893 19947 3896
rect 19889 3887 19947 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 22005 3927 22063 3933
rect 22005 3924 22017 3927
rect 20680 3896 22017 3924
rect 20680 3884 20686 3896
rect 22005 3893 22017 3896
rect 22051 3924 22063 3927
rect 22097 3927 22155 3933
rect 22097 3924 22109 3927
rect 22051 3896 22109 3924
rect 22051 3893 22063 3896
rect 22005 3887 22063 3893
rect 22097 3893 22109 3896
rect 22143 3893 22155 3927
rect 22097 3887 22155 3893
rect 22186 3884 22192 3936
rect 22244 3924 22250 3936
rect 22419 3927 22477 3933
rect 22419 3924 22431 3927
rect 22244 3896 22431 3924
rect 22244 3884 22250 3896
rect 22419 3893 22431 3896
rect 22465 3893 22477 3927
rect 22419 3887 22477 3893
rect 25498 3884 25504 3936
rect 25556 3924 25562 3936
rect 25731 3927 25789 3933
rect 25731 3924 25743 3927
rect 25556 3896 25743 3924
rect 25556 3884 25562 3896
rect 25731 3893 25743 3896
rect 25777 3893 25789 3927
rect 25731 3887 25789 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 7745 3723 7803 3729
rect 7745 3689 7757 3723
rect 7791 3720 7803 3723
rect 7926 3720 7932 3732
rect 7791 3692 7932 3720
rect 7791 3689 7803 3692
rect 7745 3683 7803 3689
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 10870 3720 10876 3732
rect 9916 3692 10876 3720
rect 9916 3680 9922 3692
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 16761 3723 16819 3729
rect 16761 3720 16773 3723
rect 12492 3692 16773 3720
rect 12492 3680 12498 3692
rect 16761 3689 16773 3692
rect 16807 3689 16819 3723
rect 17954 3720 17960 3732
rect 17915 3692 17960 3720
rect 16761 3683 16819 3689
rect 17954 3680 17960 3692
rect 18012 3680 18018 3732
rect 19058 3720 19064 3732
rect 19019 3692 19064 3720
rect 19058 3680 19064 3692
rect 19116 3680 19122 3732
rect 19981 3723 20039 3729
rect 19981 3689 19993 3723
rect 20027 3720 20039 3723
rect 22186 3720 22192 3732
rect 20027 3692 22192 3720
rect 20027 3689 20039 3692
rect 19981 3683 20039 3689
rect 9033 3655 9091 3661
rect 9033 3621 9045 3655
rect 9079 3652 9091 3655
rect 9398 3652 9404 3664
rect 9079 3624 9404 3652
rect 9079 3621 9091 3624
rect 9033 3615 9091 3621
rect 9398 3612 9404 3624
rect 9456 3652 9462 3664
rect 13722 3652 13728 3664
rect 9456 3624 10640 3652
rect 13683 3624 13728 3652
rect 9456 3612 9462 3624
rect 10612 3596 10640 3624
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 15470 3652 15476 3664
rect 14384 3624 15476 3652
rect 6270 3544 6276 3596
rect 6328 3584 6334 3596
rect 6917 3587 6975 3593
rect 6917 3584 6929 3587
rect 6328 3556 6929 3584
rect 6328 3544 6334 3556
rect 6917 3553 6929 3556
rect 6963 3584 6975 3587
rect 7006 3584 7012 3596
rect 6963 3556 7012 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 8938 3584 8944 3596
rect 8251 3556 8944 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 9306 3544 9312 3596
rect 9364 3584 9370 3596
rect 9490 3584 9496 3596
rect 9364 3556 9496 3584
rect 9364 3544 9370 3556
rect 9490 3544 9496 3556
rect 9548 3584 9554 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9548 3556 9689 3584
rect 9548 3544 9554 3556
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 10134 3544 10140 3596
rect 10192 3584 10198 3596
rect 10413 3587 10471 3593
rect 10413 3584 10425 3587
rect 10192 3556 10425 3584
rect 10192 3544 10198 3556
rect 10413 3553 10425 3556
rect 10459 3553 10471 3587
rect 10594 3584 10600 3596
rect 10555 3556 10600 3584
rect 10413 3547 10471 3553
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3516 5963 3519
rect 10042 3516 10048 3528
rect 5951 3488 10048 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 10428 3516 10456 3547
rect 10594 3544 10600 3556
rect 10652 3544 10658 3596
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3584 11115 3587
rect 11422 3584 11428 3596
rect 11103 3556 11428 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 11422 3544 11428 3556
rect 11480 3544 11486 3596
rect 11974 3584 11980 3596
rect 11935 3556 11980 3584
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 13449 3587 13507 3593
rect 13449 3584 13461 3587
rect 12400 3556 13461 3584
rect 12400 3544 12406 3556
rect 13449 3553 13461 3556
rect 13495 3584 13507 3587
rect 14182 3584 14188 3596
rect 13495 3556 14188 3584
rect 13495 3553 13507 3556
rect 13449 3547 13507 3553
rect 14182 3544 14188 3556
rect 14240 3544 14246 3596
rect 14384 3593 14412 3624
rect 15470 3612 15476 3624
rect 15528 3612 15534 3664
rect 16022 3652 16028 3664
rect 15983 3624 16028 3652
rect 16022 3612 16028 3624
rect 16080 3612 16086 3664
rect 19518 3652 19524 3664
rect 16132 3624 19524 3652
rect 14369 3587 14427 3593
rect 14369 3553 14381 3587
rect 14415 3553 14427 3587
rect 14369 3547 14427 3553
rect 11146 3516 11152 3528
rect 10428 3488 10732 3516
rect 11107 3488 11152 3516
rect 7101 3451 7159 3457
rect 7101 3417 7113 3451
rect 7147 3448 7159 3451
rect 8202 3448 8208 3460
rect 7147 3420 8208 3448
rect 7147 3417 7159 3420
rect 7101 3411 7159 3417
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 10704 3448 10732 3488
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 12250 3476 12256 3528
rect 12308 3516 12314 3528
rect 15381 3519 15439 3525
rect 12308 3488 12940 3516
rect 12308 3476 12314 3488
rect 12161 3451 12219 3457
rect 10704 3420 11652 3448
rect 11624 3392 11652 3420
rect 12161 3417 12173 3451
rect 12207 3448 12219 3451
rect 12710 3448 12716 3460
rect 12207 3420 12716 3448
rect 12207 3417 12219 3420
rect 12161 3411 12219 3417
rect 12710 3408 12716 3420
rect 12768 3408 12774 3460
rect 12912 3392 12940 3488
rect 15381 3485 15393 3519
rect 15427 3485 15439 3519
rect 15381 3479 15439 3485
rect 15396 3448 15424 3479
rect 15654 3476 15660 3528
rect 15712 3516 15718 3528
rect 16132 3516 16160 3624
rect 19518 3612 19524 3624
rect 19576 3612 19582 3664
rect 19337 3587 19395 3593
rect 19337 3553 19349 3587
rect 19383 3584 19395 3587
rect 19996 3584 20024 3683
rect 22186 3680 22192 3692
rect 22244 3680 22250 3732
rect 22278 3680 22284 3732
rect 22336 3720 22342 3732
rect 24627 3723 24685 3729
rect 24627 3720 24639 3723
rect 22336 3692 24639 3720
rect 22336 3680 22342 3692
rect 24627 3689 24639 3692
rect 24673 3689 24685 3723
rect 24627 3683 24685 3689
rect 20717 3655 20775 3661
rect 20717 3621 20729 3655
rect 20763 3652 20775 3655
rect 20990 3652 20996 3664
rect 20763 3624 20996 3652
rect 20763 3621 20775 3624
rect 20717 3615 20775 3621
rect 20990 3612 20996 3624
rect 21048 3612 21054 3664
rect 21085 3655 21143 3661
rect 21085 3621 21097 3655
rect 21131 3652 21143 3655
rect 21174 3652 21180 3664
rect 21131 3624 21180 3652
rect 21131 3621 21143 3624
rect 21085 3615 21143 3621
rect 21174 3612 21180 3624
rect 21232 3612 21238 3664
rect 21726 3612 21732 3664
rect 21784 3652 21790 3664
rect 22005 3655 22063 3661
rect 22005 3652 22017 3655
rect 21784 3624 22017 3652
rect 21784 3612 21790 3624
rect 22005 3621 22017 3624
rect 22051 3652 22063 3655
rect 25498 3652 25504 3664
rect 22051 3624 25504 3652
rect 22051 3621 22063 3624
rect 22005 3615 22063 3621
rect 25498 3612 25504 3624
rect 25556 3612 25562 3664
rect 22462 3584 22468 3596
rect 19383 3556 20024 3584
rect 22423 3556 22468 3584
rect 19383 3553 19395 3556
rect 19337 3547 19395 3553
rect 22462 3544 22468 3556
rect 22520 3544 22526 3596
rect 23544 3587 23602 3593
rect 23544 3553 23556 3587
rect 23590 3584 23602 3587
rect 24118 3584 24124 3596
rect 23590 3556 24124 3584
rect 23590 3553 23602 3556
rect 23544 3547 23602 3553
rect 24118 3544 24124 3556
rect 24176 3544 24182 3596
rect 24556 3587 24614 3593
rect 24556 3553 24568 3587
rect 24602 3584 24614 3587
rect 24670 3584 24676 3596
rect 24602 3556 24676 3584
rect 24602 3553 24614 3556
rect 24556 3547 24614 3553
rect 24670 3544 24676 3556
rect 24728 3544 24734 3596
rect 17586 3516 17592 3528
rect 15712 3488 16160 3516
rect 17499 3488 17592 3516
rect 15712 3476 15718 3488
rect 17586 3476 17592 3488
rect 17644 3516 17650 3528
rect 21450 3516 21456 3528
rect 17644 3488 21456 3516
rect 17644 3476 17650 3488
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 21637 3519 21695 3525
rect 21637 3485 21649 3519
rect 21683 3516 21695 3519
rect 21818 3516 21824 3528
rect 21683 3488 21824 3516
rect 21683 3485 21695 3488
rect 21637 3479 21695 3485
rect 21818 3476 21824 3488
rect 21876 3476 21882 3528
rect 15930 3448 15936 3460
rect 15396 3420 15936 3448
rect 15930 3408 15936 3420
rect 15988 3448 15994 3460
rect 15988 3420 19656 3448
rect 15988 3408 15994 3420
rect 8018 3380 8024 3392
rect 7979 3352 8024 3380
rect 8018 3340 8024 3352
rect 8076 3380 8082 3392
rect 8294 3380 8300 3392
rect 8076 3352 8300 3380
rect 8076 3340 8082 3352
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 8389 3383 8447 3389
rect 8389 3349 8401 3383
rect 8435 3380 8447 3383
rect 8846 3380 8852 3392
rect 8435 3352 8852 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 11425 3383 11483 3389
rect 11425 3380 11437 3383
rect 9364 3352 11437 3380
rect 9364 3340 9370 3352
rect 11425 3349 11437 3352
rect 11471 3380 11483 3383
rect 11514 3380 11520 3392
rect 11471 3352 11520 3380
rect 11471 3349 11483 3352
rect 11425 3343 11483 3349
rect 11514 3340 11520 3352
rect 11572 3340 11578 3392
rect 11606 3340 11612 3392
rect 11664 3380 11670 3392
rect 11793 3383 11851 3389
rect 11793 3380 11805 3383
rect 11664 3352 11805 3380
rect 11664 3340 11670 3352
rect 11793 3349 11805 3352
rect 11839 3349 11851 3383
rect 12618 3380 12624 3392
rect 12579 3352 12624 3380
rect 11793 3343 11851 3349
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 12894 3380 12900 3392
rect 12855 3352 12900 3380
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13262 3380 13268 3392
rect 13223 3352 13268 3380
rect 13262 3340 13268 3352
rect 13320 3340 13326 3392
rect 14642 3380 14648 3392
rect 14603 3352 14648 3380
rect 14642 3340 14648 3352
rect 14700 3340 14706 3392
rect 15105 3383 15163 3389
rect 15105 3349 15117 3383
rect 15151 3380 15163 3383
rect 15286 3380 15292 3392
rect 15151 3352 15292 3380
rect 15151 3349 15163 3352
rect 15105 3343 15163 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 16485 3383 16543 3389
rect 16485 3349 16497 3383
rect 16531 3380 16543 3383
rect 16574 3380 16580 3392
rect 16531 3352 16580 3380
rect 16531 3349 16543 3352
rect 16485 3343 16543 3349
rect 16574 3340 16580 3352
rect 16632 3340 16638 3392
rect 18506 3380 18512 3392
rect 18467 3352 18512 3380
rect 18506 3340 18512 3352
rect 18564 3340 18570 3392
rect 19518 3380 19524 3392
rect 19479 3352 19524 3380
rect 19518 3340 19524 3352
rect 19576 3340 19582 3392
rect 19628 3380 19656 3420
rect 20346 3408 20352 3460
rect 20404 3448 20410 3460
rect 22603 3451 22661 3457
rect 22603 3448 22615 3451
rect 20404 3420 22615 3448
rect 20404 3408 20410 3420
rect 22603 3417 22615 3420
rect 22649 3417 22661 3451
rect 22603 3411 22661 3417
rect 23615 3383 23673 3389
rect 23615 3380 23627 3383
rect 19628 3352 23627 3380
rect 23615 3349 23627 3352
rect 23661 3349 23673 3383
rect 23615 3343 23673 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 7006 3176 7012 3188
rect 6967 3148 7012 3176
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 8849 3179 8907 3185
rect 8849 3145 8861 3179
rect 8895 3176 8907 3179
rect 8938 3176 8944 3188
rect 8895 3148 8944 3176
rect 8895 3145 8907 3148
rect 8849 3139 8907 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9217 3179 9275 3185
rect 9217 3145 9229 3179
rect 9263 3176 9275 3179
rect 9858 3176 9864 3188
rect 9263 3148 9864 3176
rect 9263 3145 9275 3148
rect 9217 3139 9275 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 11422 3176 11428 3188
rect 11383 3148 11428 3176
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 11974 3176 11980 3188
rect 11935 3148 11980 3176
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 15470 3176 15476 3188
rect 15431 3148 15476 3176
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 15930 3176 15936 3188
rect 15891 3148 15936 3176
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 16758 3136 16764 3188
rect 16816 3176 16822 3188
rect 17589 3179 17647 3185
rect 17589 3176 17601 3179
rect 16816 3148 17601 3176
rect 16816 3136 16822 3148
rect 17589 3145 17601 3148
rect 17635 3176 17647 3179
rect 17954 3176 17960 3188
rect 17635 3148 17960 3176
rect 17635 3145 17647 3148
rect 17589 3139 17647 3145
rect 17954 3136 17960 3148
rect 18012 3136 18018 3188
rect 18417 3179 18475 3185
rect 18417 3145 18429 3179
rect 18463 3176 18475 3179
rect 18506 3176 18512 3188
rect 18463 3148 18512 3176
rect 18463 3145 18475 3148
rect 18417 3139 18475 3145
rect 18506 3136 18512 3148
rect 18564 3136 18570 3188
rect 19978 3176 19984 3188
rect 19939 3148 19984 3176
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 21542 3176 21548 3188
rect 21503 3148 21548 3176
rect 21542 3136 21548 3148
rect 21600 3136 21606 3188
rect 23198 3136 23204 3188
rect 23256 3176 23262 3188
rect 24811 3179 24869 3185
rect 24811 3176 24823 3179
rect 23256 3148 24823 3176
rect 23256 3136 23262 3148
rect 24811 3145 24823 3148
rect 24857 3145 24869 3179
rect 24811 3139 24869 3145
rect 6273 3111 6331 3117
rect 6273 3077 6285 3111
rect 6319 3108 6331 3111
rect 7190 3108 7196 3120
rect 6319 3080 7196 3108
rect 6319 3077 6331 3080
rect 6273 3071 6331 3077
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3040 4767 3043
rect 6178 3040 6184 3052
rect 4755 3012 6184 3040
rect 4755 3009 4767 3012
rect 4709 3003 4767 3009
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 5788 2975 5846 2981
rect 5788 2941 5800 2975
rect 5834 2972 5846 2975
rect 6288 2972 6316 3071
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 13357 3111 13415 3117
rect 13357 3108 13369 3111
rect 7852 3080 13369 3108
rect 7852 2981 7880 3080
rect 13357 3077 13369 3080
rect 13403 3108 13415 3111
rect 15194 3108 15200 3120
rect 13403 3080 15200 3108
rect 13403 3077 13415 3080
rect 13357 3071 13415 3077
rect 15194 3068 15200 3080
rect 15252 3068 15258 3120
rect 16850 3108 16856 3120
rect 15488 3080 16856 3108
rect 9122 3000 9128 3052
rect 9180 3040 9186 3052
rect 10594 3040 10600 3052
rect 9180 3012 9674 3040
rect 9180 3000 9186 3012
rect 5834 2944 6316 2972
rect 6641 2975 6699 2981
rect 5834 2941 5846 2944
rect 5788 2935 5846 2941
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 7837 2975 7895 2981
rect 7837 2972 7849 2975
rect 6687 2944 7849 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 7837 2941 7849 2944
rect 7883 2941 7895 2975
rect 9306 2972 9312 2984
rect 9219 2944 9312 2972
rect 7837 2935 7895 2941
rect 9306 2932 9312 2944
rect 9364 2932 9370 2984
rect 8478 2904 8484 2916
rect 8439 2876 8484 2904
rect 8478 2864 8484 2876
rect 8536 2864 8542 2916
rect 5859 2839 5917 2845
rect 5859 2805 5871 2839
rect 5905 2836 5917 2839
rect 7466 2836 7472 2848
rect 5905 2808 7472 2836
rect 5905 2805 5917 2808
rect 5859 2799 5917 2805
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 7653 2839 7711 2845
rect 7653 2805 7665 2839
rect 7699 2836 7711 2839
rect 7926 2836 7932 2848
rect 7699 2808 7932 2836
rect 7699 2805 7711 2808
rect 7653 2799 7711 2805
rect 7926 2796 7932 2808
rect 7984 2836 7990 2848
rect 9324 2836 9352 2932
rect 9646 2904 9674 3012
rect 10336 3012 10600 3040
rect 10336 2981 10364 3012
rect 10594 3000 10600 3012
rect 10652 3040 10658 3052
rect 11057 3043 11115 3049
rect 11057 3040 11069 3043
rect 10652 3012 11069 3040
rect 10652 3000 10658 3012
rect 11057 3009 11069 3012
rect 11103 3009 11115 3043
rect 11057 3003 11115 3009
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 11204 3012 13814 3040
rect 11204 3000 11210 3012
rect 9861 2975 9919 2981
rect 9861 2941 9873 2975
rect 9907 2941 9919 2975
rect 9861 2935 9919 2941
rect 10321 2975 10379 2981
rect 10321 2941 10333 2975
rect 10367 2941 10379 2975
rect 10321 2935 10379 2941
rect 10689 2975 10747 2981
rect 10689 2941 10701 2975
rect 10735 2972 10747 2975
rect 10870 2972 10876 2984
rect 10735 2944 10876 2972
rect 10735 2941 10747 2944
rect 10689 2935 10747 2941
rect 9876 2904 9904 2935
rect 10870 2932 10876 2944
rect 10928 2932 10934 2984
rect 11238 2932 11244 2984
rect 11296 2972 11302 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 11296 2944 12449 2972
rect 11296 2932 11302 2944
rect 12437 2941 12449 2944
rect 12483 2972 12495 2975
rect 13262 2972 13268 2984
rect 12483 2944 13268 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 13786 2972 13814 3012
rect 14274 2972 14280 2984
rect 13786 2944 14280 2972
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 14366 2932 14372 2984
rect 14424 2972 14430 2984
rect 15197 2975 15255 2981
rect 15197 2972 15209 2975
rect 14424 2944 15209 2972
rect 14424 2932 14430 2944
rect 15197 2941 15209 2944
rect 15243 2972 15255 2975
rect 15488 2972 15516 3080
rect 16850 3068 16856 3080
rect 16908 3068 16914 3120
rect 19153 3111 19211 3117
rect 19153 3077 19165 3111
rect 19199 3108 19211 3111
rect 20622 3108 20628 3120
rect 19199 3080 20628 3108
rect 19199 3077 19211 3080
rect 19153 3071 19211 3077
rect 16485 3043 16543 3049
rect 16485 3009 16497 3043
rect 16531 3040 16543 3043
rect 16574 3040 16580 3052
rect 16531 3012 16580 3040
rect 16531 3009 16543 3012
rect 16485 3003 16543 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 17129 3043 17187 3049
rect 17129 3009 17141 3043
rect 17175 3040 17187 3043
rect 18414 3040 18420 3052
rect 17175 3012 18420 3040
rect 17175 3009 17187 3012
rect 17129 3003 17187 3009
rect 18414 3000 18420 3012
rect 18472 3040 18478 3052
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 18472 3012 18613 3040
rect 18472 3000 18478 3012
rect 18601 3009 18613 3012
rect 18647 3040 18659 3043
rect 19242 3040 19248 3052
rect 18647 3012 19248 3040
rect 18647 3009 18659 3012
rect 18601 3003 18659 3009
rect 19242 3000 19248 3012
rect 19300 3040 19306 3052
rect 20456 3049 20484 3080
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 21082 3068 21088 3120
rect 21140 3108 21146 3120
rect 22462 3108 22468 3120
rect 21140 3080 22468 3108
rect 21140 3068 21146 3080
rect 22462 3068 22468 3080
rect 22520 3108 22526 3120
rect 22649 3111 22707 3117
rect 22649 3108 22661 3111
rect 22520 3080 22661 3108
rect 22520 3068 22526 3080
rect 22649 3077 22661 3080
rect 22695 3077 22707 3111
rect 24118 3108 24124 3120
rect 24079 3080 24124 3108
rect 22649 3071 22707 3077
rect 24118 3068 24124 3080
rect 24176 3068 24182 3120
rect 19521 3043 19579 3049
rect 19521 3040 19533 3043
rect 19300 3012 19533 3040
rect 19300 3000 19306 3012
rect 19521 3009 19533 3012
rect 19567 3009 19579 3043
rect 19521 3003 19579 3009
rect 20441 3043 20499 3049
rect 20441 3009 20453 3043
rect 20487 3009 20499 3043
rect 21726 3040 21732 3052
rect 21687 3012 21732 3040
rect 20441 3003 20499 3009
rect 21726 3000 21732 3012
rect 21784 3000 21790 3052
rect 21818 3000 21824 3052
rect 21876 3040 21882 3052
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 21876 3012 22017 3040
rect 21876 3000 21882 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 15243 2944 15516 2972
rect 15243 2941 15255 2944
rect 15197 2935 15255 2941
rect 22370 2932 22376 2984
rect 22428 2972 22434 2984
rect 23385 2975 23443 2981
rect 23385 2972 23397 2975
rect 22428 2944 23397 2972
rect 22428 2932 22434 2944
rect 23385 2941 23397 2944
rect 23431 2972 23443 2975
rect 23569 2975 23627 2981
rect 23569 2972 23581 2975
rect 23431 2944 23581 2972
rect 23431 2941 23443 2944
rect 23385 2935 23443 2941
rect 23569 2941 23581 2944
rect 23615 2941 23627 2975
rect 23569 2935 23627 2941
rect 24740 2975 24798 2981
rect 24740 2941 24752 2975
rect 24786 2972 24798 2975
rect 24854 2972 24860 2984
rect 24786 2944 24860 2972
rect 24786 2941 24798 2944
rect 24740 2935 24798 2941
rect 24854 2932 24860 2944
rect 24912 2972 24918 2984
rect 25133 2975 25191 2981
rect 25133 2972 25145 2975
rect 24912 2944 25145 2972
rect 24912 2932 24918 2944
rect 25133 2941 25145 2944
rect 25179 2941 25191 2975
rect 25133 2935 25191 2941
rect 10778 2904 10784 2916
rect 9646 2876 9904 2904
rect 10739 2876 10784 2904
rect 10778 2864 10784 2876
rect 10836 2864 10842 2916
rect 11422 2864 11428 2916
rect 11480 2904 11486 2916
rect 11790 2904 11796 2916
rect 11480 2876 11796 2904
rect 11480 2864 11486 2876
rect 11790 2864 11796 2876
rect 11848 2904 11854 2916
rect 12618 2904 12624 2916
rect 11848 2876 12624 2904
rect 11848 2864 11854 2876
rect 12618 2864 12624 2876
rect 12676 2904 12682 2916
rect 12758 2907 12816 2913
rect 12758 2904 12770 2907
rect 12676 2876 12770 2904
rect 12676 2864 12682 2876
rect 12758 2873 12770 2876
rect 12804 2904 12816 2907
rect 13633 2907 13691 2913
rect 13633 2904 13645 2907
rect 12804 2876 13645 2904
rect 12804 2873 12816 2876
rect 12758 2867 12816 2873
rect 13633 2873 13645 2876
rect 13679 2904 13691 2907
rect 13722 2904 13728 2916
rect 13679 2876 13728 2904
rect 13679 2873 13691 2876
rect 13633 2867 13691 2873
rect 13722 2864 13728 2876
rect 13780 2904 13786 2916
rect 14093 2907 14151 2913
rect 14093 2904 14105 2907
rect 13780 2876 14105 2904
rect 13780 2864 13786 2876
rect 14093 2873 14105 2876
rect 14139 2904 14151 2907
rect 14598 2907 14656 2913
rect 14598 2904 14610 2907
rect 14139 2876 14610 2904
rect 14139 2873 14151 2876
rect 14093 2867 14151 2873
rect 14598 2873 14610 2876
rect 14644 2873 14656 2907
rect 14598 2867 14656 2873
rect 16301 2907 16359 2913
rect 16301 2873 16313 2907
rect 16347 2904 16359 2907
rect 16577 2907 16635 2913
rect 16577 2904 16589 2907
rect 16347 2876 16589 2904
rect 16347 2873 16359 2876
rect 16301 2867 16359 2873
rect 16577 2873 16589 2876
rect 16623 2904 16635 2907
rect 17770 2904 17776 2916
rect 16623 2876 17776 2904
rect 16623 2873 16635 2876
rect 16577 2867 16635 2873
rect 17770 2864 17776 2876
rect 17828 2864 17834 2916
rect 18693 2907 18751 2913
rect 18693 2873 18705 2907
rect 18739 2873 18751 2907
rect 20162 2904 20168 2916
rect 20123 2876 20168 2904
rect 18693 2867 18751 2873
rect 7984 2808 9352 2836
rect 7984 2796 7990 2808
rect 18506 2796 18512 2848
rect 18564 2836 18570 2848
rect 18708 2836 18736 2867
rect 20162 2864 20168 2876
rect 20220 2864 20226 2916
rect 20257 2907 20315 2913
rect 20257 2873 20269 2907
rect 20303 2873 20315 2907
rect 20257 2867 20315 2873
rect 21821 2907 21879 2913
rect 21821 2873 21833 2907
rect 21867 2873 21879 2907
rect 21821 2867 21879 2873
rect 18564 2808 18736 2836
rect 18564 2796 18570 2808
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 20272 2836 20300 2867
rect 20036 2808 20300 2836
rect 20036 2796 20042 2808
rect 20530 2796 20536 2848
rect 20588 2836 20594 2848
rect 21085 2839 21143 2845
rect 21085 2836 21097 2839
rect 20588 2808 21097 2836
rect 20588 2796 20594 2808
rect 21085 2805 21097 2808
rect 21131 2836 21143 2839
rect 21174 2836 21180 2848
rect 21131 2808 21180 2836
rect 21131 2805 21143 2808
rect 21085 2799 21143 2805
rect 21174 2796 21180 2808
rect 21232 2796 21238 2848
rect 21542 2796 21548 2848
rect 21600 2836 21606 2848
rect 21836 2836 21864 2867
rect 21600 2808 21864 2836
rect 21600 2796 21606 2808
rect 23566 2796 23572 2848
rect 23624 2836 23630 2848
rect 23799 2839 23857 2845
rect 23799 2836 23811 2839
rect 23624 2808 23811 2836
rect 23624 2796 23630 2808
rect 23799 2805 23811 2808
rect 23845 2805 23857 2839
rect 23799 2799 23857 2805
rect 24581 2839 24639 2845
rect 24581 2805 24593 2839
rect 24627 2836 24639 2839
rect 24670 2836 24676 2848
rect 24627 2808 24676 2836
rect 24627 2805 24639 2808
rect 24581 2799 24639 2805
rect 24670 2796 24676 2808
rect 24728 2836 24734 2848
rect 26142 2836 26148 2848
rect 24728 2808 26148 2836
rect 24728 2796 24734 2808
rect 26142 2796 26148 2808
rect 26200 2796 26206 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 5951 2635 6009 2641
rect 5951 2601 5963 2635
rect 5997 2632 6009 2635
rect 7742 2632 7748 2644
rect 5997 2604 7748 2632
rect 5997 2601 6009 2604
rect 5951 2595 6009 2601
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 7926 2632 7932 2644
rect 7887 2604 7932 2632
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 8478 2592 8484 2644
rect 8536 2632 8542 2644
rect 12989 2635 13047 2641
rect 12989 2632 13001 2635
rect 8536 2604 13001 2632
rect 8536 2592 8542 2604
rect 12989 2601 13001 2604
rect 13035 2632 13047 2635
rect 14182 2632 14188 2644
rect 13035 2604 13400 2632
rect 14143 2604 14188 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 6733 2567 6791 2573
rect 6733 2533 6745 2567
rect 6779 2564 6791 2567
rect 8849 2567 8907 2573
rect 6779 2536 8248 2564
rect 6779 2533 6791 2536
rect 6733 2527 6791 2533
rect 4868 2499 4926 2505
rect 4868 2465 4880 2499
rect 4914 2465 4926 2499
rect 4868 2459 4926 2465
rect 4883 2428 4911 2459
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 8220 2505 8248 2536
rect 8849 2533 8861 2567
rect 8895 2564 8907 2567
rect 9674 2564 9680 2576
rect 8895 2536 9680 2564
rect 8895 2533 8907 2536
rect 8849 2527 8907 2533
rect 9674 2524 9680 2536
rect 9732 2524 9738 2576
rect 10642 2567 10700 2573
rect 10642 2564 10654 2567
rect 10152 2536 10654 2564
rect 5848 2499 5906 2505
rect 5848 2496 5860 2499
rect 5592 2468 5860 2496
rect 5592 2456 5598 2468
rect 5848 2465 5860 2468
rect 5894 2496 5906 2499
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 5894 2468 6285 2496
rect 5894 2465 5906 2468
rect 5848 2459 5906 2465
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7377 2499 7435 2505
rect 7377 2496 7389 2499
rect 6963 2468 7389 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7377 2465 7389 2468
rect 7423 2465 7435 2499
rect 7377 2459 7435 2465
rect 8205 2499 8263 2505
rect 8205 2465 8217 2499
rect 8251 2496 8263 2499
rect 9030 2496 9036 2508
rect 8251 2468 9036 2496
rect 8251 2465 8263 2468
rect 8205 2459 8263 2465
rect 9030 2456 9036 2468
rect 9088 2456 9094 2508
rect 9122 2456 9128 2508
rect 9180 2496 9186 2508
rect 9309 2499 9367 2505
rect 9309 2496 9321 2499
rect 9180 2468 9321 2496
rect 9180 2456 9186 2468
rect 9309 2465 9321 2468
rect 9355 2465 9367 2499
rect 9309 2459 9367 2465
rect 9398 2456 9404 2508
rect 9456 2496 9462 2508
rect 10152 2505 10180 2536
rect 10642 2533 10654 2536
rect 10688 2564 10700 2567
rect 11422 2564 11428 2576
rect 10688 2536 11428 2564
rect 10688 2533 10700 2536
rect 10642 2527 10700 2533
rect 11422 2524 11428 2536
rect 11480 2524 11486 2576
rect 11606 2564 11612 2576
rect 11567 2536 11612 2564
rect 11606 2524 11612 2536
rect 11664 2524 11670 2576
rect 13372 2573 13400 2604
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 14274 2592 14280 2644
rect 14332 2632 14338 2644
rect 14553 2635 14611 2641
rect 14553 2632 14565 2635
rect 14332 2604 14565 2632
rect 14332 2592 14338 2604
rect 14553 2601 14565 2604
rect 14599 2601 14611 2635
rect 15194 2632 15200 2644
rect 15155 2604 15200 2632
rect 14553 2595 14611 2601
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 17586 2632 17592 2644
rect 17547 2604 17592 2632
rect 17586 2592 17592 2604
rect 17644 2592 17650 2644
rect 18782 2632 18788 2644
rect 18743 2604 18788 2632
rect 18782 2592 18788 2604
rect 18840 2592 18846 2644
rect 20162 2632 20168 2644
rect 20123 2604 20168 2632
rect 20162 2592 20168 2604
rect 20220 2632 20226 2644
rect 21818 2632 21824 2644
rect 20220 2604 21824 2632
rect 20220 2592 20226 2604
rect 21818 2592 21824 2604
rect 21876 2592 21882 2644
rect 23385 2635 23443 2641
rect 23385 2601 23397 2635
rect 23431 2632 23443 2635
rect 23566 2632 23572 2644
rect 23431 2604 23572 2632
rect 23431 2601 23443 2604
rect 23385 2595 23443 2601
rect 13357 2567 13415 2573
rect 13357 2533 13369 2567
rect 13403 2533 13415 2567
rect 15212 2564 15240 2592
rect 15657 2567 15715 2573
rect 15657 2564 15669 2567
rect 15212 2536 15669 2564
rect 13357 2527 13415 2533
rect 15657 2533 15669 2536
rect 15703 2533 15715 2567
rect 15657 2527 15715 2533
rect 18141 2567 18199 2573
rect 18141 2533 18153 2567
rect 18187 2564 18199 2567
rect 19061 2567 19119 2573
rect 19061 2564 19073 2567
rect 18187 2536 19073 2564
rect 18187 2533 18199 2536
rect 18141 2527 18199 2533
rect 19061 2533 19073 2536
rect 19107 2564 19119 2567
rect 20530 2564 20536 2576
rect 19107 2536 20536 2564
rect 19107 2533 19119 2536
rect 19061 2527 19119 2533
rect 20530 2524 20536 2536
rect 20588 2524 20594 2576
rect 20625 2567 20683 2573
rect 20625 2533 20637 2567
rect 20671 2564 20683 2567
rect 21266 2564 21272 2576
rect 20671 2536 21272 2564
rect 20671 2533 20683 2536
rect 20625 2527 20683 2533
rect 21266 2524 21272 2536
rect 21324 2524 21330 2576
rect 21358 2524 21364 2576
rect 21416 2564 21422 2576
rect 21416 2536 21461 2564
rect 21416 2524 21422 2536
rect 10137 2499 10195 2505
rect 10137 2496 10149 2499
rect 9456 2468 10149 2496
rect 9456 2456 9462 2468
rect 10137 2465 10149 2468
rect 10183 2465 10195 2499
rect 10137 2459 10195 2465
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 10778 2496 10784 2508
rect 10367 2468 10784 2496
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 10778 2456 10784 2468
rect 10836 2496 10842 2508
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 10836 2468 11897 2496
rect 10836 2456 10842 2468
rect 11885 2465 11897 2468
rect 11931 2465 11943 2499
rect 11885 2459 11943 2465
rect 16850 2456 16856 2508
rect 16908 2496 16914 2508
rect 17037 2499 17095 2505
rect 17037 2496 17049 2499
rect 16908 2468 17049 2496
rect 16908 2456 16914 2468
rect 17037 2465 17049 2468
rect 17083 2465 17095 2499
rect 17037 2459 17095 2465
rect 22741 2499 22799 2505
rect 22741 2465 22753 2499
rect 22787 2496 22799 2499
rect 23400 2496 23428 2595
rect 23566 2592 23572 2604
rect 23624 2592 23630 2644
rect 23750 2592 23756 2644
rect 23808 2632 23814 2644
rect 25179 2635 25237 2641
rect 25179 2632 25191 2635
rect 23808 2604 25191 2632
rect 23808 2592 23814 2604
rect 25179 2601 25191 2604
rect 25225 2601 25237 2635
rect 25179 2595 25237 2601
rect 24026 2496 24032 2508
rect 24084 2505 24090 2508
rect 24084 2499 24122 2505
rect 22787 2468 23428 2496
rect 23974 2468 24032 2496
rect 22787 2465 22799 2468
rect 22741 2459 22799 2465
rect 24026 2456 24032 2468
rect 24110 2496 24122 2499
rect 24489 2499 24547 2505
rect 24489 2496 24501 2499
rect 24110 2468 24501 2496
rect 24110 2465 24122 2468
rect 24084 2459 24122 2465
rect 24489 2465 24501 2468
rect 24535 2465 24547 2499
rect 24489 2459 24547 2465
rect 25076 2499 25134 2505
rect 25076 2465 25088 2499
rect 25122 2465 25134 2499
rect 25076 2459 25134 2465
rect 24084 2456 24090 2459
rect 5353 2431 5411 2437
rect 5353 2428 5365 2431
rect 4883 2400 5365 2428
rect 5353 2397 5365 2400
rect 5399 2428 5411 2431
rect 10686 2428 10692 2440
rect 5399 2400 10692 2428
rect 5399 2397 5411 2400
rect 5353 2391 5411 2397
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 4939 2363 4997 2369
rect 4939 2329 4951 2363
rect 4985 2360 4997 2363
rect 5810 2360 5816 2372
rect 4985 2332 5816 2360
rect 4985 2329 4997 2332
rect 4939 2323 4997 2329
rect 5810 2320 5816 2332
rect 5868 2320 5874 2372
rect 7377 2363 7435 2369
rect 7377 2329 7389 2363
rect 7423 2360 7435 2363
rect 7561 2363 7619 2369
rect 7561 2360 7573 2363
rect 7423 2332 7573 2360
rect 7423 2329 7435 2332
rect 7377 2323 7435 2329
rect 7561 2329 7573 2332
rect 7607 2360 7619 2363
rect 8570 2360 8576 2372
rect 7607 2332 8576 2360
rect 7607 2329 7619 2332
rect 7561 2323 7619 2329
rect 8570 2320 8576 2332
rect 8628 2360 8634 2372
rect 9766 2360 9772 2372
rect 8628 2332 9772 2360
rect 8628 2320 8634 2332
rect 9766 2320 9772 2332
rect 9824 2320 9830 2372
rect 10042 2320 10048 2372
rect 10100 2360 10106 2372
rect 12345 2363 12403 2369
rect 12345 2360 12357 2363
rect 10100 2332 12357 2360
rect 10100 2320 10106 2332
rect 12345 2329 12357 2332
rect 12391 2360 12403 2363
rect 13280 2360 13308 2391
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 13964 2400 15577 2428
rect 13964 2388 13970 2400
rect 15565 2397 15577 2400
rect 15611 2428 15623 2431
rect 16485 2431 16543 2437
rect 16485 2428 16497 2431
rect 15611 2400 16497 2428
rect 15611 2397 15623 2400
rect 15565 2391 15623 2397
rect 16485 2397 16497 2400
rect 16531 2397 16543 2431
rect 16485 2391 16543 2397
rect 18782 2388 18788 2440
rect 18840 2428 18846 2440
rect 18969 2431 19027 2437
rect 18969 2428 18981 2431
rect 18840 2400 18981 2428
rect 18840 2388 18846 2400
rect 18969 2397 18981 2400
rect 19015 2397 19027 2431
rect 19242 2428 19248 2440
rect 19203 2400 19248 2428
rect 18969 2391 19027 2397
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2428 21051 2431
rect 21358 2428 21364 2440
rect 21039 2400 21364 2428
rect 21039 2397 21051 2400
rect 20993 2391 21051 2397
rect 21358 2388 21364 2400
rect 21416 2388 21422 2440
rect 21450 2388 21456 2440
rect 21508 2428 21514 2440
rect 24167 2431 24225 2437
rect 24167 2428 24179 2431
rect 21508 2400 24179 2428
rect 21508 2388 21514 2400
rect 24167 2397 24179 2400
rect 24213 2397 24225 2431
rect 24167 2391 24225 2397
rect 12391 2332 13308 2360
rect 13817 2363 13875 2369
rect 12391 2329 12403 2332
rect 12345 2323 12403 2329
rect 13817 2329 13829 2363
rect 13863 2360 13875 2363
rect 16114 2360 16120 2372
rect 13863 2332 16120 2360
rect 13863 2329 13875 2332
rect 13817 2323 13875 2329
rect 16114 2320 16120 2332
rect 16172 2320 16178 2372
rect 16758 2320 16764 2372
rect 16816 2360 16822 2372
rect 17221 2363 17279 2369
rect 17221 2360 17233 2363
rect 16816 2332 17233 2360
rect 16816 2320 16822 2332
rect 17221 2329 17233 2332
rect 17267 2329 17279 2363
rect 17221 2323 17279 2329
rect 19978 2320 19984 2372
rect 20036 2360 20042 2372
rect 21818 2360 21824 2372
rect 20036 2332 21128 2360
rect 21779 2332 21824 2360
rect 20036 2320 20042 2332
rect 7101 2295 7159 2301
rect 7101 2261 7113 2295
rect 7147 2292 7159 2295
rect 7282 2292 7288 2304
rect 7147 2264 7288 2292
rect 7147 2261 7159 2264
rect 7101 2255 7159 2261
rect 7282 2252 7288 2264
rect 7340 2252 7346 2304
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 11241 2295 11299 2301
rect 11241 2292 11253 2295
rect 9088 2264 11253 2292
rect 9088 2252 9094 2264
rect 11241 2261 11253 2264
rect 11287 2292 11299 2295
rect 12894 2292 12900 2304
rect 11287 2264 12900 2292
rect 11287 2261 11299 2264
rect 11241 2255 11299 2261
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 16850 2292 16856 2304
rect 16811 2264 16856 2292
rect 16850 2252 16856 2264
rect 16908 2252 16914 2304
rect 21100 2292 21128 2332
rect 21818 2320 21824 2332
rect 21876 2320 21882 2372
rect 22830 2320 22836 2372
rect 22888 2360 22894 2372
rect 25091 2360 25119 2459
rect 25501 2363 25559 2369
rect 25501 2360 25513 2363
rect 22888 2332 25513 2360
rect 22888 2320 22894 2332
rect 25501 2329 25513 2332
rect 25547 2329 25559 2363
rect 25501 2323 25559 2329
rect 22925 2295 22983 2301
rect 22925 2292 22937 2295
rect 21100 2264 22937 2292
rect 22925 2261 22937 2264
rect 22971 2261 22983 2295
rect 22925 2255 22983 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 1670 2048 1676 2100
rect 1728 2088 1734 2100
rect 6086 2088 6092 2100
rect 1728 2060 6092 2088
rect 1728 2048 1734 2060
rect 6086 2048 6092 2060
rect 6144 2088 6150 2100
rect 9398 2088 9404 2100
rect 6144 2060 9404 2088
rect 6144 2048 6150 2060
rect 9398 2048 9404 2060
rect 9456 2048 9462 2100
rect 2222 1980 2228 2032
rect 2280 2020 2286 2032
rect 6822 2020 6828 2032
rect 2280 1992 6828 2020
rect 2280 1980 2286 1992
rect 6822 1980 6828 1992
rect 6880 1980 6886 2032
rect 15838 76 15844 128
rect 15896 116 15902 128
rect 16482 116 16488 128
rect 15896 88 16488 116
rect 15896 76 15902 88
rect 16482 76 16488 88
rect 16540 76 16546 128
rect 13906 8 13912 60
rect 13964 48 13970 60
rect 19518 48 19524 60
rect 13964 20 19524 48
rect 13964 8 13970 20
rect 19518 8 19524 20
rect 19576 8 19582 60
<< via1 >>
rect 20 27480 72 27532
rect 664 27480 716 27532
rect 2780 27480 2832 27532
rect 3424 27480 3476 27532
rect 19524 27480 19576 27532
rect 21640 27480 21692 27532
rect 22468 27480 22520 27532
rect 23020 27480 23072 27532
rect 24860 27480 24912 27532
rect 25780 27480 25832 27532
rect 26240 27480 26292 27532
rect 27160 27480 27212 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 18788 24352 18840 24404
rect 10784 24216 10836 24268
rect 17592 24259 17644 24268
rect 17592 24225 17601 24259
rect 17601 24225 17635 24259
rect 17635 24225 17644 24259
rect 17592 24216 17644 24225
rect 23296 24216 23348 24268
rect 22928 24012 22980 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 6184 23808 6236 23860
rect 13176 23808 13228 23860
rect 14648 23808 14700 23860
rect 17408 23808 17460 23860
rect 17592 23851 17644 23860
rect 17592 23817 17601 23851
rect 17601 23817 17635 23851
rect 17635 23817 17644 23851
rect 17592 23808 17644 23817
rect 20168 23808 20220 23860
rect 23296 23851 23348 23860
rect 23296 23817 23305 23851
rect 23305 23817 23339 23851
rect 23339 23817 23348 23851
rect 23296 23808 23348 23817
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 8024 23672 8076 23724
rect 1216 23604 1268 23656
rect 4712 23647 4764 23656
rect 4712 23613 4721 23647
rect 4721 23613 4755 23647
rect 4755 23613 4764 23647
rect 4712 23604 4764 23613
rect 12440 23647 12492 23656
rect 4068 23468 4120 23520
rect 12440 23613 12449 23647
rect 12449 23613 12483 23647
rect 12483 23613 12492 23647
rect 12440 23604 12492 23613
rect 15936 23647 15988 23656
rect 7748 23468 7800 23520
rect 15936 23613 15945 23647
rect 15945 23613 15979 23647
rect 15979 23613 15988 23647
rect 15936 23604 15988 23613
rect 16948 23604 17000 23656
rect 17224 23604 17276 23656
rect 24216 23740 24268 23792
rect 25136 23604 25188 23656
rect 21456 23536 21508 23588
rect 22836 23536 22888 23588
rect 14832 23468 14884 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 112 23264 164 23316
rect 1400 23171 1452 23180
rect 1400 23137 1409 23171
rect 1409 23137 1443 23171
rect 1443 23137 1452 23171
rect 1400 23128 1452 23137
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 25136 22763 25188 22772
rect 25136 22729 25145 22763
rect 25145 22729 25179 22763
rect 25179 22729 25188 22763
rect 25136 22720 25188 22729
rect 11980 22652 12032 22704
rect 12440 22652 12492 22704
rect 1400 22516 1452 22568
rect 11980 22516 12032 22568
rect 25136 22516 25188 22568
rect 22008 22380 22060 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 24676 20952 24728 21004
rect 18604 20748 18656 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 24676 20587 24728 20596
rect 24676 20553 24685 20587
rect 24685 20553 24719 20587
rect 24719 20553 24728 20587
rect 24676 20544 24728 20553
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 12072 19864 12124 19916
rect 11612 19660 11664 19712
rect 13912 19703 13964 19712
rect 13912 19669 13921 19703
rect 13921 19669 13955 19703
rect 13955 19669 13964 19703
rect 13912 19660 13964 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 14832 19456 14884 19508
rect 11336 19363 11388 19372
rect 11336 19329 11345 19363
rect 11345 19329 11379 19363
rect 11379 19329 11388 19363
rect 11336 19320 11388 19329
rect 13912 19320 13964 19372
rect 17684 19320 17736 19372
rect 15844 19295 15896 19304
rect 8576 19184 8628 19236
rect 13544 19184 13596 19236
rect 15844 19261 15853 19295
rect 15853 19261 15887 19295
rect 15887 19261 15896 19295
rect 15844 19252 15896 19261
rect 10876 19116 10928 19168
rect 12072 19159 12124 19168
rect 12072 19125 12081 19159
rect 12081 19125 12115 19159
rect 12115 19125 12124 19159
rect 12072 19116 12124 19125
rect 12900 19116 12952 19168
rect 14832 19184 14884 19236
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 10876 18955 10928 18964
rect 10876 18921 10885 18955
rect 10885 18921 10919 18955
rect 10919 18921 10928 18955
rect 10876 18912 10928 18921
rect 12072 18912 12124 18964
rect 16764 18912 16816 18964
rect 9864 18887 9916 18896
rect 9864 18853 9873 18887
rect 9873 18853 9907 18887
rect 9907 18853 9916 18887
rect 9864 18844 9916 18853
rect 13728 18844 13780 18896
rect 15568 18887 15620 18896
rect 15568 18853 15577 18887
rect 15577 18853 15611 18887
rect 15611 18853 15620 18887
rect 15568 18844 15620 18853
rect 8576 18776 8628 18828
rect 11336 18776 11388 18828
rect 12164 18776 12216 18828
rect 21548 18819 21600 18828
rect 21548 18785 21566 18819
rect 21566 18785 21600 18819
rect 21548 18776 21600 18785
rect 22100 18776 22152 18828
rect 10232 18708 10284 18760
rect 11244 18751 11296 18760
rect 11244 18717 11253 18751
rect 11253 18717 11287 18751
rect 11287 18717 11296 18751
rect 11244 18708 11296 18717
rect 10048 18640 10100 18692
rect 14556 18708 14608 18760
rect 15660 18708 15712 18760
rect 16120 18751 16172 18760
rect 16120 18717 16129 18751
rect 16129 18717 16163 18751
rect 16163 18717 16172 18751
rect 16120 18708 16172 18717
rect 12808 18615 12860 18624
rect 12808 18581 12817 18615
rect 12817 18581 12851 18615
rect 12851 18581 12860 18615
rect 12808 18572 12860 18581
rect 22652 18572 22704 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 7748 18411 7800 18420
rect 7748 18377 7757 18411
rect 7757 18377 7791 18411
rect 7791 18377 7800 18411
rect 7748 18368 7800 18377
rect 8576 18411 8628 18420
rect 8576 18377 8585 18411
rect 8585 18377 8619 18411
rect 8619 18377 8628 18411
rect 8576 18368 8628 18377
rect 10232 18411 10284 18420
rect 10232 18377 10241 18411
rect 10241 18377 10275 18411
rect 10275 18377 10284 18411
rect 10232 18368 10284 18377
rect 12164 18411 12216 18420
rect 12164 18377 12173 18411
rect 12173 18377 12207 18411
rect 12207 18377 12216 18411
rect 12164 18368 12216 18377
rect 21548 18411 21600 18420
rect 21548 18377 21557 18411
rect 21557 18377 21591 18411
rect 21591 18377 21600 18411
rect 21548 18368 21600 18377
rect 22468 18411 22520 18420
rect 22468 18377 22477 18411
rect 22477 18377 22511 18411
rect 22511 18377 22520 18411
rect 22468 18368 22520 18377
rect 13728 18300 13780 18352
rect 15568 18300 15620 18352
rect 15660 18300 15712 18352
rect 21456 18300 21508 18352
rect 8024 18232 8076 18284
rect 9036 18232 9088 18284
rect 10876 18275 10928 18284
rect 10876 18241 10885 18275
rect 10885 18241 10919 18275
rect 10919 18241 10928 18275
rect 10876 18232 10928 18241
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 15936 18232 15988 18284
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 8760 18164 8812 18216
rect 12808 18207 12860 18216
rect 12808 18173 12817 18207
rect 12817 18173 12851 18207
rect 12851 18173 12860 18207
rect 12808 18164 12860 18173
rect 12900 18164 12952 18216
rect 19524 18207 19576 18216
rect 19524 18173 19542 18207
rect 19542 18173 19576 18207
rect 19524 18164 19576 18173
rect 22468 18164 22520 18216
rect 9588 18139 9640 18148
rect 8208 18071 8260 18080
rect 8208 18037 8217 18071
rect 8217 18037 8251 18071
rect 8251 18037 8260 18071
rect 8208 18028 8260 18037
rect 9588 18105 9597 18139
rect 9597 18105 9631 18139
rect 9631 18105 9640 18139
rect 9588 18096 9640 18105
rect 10968 18139 11020 18148
rect 10968 18105 10977 18139
rect 10977 18105 11011 18139
rect 11011 18105 11020 18139
rect 10968 18096 11020 18105
rect 11888 18096 11940 18148
rect 13360 18139 13412 18148
rect 13360 18105 13369 18139
rect 13369 18105 13403 18139
rect 13403 18105 13412 18139
rect 13360 18096 13412 18105
rect 14280 18139 14332 18148
rect 14280 18105 14289 18139
rect 14289 18105 14323 18139
rect 14323 18105 14332 18139
rect 14280 18096 14332 18105
rect 20536 18139 20588 18148
rect 9496 18028 9548 18080
rect 9864 18071 9916 18080
rect 9864 18037 9873 18071
rect 9873 18037 9907 18071
rect 9907 18037 9916 18071
rect 9864 18028 9916 18037
rect 13728 18071 13780 18080
rect 13728 18037 13737 18071
rect 13737 18037 13771 18071
rect 13771 18037 13780 18071
rect 13728 18028 13780 18037
rect 15384 18028 15436 18080
rect 20536 18105 20545 18139
rect 20545 18105 20579 18139
rect 20579 18105 20588 18139
rect 20536 18096 20588 18105
rect 19432 18028 19484 18080
rect 21456 18096 21508 18148
rect 21088 18028 21140 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 9036 17867 9088 17876
rect 9036 17833 9045 17867
rect 9045 17833 9079 17867
rect 9079 17833 9088 17867
rect 9036 17824 9088 17833
rect 11704 17824 11756 17876
rect 7472 17756 7524 17808
rect 8208 17799 8260 17808
rect 8208 17765 8217 17799
rect 8217 17765 8251 17799
rect 8251 17765 8260 17799
rect 8208 17756 8260 17765
rect 10692 17756 10744 17808
rect 11244 17756 11296 17808
rect 11796 17799 11848 17808
rect 11796 17765 11805 17799
rect 11805 17765 11839 17799
rect 11839 17765 11848 17799
rect 11796 17756 11848 17765
rect 13360 17824 13412 17876
rect 14096 17824 14148 17876
rect 20536 17867 20588 17876
rect 20536 17833 20545 17867
rect 20545 17833 20579 17867
rect 20579 17833 20588 17867
rect 20536 17824 20588 17833
rect 24768 17867 24820 17876
rect 24768 17833 24777 17867
rect 24777 17833 24811 17867
rect 24811 17833 24820 17867
rect 24768 17824 24820 17833
rect 15476 17799 15528 17808
rect 15476 17765 15485 17799
rect 15485 17765 15519 17799
rect 15519 17765 15528 17799
rect 15476 17756 15528 17765
rect 19432 17799 19484 17808
rect 19432 17765 19441 17799
rect 19441 17765 19475 17799
rect 19475 17765 19484 17799
rect 19432 17756 19484 17765
rect 21088 17799 21140 17808
rect 21088 17765 21097 17799
rect 21097 17765 21131 17799
rect 21131 17765 21140 17799
rect 21088 17756 21140 17765
rect 21548 17756 21600 17808
rect 22652 17799 22704 17808
rect 22652 17765 22661 17799
rect 22661 17765 22695 17799
rect 22695 17765 22704 17799
rect 22652 17756 22704 17765
rect 23112 17756 23164 17808
rect 17684 17731 17736 17740
rect 17684 17697 17693 17731
rect 17693 17697 17727 17731
rect 17727 17697 17736 17731
rect 17684 17688 17736 17697
rect 17960 17688 18012 17740
rect 24216 17688 24268 17740
rect 8116 17663 8168 17672
rect 8116 17629 8125 17663
rect 8125 17629 8159 17663
rect 8159 17629 8168 17663
rect 8116 17620 8168 17629
rect 10048 17663 10100 17672
rect 10048 17629 10057 17663
rect 10057 17629 10091 17663
rect 10091 17629 10100 17663
rect 10048 17620 10100 17629
rect 11888 17620 11940 17672
rect 12072 17663 12124 17672
rect 12072 17629 12081 17663
rect 12081 17629 12115 17663
rect 12115 17629 12124 17663
rect 12072 17620 12124 17629
rect 13360 17663 13412 17672
rect 13360 17629 13369 17663
rect 13369 17629 13403 17663
rect 13403 17629 13412 17663
rect 13360 17620 13412 17629
rect 8760 17552 8812 17604
rect 10784 17595 10836 17604
rect 10784 17561 10793 17595
rect 10793 17561 10827 17595
rect 10827 17561 10836 17595
rect 10784 17552 10836 17561
rect 14556 17620 14608 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 18420 17663 18472 17672
rect 18420 17629 18429 17663
rect 18429 17629 18463 17663
rect 18463 17629 18472 17663
rect 18420 17620 18472 17629
rect 19340 17663 19392 17672
rect 19340 17629 19349 17663
rect 19349 17629 19383 17663
rect 19383 17629 19392 17663
rect 19340 17620 19392 17629
rect 21180 17620 21232 17672
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 22376 17620 22428 17672
rect 9864 17484 9916 17536
rect 15936 17552 15988 17604
rect 22744 17552 22796 17604
rect 12900 17484 12952 17536
rect 14280 17484 14332 17536
rect 15568 17484 15620 17536
rect 17592 17484 17644 17536
rect 22468 17484 22520 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 7472 17323 7524 17332
rect 7472 17289 7481 17323
rect 7481 17289 7515 17323
rect 7515 17289 7524 17323
rect 7472 17280 7524 17289
rect 8116 17280 8168 17332
rect 9496 17280 9548 17332
rect 11796 17323 11848 17332
rect 11796 17289 11805 17323
rect 11805 17289 11839 17323
rect 11839 17289 11848 17323
rect 11796 17280 11848 17289
rect 15384 17323 15436 17332
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 15568 17280 15620 17332
rect 22652 17280 22704 17332
rect 15476 17212 15528 17264
rect 20904 17212 20956 17264
rect 23112 17255 23164 17264
rect 23112 17221 23121 17255
rect 23121 17221 23155 17255
rect 23155 17221 23164 17255
rect 23112 17212 23164 17221
rect 7196 17144 7248 17196
rect 14096 17187 14148 17196
rect 14096 17153 14105 17187
rect 14105 17153 14139 17187
rect 14139 17153 14148 17187
rect 14096 17144 14148 17153
rect 15568 17144 15620 17196
rect 17408 17144 17460 17196
rect 17960 17144 18012 17196
rect 6092 17076 6144 17128
rect 7656 17119 7708 17128
rect 7656 17085 7674 17119
rect 7674 17085 7708 17119
rect 7656 17076 7708 17085
rect 8668 17119 8720 17128
rect 8668 17085 8677 17119
rect 8677 17085 8711 17119
rect 8711 17085 8720 17119
rect 8668 17076 8720 17085
rect 12624 17119 12676 17128
rect 12624 17085 12633 17119
rect 12633 17085 12667 17119
rect 12667 17085 12676 17119
rect 12624 17076 12676 17085
rect 12900 17119 12952 17128
rect 12900 17085 12909 17119
rect 12909 17085 12943 17119
rect 12943 17085 12952 17119
rect 12900 17076 12952 17085
rect 16764 17076 16816 17128
rect 10048 17008 10100 17060
rect 13176 17051 13228 17060
rect 13176 17017 13185 17051
rect 13185 17017 13219 17051
rect 13219 17017 13228 17051
rect 13176 17008 13228 17017
rect 15936 17051 15988 17060
rect 11704 16940 11756 16992
rect 13452 16983 13504 16992
rect 13452 16949 13461 16983
rect 13461 16949 13495 16983
rect 13495 16949 13504 16983
rect 13452 16940 13504 16949
rect 13912 16983 13964 16992
rect 13912 16949 13921 16983
rect 13921 16949 13955 16983
rect 13955 16949 13964 16983
rect 15936 17017 15945 17051
rect 15945 17017 15979 17051
rect 15979 17017 15988 17051
rect 15936 17008 15988 17017
rect 13912 16940 13964 16949
rect 15384 16940 15436 16992
rect 16212 16940 16264 16992
rect 17592 16940 17644 16992
rect 22468 17076 22520 17128
rect 23848 17076 23900 17128
rect 18788 17008 18840 17060
rect 18696 16940 18748 16992
rect 18972 16983 19024 16992
rect 18972 16949 18981 16983
rect 18981 16949 19015 16983
rect 19015 16949 19024 16983
rect 19432 17008 19484 17060
rect 20628 17008 20680 17060
rect 20904 17051 20956 17060
rect 20904 17017 20913 17051
rect 20913 17017 20947 17051
rect 20947 17017 20956 17051
rect 20904 17008 20956 17017
rect 21456 17051 21508 17060
rect 21456 17017 21465 17051
rect 21465 17017 21499 17051
rect 21499 17017 21508 17051
rect 21456 17008 21508 17017
rect 18972 16940 19024 16949
rect 21548 16940 21600 16992
rect 22560 16940 22612 16992
rect 24216 16940 24268 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 8116 16736 8168 16788
rect 10048 16779 10100 16788
rect 10048 16745 10057 16779
rect 10057 16745 10091 16779
rect 10091 16745 10100 16779
rect 10048 16736 10100 16745
rect 10692 16736 10744 16788
rect 14556 16736 14608 16788
rect 16212 16779 16264 16788
rect 16212 16745 16221 16779
rect 16221 16745 16255 16779
rect 16255 16745 16264 16779
rect 16212 16736 16264 16745
rect 19248 16736 19300 16788
rect 7196 16711 7248 16720
rect 7196 16677 7205 16711
rect 7205 16677 7239 16711
rect 7239 16677 7248 16711
rect 7196 16668 7248 16677
rect 8668 16668 8720 16720
rect 11612 16711 11664 16720
rect 11612 16677 11621 16711
rect 11621 16677 11655 16711
rect 11655 16677 11664 16711
rect 11612 16668 11664 16677
rect 11704 16711 11756 16720
rect 11704 16677 11713 16711
rect 11713 16677 11747 16711
rect 11747 16677 11756 16711
rect 11704 16668 11756 16677
rect 13452 16668 13504 16720
rect 13544 16668 13596 16720
rect 13820 16711 13872 16720
rect 13820 16677 13829 16711
rect 13829 16677 13863 16711
rect 13863 16677 13872 16711
rect 13820 16668 13872 16677
rect 15292 16668 15344 16720
rect 20996 16736 21048 16788
rect 21548 16736 21600 16788
rect 20812 16668 20864 16720
rect 21180 16668 21232 16720
rect 22560 16711 22612 16720
rect 22560 16677 22569 16711
rect 22569 16677 22603 16711
rect 22603 16677 22612 16711
rect 22560 16668 22612 16677
rect 23204 16668 23256 16720
rect 6736 16643 6788 16652
rect 6736 16609 6745 16643
rect 6745 16609 6779 16643
rect 6779 16609 6788 16643
rect 6736 16600 6788 16609
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 8392 16600 8444 16652
rect 17040 16643 17092 16652
rect 17040 16609 17049 16643
rect 17049 16609 17083 16643
rect 17083 16609 17092 16643
rect 17040 16600 17092 16609
rect 17408 16600 17460 16652
rect 18420 16600 18472 16652
rect 19616 16600 19668 16652
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 11888 16575 11940 16584
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 11888 16532 11940 16541
rect 14832 16532 14884 16584
rect 18052 16575 18104 16584
rect 18052 16541 18061 16575
rect 18061 16541 18095 16575
rect 18095 16541 18104 16575
rect 18052 16532 18104 16541
rect 22192 16532 22244 16584
rect 22376 16532 22428 16584
rect 12624 16439 12676 16448
rect 12624 16405 12633 16439
rect 12633 16405 12667 16439
rect 12667 16405 12676 16439
rect 12624 16396 12676 16405
rect 18788 16439 18840 16448
rect 18788 16405 18797 16439
rect 18797 16405 18831 16439
rect 18831 16405 18840 16439
rect 18788 16396 18840 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 8116 16235 8168 16244
rect 8116 16201 8125 16235
rect 8125 16201 8159 16235
rect 8159 16201 8168 16235
rect 8116 16192 8168 16201
rect 9680 16192 9732 16244
rect 9772 16235 9824 16244
rect 9772 16201 9781 16235
rect 9781 16201 9815 16235
rect 9815 16201 9824 16235
rect 9772 16192 9824 16201
rect 10048 16192 10100 16244
rect 10784 16124 10836 16176
rect 11612 16192 11664 16244
rect 13820 16192 13872 16244
rect 14832 16192 14884 16244
rect 16028 16192 16080 16244
rect 18972 16235 19024 16244
rect 9588 16056 9640 16108
rect 11704 16056 11756 16108
rect 8300 16031 8352 16040
rect 8300 15997 8309 16031
rect 8309 15997 8343 16031
rect 8343 15997 8352 16031
rect 8300 15988 8352 15997
rect 8392 15988 8444 16040
rect 6736 15920 6788 15972
rect 8944 15920 8996 15972
rect 9956 15963 10008 15972
rect 9956 15929 9965 15963
rect 9965 15929 9999 15963
rect 9999 15929 10008 15963
rect 9956 15920 10008 15929
rect 13176 16056 13228 16108
rect 16120 16124 16172 16176
rect 15844 16099 15896 16108
rect 15844 16065 15853 16099
rect 15853 16065 15887 16099
rect 15887 16065 15896 16099
rect 15844 16056 15896 16065
rect 18052 16099 18104 16108
rect 18052 16065 18061 16099
rect 18061 16065 18095 16099
rect 18095 16065 18104 16099
rect 18052 16056 18104 16065
rect 18972 16201 18981 16235
rect 18981 16201 19015 16235
rect 19015 16201 19024 16235
rect 18972 16192 19024 16201
rect 19340 16192 19392 16244
rect 20812 16192 20864 16244
rect 22192 16235 22244 16244
rect 22192 16201 22201 16235
rect 22201 16201 22235 16235
rect 22235 16201 22244 16235
rect 22192 16192 22244 16201
rect 22928 16235 22980 16244
rect 22928 16201 22937 16235
rect 22937 16201 22971 16235
rect 22971 16201 22980 16235
rect 22928 16192 22980 16201
rect 23204 16235 23256 16244
rect 23204 16201 23213 16235
rect 23213 16201 23247 16235
rect 23247 16201 23256 16235
rect 23204 16192 23256 16201
rect 19616 16167 19668 16176
rect 19616 16133 19625 16167
rect 19625 16133 19659 16167
rect 19659 16133 19668 16167
rect 19616 16124 19668 16133
rect 18604 16056 18656 16108
rect 17224 15988 17276 16040
rect 18972 15988 19024 16040
rect 21180 16056 21232 16108
rect 22928 15988 22980 16040
rect 13452 15920 13504 15972
rect 13912 15920 13964 15972
rect 15292 15963 15344 15972
rect 15292 15929 15301 15963
rect 15301 15929 15335 15963
rect 15335 15929 15344 15963
rect 15292 15920 15344 15929
rect 10140 15852 10192 15904
rect 13728 15852 13780 15904
rect 16028 15920 16080 15972
rect 17040 15963 17092 15972
rect 17040 15929 17049 15963
rect 17049 15929 17083 15963
rect 17083 15929 17092 15963
rect 17040 15920 17092 15929
rect 20996 15963 21048 15972
rect 20996 15929 21005 15963
rect 21005 15929 21039 15963
rect 21039 15929 21048 15963
rect 20996 15920 21048 15929
rect 21732 15920 21784 15972
rect 16120 15852 16172 15904
rect 17408 15895 17460 15904
rect 17408 15861 17417 15895
rect 17417 15861 17451 15895
rect 17451 15861 17460 15895
rect 17408 15852 17460 15861
rect 17776 15895 17828 15904
rect 17776 15861 17785 15895
rect 17785 15861 17819 15895
rect 17819 15861 17828 15895
rect 17776 15852 17828 15861
rect 19340 15895 19392 15904
rect 19340 15861 19349 15895
rect 19349 15861 19383 15895
rect 19383 15861 19392 15895
rect 19340 15852 19392 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 13176 15691 13228 15700
rect 13176 15657 13185 15691
rect 13185 15657 13219 15691
rect 13219 15657 13228 15691
rect 13176 15648 13228 15657
rect 13544 15691 13596 15700
rect 13544 15657 13553 15691
rect 13553 15657 13587 15691
rect 13587 15657 13596 15691
rect 13544 15648 13596 15657
rect 15936 15648 15988 15700
rect 21180 15648 21232 15700
rect 22560 15691 22612 15700
rect 22560 15657 22569 15691
rect 22569 15657 22603 15691
rect 22603 15657 22612 15691
rect 22560 15648 22612 15657
rect 10048 15580 10100 15632
rect 10508 15580 10560 15632
rect 10968 15580 11020 15632
rect 13728 15580 13780 15632
rect 15476 15623 15528 15632
rect 15476 15589 15485 15623
rect 15485 15589 15519 15623
rect 15519 15589 15528 15623
rect 15476 15580 15528 15589
rect 16212 15580 16264 15632
rect 17776 15580 17828 15632
rect 20812 15580 20864 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 10784 15512 10836 15564
rect 12072 15555 12124 15564
rect 12072 15521 12081 15555
rect 12081 15521 12115 15555
rect 12115 15521 12124 15555
rect 12072 15512 12124 15521
rect 20260 15512 20312 15564
rect 9864 15444 9916 15496
rect 11704 15444 11756 15496
rect 12992 15444 13044 15496
rect 15568 15444 15620 15496
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 17960 15487 18012 15496
rect 17960 15453 17969 15487
rect 17969 15453 18003 15487
rect 18003 15453 18012 15487
rect 17960 15444 18012 15453
rect 20628 15444 20680 15496
rect 21364 15444 21416 15496
rect 21732 15444 21784 15496
rect 1492 15376 1544 15428
rect 2044 15376 2096 15428
rect 8300 15376 8352 15428
rect 12808 15376 12860 15428
rect 21088 15376 21140 15428
rect 21548 15376 21600 15428
rect 8392 15351 8444 15360
rect 8392 15317 8401 15351
rect 8401 15317 8435 15351
rect 8435 15317 8444 15351
rect 8392 15308 8444 15317
rect 9312 15351 9364 15360
rect 9312 15317 9321 15351
rect 9321 15317 9355 15351
rect 9355 15317 9364 15351
rect 9312 15308 9364 15317
rect 9956 15308 10008 15360
rect 12072 15308 12124 15360
rect 19156 15351 19208 15360
rect 19156 15317 19165 15351
rect 19165 15317 19199 15351
rect 19199 15317 19208 15351
rect 19156 15308 19208 15317
rect 20444 15308 20496 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 9772 15104 9824 15156
rect 10140 15104 10192 15156
rect 10508 15147 10560 15156
rect 10508 15113 10517 15147
rect 10517 15113 10551 15147
rect 10551 15113 10560 15147
rect 10508 15104 10560 15113
rect 10968 15104 11020 15156
rect 13728 15104 13780 15156
rect 13820 15104 13872 15156
rect 15476 15104 15528 15156
rect 15568 15104 15620 15156
rect 17960 15104 18012 15156
rect 18788 15104 18840 15156
rect 20996 15104 21048 15156
rect 21364 15104 21416 15156
rect 22376 15147 22428 15156
rect 22376 15113 22385 15147
rect 22385 15113 22419 15147
rect 22419 15113 22428 15147
rect 22376 15104 22428 15113
rect 9128 15036 9180 15088
rect 22284 15036 22336 15088
rect 8116 14968 8168 15020
rect 12164 15011 12216 15020
rect 12164 14977 12173 15011
rect 12173 14977 12207 15011
rect 12207 14977 12216 15011
rect 12164 14968 12216 14977
rect 9312 14943 9364 14952
rect 9312 14909 9321 14943
rect 9321 14909 9355 14943
rect 9355 14909 9364 14943
rect 9312 14900 9364 14909
rect 9772 14900 9824 14952
rect 16028 14968 16080 15020
rect 16212 15011 16264 15020
rect 16212 14977 16221 15011
rect 16221 14977 16255 15011
rect 16255 14977 16264 15011
rect 16212 14968 16264 14977
rect 19156 14968 19208 15020
rect 21456 14968 21508 15020
rect 12532 14900 12584 14952
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 12900 14900 12952 14909
rect 17684 14900 17736 14952
rect 19340 14900 19392 14952
rect 12992 14832 13044 14884
rect 13176 14875 13228 14884
rect 13176 14841 13185 14875
rect 13185 14841 13219 14875
rect 13219 14841 13228 14875
rect 13176 14832 13228 14841
rect 14188 14875 14240 14884
rect 14188 14841 14197 14875
rect 14197 14841 14231 14875
rect 14231 14841 14240 14875
rect 14188 14832 14240 14841
rect 15752 14875 15804 14884
rect 1400 14764 1452 14816
rect 5264 14764 5316 14816
rect 8576 14764 8628 14816
rect 9680 14807 9732 14816
rect 9680 14773 9689 14807
rect 9689 14773 9723 14807
rect 9723 14773 9732 14807
rect 9680 14764 9732 14773
rect 13820 14764 13872 14816
rect 15752 14841 15761 14875
rect 15761 14841 15795 14875
rect 15795 14841 15804 14875
rect 15752 14832 15804 14841
rect 15936 14764 15988 14816
rect 16856 14764 16908 14816
rect 17776 14807 17828 14816
rect 17776 14773 17785 14807
rect 17785 14773 17819 14807
rect 17819 14773 17828 14807
rect 17776 14764 17828 14773
rect 20168 14832 20220 14884
rect 21732 14875 21784 14884
rect 20260 14807 20312 14816
rect 20260 14773 20269 14807
rect 20269 14773 20303 14807
rect 20303 14773 20312 14807
rect 20260 14764 20312 14773
rect 20352 14764 20404 14816
rect 20812 14807 20864 14816
rect 20812 14773 20821 14807
rect 20821 14773 20855 14807
rect 20855 14773 20864 14807
rect 20812 14764 20864 14773
rect 21732 14841 21741 14875
rect 21741 14841 21775 14875
rect 21775 14841 21784 14875
rect 21732 14832 21784 14841
rect 24032 14832 24084 14884
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 9864 14603 9916 14612
rect 9864 14569 9873 14603
rect 9873 14569 9907 14603
rect 9907 14569 9916 14603
rect 9864 14560 9916 14569
rect 10968 14560 11020 14612
rect 11520 14560 11572 14612
rect 11704 14603 11756 14612
rect 11704 14569 11713 14603
rect 11713 14569 11747 14603
rect 11747 14569 11756 14603
rect 11704 14560 11756 14569
rect 12256 14560 12308 14612
rect 12992 14603 13044 14612
rect 12992 14569 13001 14603
rect 13001 14569 13035 14603
rect 13035 14569 13044 14603
rect 12992 14560 13044 14569
rect 13452 14603 13504 14612
rect 13452 14569 13461 14603
rect 13461 14569 13495 14603
rect 13495 14569 13504 14603
rect 13452 14560 13504 14569
rect 13820 14560 13872 14612
rect 15660 14603 15712 14612
rect 15660 14569 15669 14603
rect 15669 14569 15703 14603
rect 15703 14569 15712 14603
rect 15660 14560 15712 14569
rect 16120 14560 16172 14612
rect 19340 14560 19392 14612
rect 20352 14560 20404 14612
rect 20444 14560 20496 14612
rect 9680 14492 9732 14544
rect 17960 14492 18012 14544
rect 21364 14560 21416 14612
rect 21088 14535 21140 14544
rect 21088 14501 21097 14535
rect 21097 14501 21131 14535
rect 21131 14501 21140 14535
rect 21088 14492 21140 14501
rect 22284 14492 22336 14544
rect 8208 14467 8260 14476
rect 8208 14433 8217 14467
rect 8217 14433 8251 14467
rect 8251 14433 8260 14467
rect 8208 14424 8260 14433
rect 8392 14424 8444 14476
rect 9036 14424 9088 14476
rect 17316 14467 17368 14476
rect 17316 14433 17325 14467
rect 17325 14433 17359 14467
rect 17359 14433 17368 14467
rect 17316 14424 17368 14433
rect 17408 14424 17460 14476
rect 20812 14424 20864 14476
rect 21916 14424 21968 14476
rect 24032 14467 24084 14476
rect 24032 14433 24041 14467
rect 24041 14433 24075 14467
rect 24075 14433 24084 14467
rect 24032 14424 24084 14433
rect 10692 14356 10744 14408
rect 13176 14356 13228 14408
rect 15384 14356 15436 14408
rect 21272 14399 21324 14408
rect 9220 14263 9272 14272
rect 9220 14229 9229 14263
rect 9229 14229 9263 14263
rect 9263 14229 9272 14263
rect 9220 14220 9272 14229
rect 12440 14263 12492 14272
rect 12440 14229 12449 14263
rect 12449 14229 12483 14263
rect 12483 14229 12492 14263
rect 12440 14220 12492 14229
rect 14188 14220 14240 14272
rect 18052 14263 18104 14272
rect 18052 14229 18061 14263
rect 18061 14229 18095 14263
rect 18095 14229 18104 14263
rect 18052 14220 18104 14229
rect 18880 14263 18932 14272
rect 18880 14229 18889 14263
rect 18889 14229 18923 14263
rect 18923 14229 18932 14263
rect 21272 14365 21281 14399
rect 21281 14365 21315 14399
rect 21315 14365 21324 14399
rect 21272 14356 21324 14365
rect 18880 14220 18932 14229
rect 23756 14220 23808 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 9680 14016 9732 14068
rect 10048 14016 10100 14068
rect 11428 14059 11480 14068
rect 11428 14025 11437 14059
rect 11437 14025 11471 14059
rect 11471 14025 11480 14059
rect 11428 14016 11480 14025
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 13452 14059 13504 14068
rect 13452 14025 13461 14059
rect 13461 14025 13495 14059
rect 13495 14025 13504 14059
rect 13452 14016 13504 14025
rect 15476 14016 15528 14068
rect 16028 14016 16080 14068
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 7932 13855 7984 13864
rect 7932 13821 7941 13855
rect 7941 13821 7975 13855
rect 7975 13821 7984 13855
rect 7932 13812 7984 13821
rect 8116 13855 8168 13864
rect 8116 13821 8125 13855
rect 8125 13821 8159 13855
rect 8159 13821 8168 13855
rect 10876 13948 10928 14000
rect 8116 13812 8168 13821
rect 8392 13787 8444 13796
rect 8392 13753 8401 13787
rect 8401 13753 8435 13787
rect 8435 13753 8444 13787
rect 8392 13744 8444 13753
rect 11428 13812 11480 13864
rect 12164 13812 12216 13864
rect 13636 13948 13688 14000
rect 13084 13880 13136 13932
rect 17316 14016 17368 14068
rect 18236 14059 18288 14068
rect 18236 14025 18245 14059
rect 18245 14025 18279 14059
rect 18279 14025 18288 14059
rect 18236 14016 18288 14025
rect 20168 14059 20220 14068
rect 14280 13855 14332 13864
rect 14280 13821 14289 13855
rect 14289 13821 14323 13855
rect 14323 13821 14332 13855
rect 14280 13812 14332 13821
rect 16672 13812 16724 13864
rect 17500 13948 17552 14000
rect 20168 14025 20177 14059
rect 20177 14025 20211 14059
rect 20211 14025 20220 14059
rect 20168 14016 20220 14025
rect 22284 14016 22336 14068
rect 22928 14016 22980 14068
rect 18880 13880 18932 13932
rect 17408 13855 17460 13864
rect 17408 13821 17417 13855
rect 17417 13821 17451 13855
rect 17451 13821 17460 13855
rect 17408 13812 17460 13821
rect 18052 13812 18104 13864
rect 11336 13744 11388 13796
rect 13084 13744 13136 13796
rect 15660 13744 15712 13796
rect 8208 13676 8260 13728
rect 9036 13676 9088 13728
rect 9634 13676 9686 13728
rect 10968 13676 11020 13728
rect 19340 13676 19392 13728
rect 20168 13676 20220 13728
rect 20812 13855 20864 13864
rect 20812 13821 20821 13855
rect 20821 13821 20855 13855
rect 20855 13821 20864 13855
rect 20812 13812 20864 13821
rect 21272 13812 21324 13864
rect 22928 13812 22980 13864
rect 24860 14016 24912 14068
rect 21916 13744 21968 13796
rect 23296 13744 23348 13796
rect 24032 13744 24084 13796
rect 22100 13676 22152 13728
rect 23664 13676 23716 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 9128 13472 9180 13524
rect 9588 13472 9640 13524
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 10968 13472 11020 13524
rect 13176 13472 13228 13524
rect 20168 13515 20220 13524
rect 20168 13481 20177 13515
rect 20177 13481 20211 13515
rect 20211 13481 20220 13515
rect 20168 13472 20220 13481
rect 20996 13472 21048 13524
rect 23664 13472 23716 13524
rect 7932 13404 7984 13456
rect 11336 13447 11388 13456
rect 8024 13379 8076 13388
rect 8024 13345 8033 13379
rect 8033 13345 8067 13379
rect 8067 13345 8076 13379
rect 8024 13336 8076 13345
rect 8116 13336 8168 13388
rect 11336 13413 11345 13447
rect 11345 13413 11379 13447
rect 11379 13413 11388 13447
rect 11336 13404 11388 13413
rect 11520 13404 11572 13456
rect 11796 13404 11848 13456
rect 9956 13379 10008 13388
rect 9956 13345 9965 13379
rect 9965 13345 9999 13379
rect 9999 13345 10008 13379
rect 9956 13336 10008 13345
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 12808 13336 12860 13388
rect 13636 13379 13688 13388
rect 8760 13311 8812 13320
rect 8760 13277 8769 13311
rect 8769 13277 8803 13311
rect 8803 13277 8812 13311
rect 8760 13268 8812 13277
rect 9220 13268 9272 13320
rect 9864 13200 9916 13252
rect 13636 13345 13645 13379
rect 13645 13345 13679 13379
rect 13679 13345 13688 13379
rect 13636 13336 13688 13345
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 19064 13404 19116 13456
rect 19340 13404 19392 13456
rect 20812 13404 20864 13456
rect 22836 13447 22888 13456
rect 22836 13413 22845 13447
rect 22845 13413 22879 13447
rect 22879 13413 22888 13447
rect 22836 13404 22888 13413
rect 22928 13447 22980 13456
rect 22928 13413 22937 13447
rect 22937 13413 22971 13447
rect 22971 13413 22980 13447
rect 22928 13404 22980 13413
rect 16028 13379 16080 13388
rect 16028 13345 16037 13379
rect 16037 13345 16071 13379
rect 16071 13345 16080 13379
rect 16028 13336 16080 13345
rect 16580 13336 16632 13388
rect 17316 13379 17368 13388
rect 17316 13345 17325 13379
rect 17325 13345 17359 13379
rect 17359 13345 17368 13379
rect 17316 13336 17368 13345
rect 17408 13336 17460 13388
rect 24768 13336 24820 13388
rect 26240 13336 26292 13388
rect 15384 13268 15436 13320
rect 18512 13268 18564 13320
rect 18880 13311 18932 13320
rect 18880 13277 18889 13311
rect 18889 13277 18923 13311
rect 18923 13277 18932 13311
rect 18880 13268 18932 13277
rect 20628 13268 20680 13320
rect 21732 13268 21784 13320
rect 24032 13268 24084 13320
rect 14280 13243 14332 13252
rect 14280 13209 14289 13243
rect 14289 13209 14323 13243
rect 14323 13209 14332 13243
rect 14280 13200 14332 13209
rect 14648 13200 14700 13252
rect 9220 13175 9272 13184
rect 9220 13141 9229 13175
rect 9229 13141 9263 13175
rect 9263 13141 9272 13175
rect 9220 13132 9272 13141
rect 18696 13132 18748 13184
rect 22652 13132 22704 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 112 12928 164 12980
rect 8116 12971 8168 12980
rect 8116 12937 8125 12971
rect 8125 12937 8159 12971
rect 8159 12937 8168 12971
rect 8116 12928 8168 12937
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 12808 12971 12860 12980
rect 12808 12937 12817 12971
rect 12817 12937 12851 12971
rect 12851 12937 12860 12971
rect 12808 12928 12860 12937
rect 12992 12928 13044 12980
rect 13636 12928 13688 12980
rect 15936 12971 15988 12980
rect 8024 12860 8076 12912
rect 9220 12860 9272 12912
rect 10968 12792 11020 12844
rect 11336 12860 11388 12912
rect 12716 12860 12768 12912
rect 15936 12937 15945 12971
rect 15945 12937 15979 12971
rect 15979 12937 15988 12971
rect 15936 12928 15988 12937
rect 17408 12971 17460 12980
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 21088 12928 21140 12980
rect 22928 12928 22980 12980
rect 24768 12971 24820 12980
rect 24768 12937 24777 12971
rect 24777 12937 24811 12971
rect 24811 12937 24820 12971
rect 24768 12928 24820 12937
rect 27620 12928 27672 12980
rect 16028 12860 16080 12912
rect 18052 12860 18104 12912
rect 19340 12903 19392 12912
rect 19340 12869 19349 12903
rect 19349 12869 19383 12903
rect 19383 12869 19392 12903
rect 20168 12903 20220 12912
rect 19340 12860 19392 12869
rect 20168 12869 20177 12903
rect 20177 12869 20211 12903
rect 20211 12869 20220 12903
rect 20168 12860 20220 12869
rect 23664 12860 23716 12912
rect 9680 12767 9732 12776
rect 9680 12733 9689 12767
rect 9689 12733 9723 12767
rect 9723 12733 9732 12767
rect 9680 12724 9732 12733
rect 9036 12656 9088 12708
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 14924 12792 14976 12801
rect 16672 12792 16724 12844
rect 16580 12767 16632 12776
rect 16580 12733 16589 12767
rect 16589 12733 16623 12767
rect 16623 12733 16632 12767
rect 16580 12724 16632 12733
rect 16764 12724 16816 12776
rect 18696 12724 18748 12776
rect 18880 12792 18932 12844
rect 20260 12792 20312 12844
rect 20352 12792 20404 12844
rect 22100 12792 22152 12844
rect 22376 12792 22428 12844
rect 10140 12656 10192 12708
rect 10968 12699 11020 12708
rect 10968 12665 10977 12699
rect 10977 12665 11011 12699
rect 11011 12665 11020 12699
rect 10968 12656 11020 12665
rect 12624 12656 12676 12708
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 9312 12631 9364 12640
rect 9312 12597 9321 12631
rect 9321 12597 9355 12631
rect 9355 12597 9364 12631
rect 9312 12588 9364 12597
rect 13452 12699 13504 12708
rect 13452 12665 13461 12699
rect 13461 12665 13495 12699
rect 13495 12665 13504 12699
rect 13452 12656 13504 12665
rect 13912 12588 13964 12640
rect 14648 12588 14700 12640
rect 14832 12588 14884 12640
rect 18144 12656 18196 12708
rect 20076 12724 20128 12776
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 24032 12835 24084 12844
rect 24032 12801 24041 12835
rect 24041 12801 24075 12835
rect 24075 12801 24084 12835
rect 24032 12792 24084 12801
rect 24860 12724 24912 12776
rect 17868 12631 17920 12640
rect 17868 12597 17877 12631
rect 17877 12597 17911 12631
rect 17911 12597 17920 12631
rect 20444 12656 20496 12708
rect 21732 12699 21784 12708
rect 17868 12588 17920 12597
rect 20168 12588 20220 12640
rect 21732 12665 21741 12699
rect 21741 12665 21775 12699
rect 21775 12665 21784 12699
rect 21732 12656 21784 12665
rect 22284 12656 22336 12708
rect 22192 12588 22244 12640
rect 22928 12588 22980 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 10876 12427 10928 12436
rect 10876 12393 10885 12427
rect 10885 12393 10919 12427
rect 10919 12393 10928 12427
rect 10876 12384 10928 12393
rect 10968 12384 11020 12436
rect 9956 12359 10008 12368
rect 9956 12325 9965 12359
rect 9965 12325 9999 12359
rect 9999 12325 10008 12359
rect 9956 12316 10008 12325
rect 11888 12316 11940 12368
rect 13544 12384 13596 12436
rect 14188 12384 14240 12436
rect 14924 12427 14976 12436
rect 14924 12393 14933 12427
rect 14933 12393 14967 12427
rect 14967 12393 14976 12427
rect 14924 12384 14976 12393
rect 16764 12427 16816 12436
rect 13636 12316 13688 12368
rect 16764 12393 16773 12427
rect 16773 12393 16807 12427
rect 16807 12393 16816 12427
rect 16764 12384 16816 12393
rect 17316 12427 17368 12436
rect 17316 12393 17325 12427
rect 17325 12393 17359 12427
rect 17359 12393 17368 12427
rect 17316 12384 17368 12393
rect 20076 12384 20128 12436
rect 20352 12427 20404 12436
rect 20352 12393 20361 12427
rect 20361 12393 20395 12427
rect 20395 12393 20404 12427
rect 20352 12384 20404 12393
rect 23020 12384 23072 12436
rect 15476 12359 15528 12368
rect 15476 12325 15485 12359
rect 15485 12325 15519 12359
rect 15519 12325 15528 12359
rect 15476 12316 15528 12325
rect 16028 12359 16080 12368
rect 16028 12325 16037 12359
rect 16037 12325 16071 12359
rect 16071 12325 16080 12359
rect 16028 12316 16080 12325
rect 8760 12112 8812 12164
rect 8852 12112 8904 12164
rect 9312 12044 9364 12096
rect 10048 12044 10100 12096
rect 13912 12248 13964 12300
rect 12348 12223 12400 12232
rect 12348 12189 12357 12223
rect 12357 12189 12391 12223
rect 12391 12189 12400 12223
rect 12348 12180 12400 12189
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 13820 12180 13872 12232
rect 15384 12223 15436 12232
rect 15384 12189 15393 12223
rect 15393 12189 15427 12223
rect 15427 12189 15436 12223
rect 15384 12180 15436 12189
rect 11428 12112 11480 12164
rect 16580 12316 16632 12368
rect 17868 12316 17920 12368
rect 20168 12316 20220 12368
rect 20996 12359 21048 12368
rect 20996 12325 21005 12359
rect 21005 12325 21039 12359
rect 21039 12325 21048 12359
rect 20996 12316 21048 12325
rect 21088 12359 21140 12368
rect 21088 12325 21097 12359
rect 21097 12325 21131 12359
rect 21131 12325 21140 12359
rect 22652 12359 22704 12368
rect 21088 12316 21140 12325
rect 22652 12325 22661 12359
rect 22661 12325 22695 12359
rect 22695 12325 22704 12359
rect 22652 12316 22704 12325
rect 22928 12316 22980 12368
rect 19984 12248 20036 12300
rect 18328 12180 18380 12232
rect 21732 12180 21784 12232
rect 22560 12223 22612 12232
rect 22560 12189 22569 12223
rect 22569 12189 22603 12223
rect 22603 12189 22612 12223
rect 22560 12180 22612 12189
rect 22836 12223 22888 12232
rect 22836 12189 22845 12223
rect 22845 12189 22879 12223
rect 22879 12189 22888 12223
rect 22836 12180 22888 12189
rect 24768 12316 24820 12368
rect 24124 12223 24176 12232
rect 24124 12189 24133 12223
rect 24133 12189 24167 12223
rect 24167 12189 24176 12223
rect 24124 12180 24176 12189
rect 24216 12180 24268 12232
rect 16764 12112 16816 12164
rect 13360 12087 13412 12096
rect 13360 12053 13369 12087
rect 13369 12053 13403 12087
rect 13403 12053 13412 12087
rect 13360 12044 13412 12053
rect 19616 12087 19668 12096
rect 19616 12053 19625 12087
rect 19625 12053 19659 12087
rect 19659 12053 19668 12087
rect 19616 12044 19668 12053
rect 20628 12087 20680 12096
rect 20628 12053 20637 12087
rect 20637 12053 20671 12087
rect 20671 12053 20680 12087
rect 20628 12044 20680 12053
rect 23112 12044 23164 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 10876 11840 10928 11892
rect 11520 11883 11572 11892
rect 11520 11849 11529 11883
rect 11529 11849 11563 11883
rect 11563 11849 11572 11883
rect 11888 11883 11940 11892
rect 11520 11840 11572 11849
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 13728 11840 13780 11892
rect 14832 11840 14884 11892
rect 20628 11840 20680 11892
rect 20904 11883 20956 11892
rect 20904 11849 20913 11883
rect 20913 11849 20947 11883
rect 20947 11849 20956 11883
rect 20904 11840 20956 11849
rect 20996 11840 21048 11892
rect 22652 11840 22704 11892
rect 24768 11883 24820 11892
rect 1492 11636 1544 11688
rect 7932 11704 7984 11756
rect 9496 11747 9548 11756
rect 9496 11713 9505 11747
rect 9505 11713 9539 11747
rect 9539 11713 9548 11747
rect 9496 11704 9548 11713
rect 10876 11704 10928 11756
rect 7564 11543 7616 11552
rect 7564 11509 7573 11543
rect 7573 11509 7607 11543
rect 7607 11509 7616 11543
rect 8852 11636 8904 11688
rect 9128 11679 9180 11688
rect 9128 11645 9137 11679
rect 9137 11645 9171 11679
rect 9171 11645 9180 11679
rect 9128 11636 9180 11645
rect 9404 11636 9456 11688
rect 8208 11611 8260 11620
rect 8208 11577 8217 11611
rect 8217 11577 8251 11611
rect 8251 11577 8260 11611
rect 8208 11568 8260 11577
rect 16028 11772 16080 11824
rect 19340 11815 19392 11824
rect 19340 11781 19349 11815
rect 19349 11781 19383 11815
rect 19383 11781 19392 11815
rect 19340 11772 19392 11781
rect 18052 11704 18104 11756
rect 19616 11772 19668 11824
rect 24768 11849 24777 11883
rect 24777 11849 24811 11883
rect 24811 11849 24820 11883
rect 24768 11840 24820 11849
rect 23572 11772 23624 11824
rect 24216 11772 24268 11824
rect 24400 11772 24452 11824
rect 21088 11704 21140 11756
rect 12716 11679 12768 11688
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 12992 11679 13044 11688
rect 12992 11645 13001 11679
rect 13001 11645 13035 11679
rect 13035 11645 13044 11679
rect 12992 11636 13044 11645
rect 13728 11636 13780 11688
rect 18604 11679 18656 11688
rect 18604 11645 18622 11679
rect 18622 11645 18656 11679
rect 18604 11636 18656 11645
rect 19340 11636 19392 11688
rect 20444 11679 20496 11688
rect 12532 11568 12584 11620
rect 13544 11568 13596 11620
rect 7564 11500 7616 11509
rect 8760 11500 8812 11552
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 18328 11611 18380 11620
rect 13820 11500 13872 11509
rect 14832 11500 14884 11552
rect 15476 11500 15528 11552
rect 18328 11577 18337 11611
rect 18337 11577 18371 11611
rect 18371 11577 18380 11611
rect 20444 11645 20453 11679
rect 20453 11645 20487 11679
rect 20487 11645 20496 11679
rect 20444 11636 20496 11645
rect 20812 11636 20864 11688
rect 18328 11568 18380 11577
rect 16212 11500 16264 11552
rect 17868 11500 17920 11552
rect 19340 11500 19392 11552
rect 21364 11500 21416 11552
rect 22100 11611 22152 11620
rect 22100 11577 22109 11611
rect 22109 11577 22143 11611
rect 22143 11577 22152 11611
rect 22100 11568 22152 11577
rect 22284 11568 22336 11620
rect 23112 11568 23164 11620
rect 23480 11500 23532 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 10048 11339 10100 11348
rect 10048 11305 10057 11339
rect 10057 11305 10091 11339
rect 10091 11305 10100 11339
rect 10048 11296 10100 11305
rect 10784 11339 10836 11348
rect 10784 11305 10793 11339
rect 10793 11305 10827 11339
rect 10827 11305 10836 11339
rect 10784 11296 10836 11305
rect 12348 11296 12400 11348
rect 16212 11339 16264 11348
rect 16212 11305 16221 11339
rect 16221 11305 16255 11339
rect 16255 11305 16264 11339
rect 16212 11296 16264 11305
rect 19340 11296 19392 11348
rect 19984 11296 20036 11348
rect 22560 11339 22612 11348
rect 11520 11271 11572 11280
rect 11520 11237 11529 11271
rect 11529 11237 11563 11271
rect 11563 11237 11572 11271
rect 11520 11228 11572 11237
rect 12440 11228 12492 11280
rect 12716 11228 12768 11280
rect 13544 11228 13596 11280
rect 15476 11228 15528 11280
rect 21180 11271 21232 11280
rect 21180 11237 21189 11271
rect 21189 11237 21223 11271
rect 21223 11237 21232 11271
rect 21180 11228 21232 11237
rect 22560 11305 22569 11339
rect 22569 11305 22603 11339
rect 22603 11305 22612 11339
rect 22560 11296 22612 11305
rect 24124 11339 24176 11348
rect 24124 11305 24133 11339
rect 24133 11305 24167 11339
rect 24167 11305 24176 11339
rect 24124 11296 24176 11305
rect 24400 11339 24452 11348
rect 24400 11305 24409 11339
rect 24409 11305 24443 11339
rect 24443 11305 24452 11339
rect 24400 11296 24452 11305
rect 21824 11228 21876 11280
rect 22836 11228 22888 11280
rect 23112 11228 23164 11280
rect 23204 11228 23256 11280
rect 24032 11228 24084 11280
rect 7288 10999 7340 11008
rect 7288 10965 7297 10999
rect 7297 10965 7331 10999
rect 7331 10965 7340 10999
rect 7288 10956 7340 10965
rect 7472 10956 7524 11008
rect 8944 11160 8996 11212
rect 10324 11203 10376 11212
rect 7748 11135 7800 11144
rect 7748 11101 7757 11135
rect 7757 11101 7791 11135
rect 7791 11101 7800 11135
rect 7748 11092 7800 11101
rect 10324 11169 10333 11203
rect 10333 11169 10367 11203
rect 10367 11169 10376 11203
rect 10324 11160 10376 11169
rect 11152 11092 11204 11144
rect 11888 11092 11940 11144
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 13728 11160 13780 11212
rect 15292 11203 15344 11212
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 15292 11160 15344 11169
rect 17500 11203 17552 11212
rect 17500 11169 17509 11203
rect 17509 11169 17543 11203
rect 17543 11169 17552 11203
rect 17500 11160 17552 11169
rect 17960 11203 18012 11212
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 18512 11160 18564 11212
rect 19248 11160 19300 11212
rect 24676 11160 24728 11212
rect 25044 11160 25096 11212
rect 15384 11092 15436 11144
rect 16028 11092 16080 11144
rect 18236 11135 18288 11144
rect 18236 11101 18245 11135
rect 18245 11101 18279 11135
rect 18279 11101 18288 11135
rect 18236 11092 18288 11101
rect 20720 11092 20772 11144
rect 21088 11135 21140 11144
rect 21088 11101 21097 11135
rect 21097 11101 21131 11135
rect 21131 11101 21140 11135
rect 21088 11092 21140 11101
rect 22284 11092 22336 11144
rect 9128 10956 9180 11008
rect 9956 10956 10008 11008
rect 10876 10956 10928 11008
rect 13360 10956 13412 11008
rect 15844 11024 15896 11076
rect 14280 10999 14332 11008
rect 14280 10965 14289 10999
rect 14289 10965 14323 10999
rect 14323 10965 14332 10999
rect 14280 10956 14332 10965
rect 15752 10956 15804 11008
rect 19984 10999 20036 11008
rect 19984 10965 19993 10999
rect 19993 10965 20027 10999
rect 20027 10965 20036 10999
rect 19984 10956 20036 10965
rect 22100 10999 22152 11008
rect 22100 10965 22109 10999
rect 22109 10965 22143 10999
rect 22143 10965 22152 10999
rect 22100 10956 22152 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2780 10752 2832 10804
rect 11520 10795 11572 10804
rect 11520 10761 11529 10795
rect 11529 10761 11563 10795
rect 11563 10761 11572 10795
rect 11520 10752 11572 10761
rect 13544 10752 13596 10804
rect 14832 10795 14884 10804
rect 14832 10761 14841 10795
rect 14841 10761 14875 10795
rect 14875 10761 14884 10795
rect 14832 10752 14884 10761
rect 17500 10752 17552 10804
rect 19984 10752 20036 10804
rect 21180 10752 21232 10804
rect 22192 10752 22244 10804
rect 23112 10752 23164 10804
rect 24676 10795 24728 10804
rect 24676 10761 24685 10795
rect 24685 10761 24719 10795
rect 24719 10761 24728 10795
rect 24676 10752 24728 10761
rect 25412 10795 25464 10804
rect 25412 10761 25421 10795
rect 25421 10761 25455 10795
rect 25455 10761 25464 10795
rect 25412 10752 25464 10761
rect 8484 10684 8536 10736
rect 21824 10727 21876 10736
rect 21824 10693 21833 10727
rect 21833 10693 21867 10727
rect 21867 10693 21876 10727
rect 21824 10684 21876 10693
rect 8024 10616 8076 10668
rect 8576 10616 8628 10668
rect 10324 10616 10376 10668
rect 10876 10659 10928 10668
rect 7472 10548 7524 10600
rect 10876 10625 10885 10659
rect 10885 10625 10919 10659
rect 10919 10625 10928 10659
rect 10876 10616 10928 10625
rect 7288 10480 7340 10532
rect 8208 10480 8260 10532
rect 9036 10480 9088 10532
rect 12532 10548 12584 10600
rect 14280 10616 14332 10668
rect 15752 10659 15804 10668
rect 15752 10625 15761 10659
rect 15761 10625 15795 10659
rect 15795 10625 15804 10659
rect 15752 10616 15804 10625
rect 16028 10659 16080 10668
rect 16028 10625 16037 10659
rect 16037 10625 16071 10659
rect 16071 10625 16080 10659
rect 16028 10616 16080 10625
rect 18052 10659 18104 10668
rect 18052 10625 18061 10659
rect 18061 10625 18095 10659
rect 18095 10625 18104 10659
rect 18052 10616 18104 10625
rect 18144 10616 18196 10668
rect 19984 10616 20036 10668
rect 20904 10616 20956 10668
rect 22008 10616 22060 10668
rect 10784 10480 10836 10532
rect 11336 10480 11388 10532
rect 12624 10480 12676 10532
rect 13544 10480 13596 10532
rect 8484 10455 8536 10464
rect 8484 10421 8493 10455
rect 8493 10421 8527 10455
rect 8527 10421 8536 10455
rect 8484 10412 8536 10421
rect 11152 10455 11204 10464
rect 11152 10421 11161 10455
rect 11161 10421 11195 10455
rect 11195 10421 11204 10455
rect 11152 10412 11204 10421
rect 11888 10455 11940 10464
rect 11888 10421 11897 10455
rect 11897 10421 11931 10455
rect 11931 10421 11940 10455
rect 11888 10412 11940 10421
rect 13452 10455 13504 10464
rect 13452 10421 13461 10455
rect 13461 10421 13495 10455
rect 13495 10421 13504 10455
rect 13452 10412 13504 10421
rect 15844 10523 15896 10532
rect 15844 10489 15853 10523
rect 15853 10489 15887 10523
rect 15887 10489 15896 10523
rect 15844 10480 15896 10489
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 17960 10412 18012 10464
rect 18144 10412 18196 10464
rect 18696 10455 18748 10464
rect 18696 10421 18705 10455
rect 18705 10421 18739 10455
rect 18739 10421 18748 10455
rect 19340 10480 19392 10532
rect 18696 10412 18748 10421
rect 22376 10548 22428 10600
rect 22744 10548 22796 10600
rect 21272 10523 21324 10532
rect 21272 10489 21281 10523
rect 21281 10489 21315 10523
rect 21315 10489 21324 10523
rect 21272 10480 21324 10489
rect 22284 10412 22336 10464
rect 23296 10412 23348 10464
rect 24124 10591 24176 10600
rect 24124 10557 24133 10591
rect 24133 10557 24167 10591
rect 24167 10557 24176 10591
rect 24124 10548 24176 10557
rect 25228 10591 25280 10600
rect 25228 10557 25237 10591
rect 25237 10557 25271 10591
rect 25271 10557 25280 10591
rect 25228 10548 25280 10557
rect 23756 10455 23808 10464
rect 23756 10421 23765 10455
rect 23765 10421 23799 10455
rect 23799 10421 23808 10455
rect 23756 10412 23808 10421
rect 25044 10455 25096 10464
rect 25044 10421 25053 10455
rect 25053 10421 25087 10455
rect 25087 10421 25096 10455
rect 25044 10412 25096 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 7748 10208 7800 10260
rect 12900 10208 12952 10260
rect 13084 10251 13136 10260
rect 13084 10217 13093 10251
rect 13093 10217 13127 10251
rect 13127 10217 13136 10251
rect 13084 10208 13136 10217
rect 15292 10208 15344 10260
rect 18236 10208 18288 10260
rect 19248 10208 19300 10260
rect 19984 10251 20036 10260
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 20720 10251 20772 10260
rect 20720 10217 20729 10251
rect 20729 10217 20763 10251
rect 20763 10217 20772 10251
rect 20720 10208 20772 10217
rect 21272 10208 21324 10260
rect 23204 10208 23256 10260
rect 5448 10183 5500 10192
rect 5448 10149 5457 10183
rect 5457 10149 5491 10183
rect 5491 10149 5500 10183
rect 5448 10140 5500 10149
rect 1492 10072 1544 10124
rect 3976 10072 4028 10124
rect 5356 10047 5408 10056
rect 5356 10013 5365 10047
rect 5365 10013 5399 10047
rect 5399 10013 5408 10047
rect 5356 10004 5408 10013
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 11888 10140 11940 10192
rect 14280 10140 14332 10192
rect 7748 10115 7800 10124
rect 7748 10081 7757 10115
rect 7757 10081 7791 10115
rect 7791 10081 7800 10115
rect 7748 10072 7800 10081
rect 7932 10115 7984 10124
rect 7932 10081 7941 10115
rect 7941 10081 7975 10115
rect 7975 10081 7984 10115
rect 7932 10072 7984 10081
rect 9036 10072 9088 10124
rect 7104 9868 7156 9920
rect 8852 10004 8904 10056
rect 10692 10072 10744 10124
rect 12532 10115 12584 10124
rect 10048 10047 10100 10056
rect 10048 10013 10057 10047
rect 10057 10013 10091 10047
rect 10091 10013 10100 10047
rect 10048 10004 10100 10013
rect 12072 10004 12124 10056
rect 12532 10081 12541 10115
rect 12541 10081 12575 10115
rect 12575 10081 12584 10115
rect 12532 10072 12584 10081
rect 13636 10115 13688 10124
rect 13636 10081 13645 10115
rect 13645 10081 13679 10115
rect 13679 10081 13688 10115
rect 13636 10072 13688 10081
rect 13728 10072 13780 10124
rect 15936 10115 15988 10124
rect 15936 10081 15945 10115
rect 15945 10081 15979 10115
rect 15979 10081 15988 10115
rect 15936 10072 15988 10081
rect 20996 10140 21048 10192
rect 16580 10072 16632 10124
rect 17500 10072 17552 10124
rect 18144 10072 18196 10124
rect 19156 10072 19208 10124
rect 23296 10140 23348 10192
rect 22928 10115 22980 10124
rect 22928 10081 22937 10115
rect 22937 10081 22971 10115
rect 22971 10081 22980 10115
rect 22928 10072 22980 10081
rect 14096 10004 14148 10056
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 16212 10047 16264 10056
rect 16212 10013 16221 10047
rect 16221 10013 16255 10047
rect 16255 10013 16264 10047
rect 16212 10004 16264 10013
rect 19432 10004 19484 10056
rect 20812 10004 20864 10056
rect 8944 9936 8996 9988
rect 12532 9936 12584 9988
rect 20260 9936 20312 9988
rect 21548 9979 21600 9988
rect 21548 9945 21557 9979
rect 21557 9945 21591 9979
rect 21591 9945 21600 9979
rect 21548 9936 21600 9945
rect 24124 10208 24176 10260
rect 9036 9911 9088 9920
rect 9036 9877 9045 9911
rect 9045 9877 9079 9911
rect 9079 9877 9088 9911
rect 9036 9868 9088 9877
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 9956 9911 10008 9920
rect 9956 9877 9965 9911
rect 9965 9877 9999 9911
rect 9999 9877 10008 9911
rect 9956 9868 10008 9877
rect 10600 9868 10652 9920
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 16856 9868 16908 9920
rect 23204 9868 23256 9920
rect 23388 9868 23440 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 3976 9707 4028 9716
rect 3976 9673 3985 9707
rect 3985 9673 4019 9707
rect 4019 9673 4028 9707
rect 3976 9664 4028 9673
rect 5356 9664 5408 9716
rect 7564 9707 7616 9716
rect 7564 9673 7573 9707
rect 7573 9673 7607 9707
rect 7607 9673 7616 9707
rect 7564 9664 7616 9673
rect 7932 9664 7984 9716
rect 9680 9707 9732 9716
rect 9680 9673 9689 9707
rect 9689 9673 9723 9707
rect 9723 9673 9732 9707
rect 9680 9664 9732 9673
rect 12440 9664 12492 9716
rect 12624 9664 12676 9716
rect 8944 9596 8996 9648
rect 9588 9596 9640 9648
rect 4068 9528 4120 9580
rect 8208 9528 8260 9580
rect 9404 9571 9456 9580
rect 9404 9537 9413 9571
rect 9413 9537 9447 9571
rect 9447 9537 9456 9571
rect 10600 9596 10652 9648
rect 15568 9664 15620 9716
rect 20996 9664 21048 9716
rect 22100 9664 22152 9716
rect 23296 9707 23348 9716
rect 23296 9673 23305 9707
rect 23305 9673 23339 9707
rect 23339 9673 23348 9707
rect 23296 9664 23348 9673
rect 15936 9596 15988 9648
rect 21272 9596 21324 9648
rect 22192 9639 22244 9648
rect 22192 9605 22201 9639
rect 22201 9605 22235 9639
rect 22235 9605 22244 9639
rect 22192 9596 22244 9605
rect 22928 9596 22980 9648
rect 9404 9528 9456 9537
rect 9956 9528 10008 9580
rect 11060 9528 11112 9580
rect 11428 9571 11480 9580
rect 11428 9537 11437 9571
rect 11437 9537 11471 9571
rect 11471 9537 11480 9571
rect 11428 9528 11480 9537
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 15752 9528 15804 9580
rect 16028 9571 16080 9580
rect 16028 9537 16037 9571
rect 16037 9537 16071 9571
rect 16071 9537 16080 9571
rect 16028 9528 16080 9537
rect 18236 9528 18288 9580
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 21180 9571 21232 9580
rect 21180 9537 21189 9571
rect 21189 9537 21223 9571
rect 21223 9537 21232 9571
rect 21180 9528 21232 9537
rect 4252 9503 4304 9512
rect 4252 9469 4270 9503
rect 4270 9469 4304 9503
rect 4252 9460 4304 9469
rect 5356 9435 5408 9444
rect 5356 9401 5365 9435
rect 5365 9401 5399 9435
rect 5399 9401 5408 9435
rect 5356 9392 5408 9401
rect 6276 9392 6328 9444
rect 9312 9460 9364 9512
rect 10692 9503 10744 9512
rect 10692 9469 10701 9503
rect 10701 9469 10735 9503
rect 10735 9469 10744 9503
rect 10692 9460 10744 9469
rect 10968 9503 11020 9512
rect 10968 9469 10977 9503
rect 10977 9469 11011 9503
rect 11011 9469 11020 9503
rect 10968 9460 11020 9469
rect 14004 9503 14056 9512
rect 14004 9469 14013 9503
rect 14013 9469 14047 9503
rect 14047 9469 14056 9503
rect 14004 9460 14056 9469
rect 22100 9460 22152 9512
rect 25228 9460 25280 9512
rect 9036 9435 9088 9444
rect 9036 9401 9045 9435
rect 9045 9401 9079 9435
rect 9079 9401 9088 9435
rect 9036 9392 9088 9401
rect 12808 9392 12860 9444
rect 13360 9392 13412 9444
rect 15568 9392 15620 9444
rect 16580 9435 16632 9444
rect 16580 9401 16589 9435
rect 16589 9401 16623 9435
rect 16623 9401 16632 9435
rect 16580 9392 16632 9401
rect 18144 9392 18196 9444
rect 20996 9435 21048 9444
rect 20996 9401 21005 9435
rect 21005 9401 21039 9435
rect 21039 9401 21048 9435
rect 20996 9392 21048 9401
rect 1492 9324 1544 9376
rect 7104 9367 7156 9376
rect 7104 9333 7113 9367
rect 7113 9333 7147 9367
rect 7147 9333 7156 9367
rect 7104 9324 7156 9333
rect 8484 9324 8536 9376
rect 9588 9324 9640 9376
rect 10048 9367 10100 9376
rect 10048 9333 10057 9367
rect 10057 9333 10091 9367
rect 10091 9333 10100 9367
rect 10048 9324 10100 9333
rect 10968 9324 11020 9376
rect 12900 9324 12952 9376
rect 13728 9324 13780 9376
rect 14188 9367 14240 9376
rect 14188 9333 14197 9367
rect 14197 9333 14231 9367
rect 14231 9333 14240 9367
rect 14188 9324 14240 9333
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 18696 9367 18748 9376
rect 18696 9333 18705 9367
rect 18705 9333 18739 9367
rect 18739 9333 18748 9367
rect 18696 9324 18748 9333
rect 20812 9324 20864 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 7748 9120 7800 9172
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 11612 9120 11664 9172
rect 12072 9120 12124 9172
rect 13636 9120 13688 9172
rect 13820 9120 13872 9172
rect 15752 9120 15804 9172
rect 19432 9120 19484 9172
rect 6184 9052 6236 9104
rect 12900 9052 12952 9104
rect 13176 9095 13228 9104
rect 13176 9061 13185 9095
rect 13185 9061 13219 9095
rect 13219 9061 13228 9095
rect 13176 9052 13228 9061
rect 15384 9052 15436 9104
rect 15844 9052 15896 9104
rect 19616 9052 19668 9104
rect 20628 9052 20680 9104
rect 7472 9027 7524 9036
rect 7472 8993 7481 9027
rect 7481 8993 7515 9027
rect 7515 8993 7524 9027
rect 7472 8984 7524 8993
rect 9036 8984 9088 9036
rect 9496 8984 9548 9036
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 9312 8916 9364 8968
rect 10140 8984 10192 9036
rect 11612 9027 11664 9036
rect 11612 8993 11621 9027
rect 11621 8993 11655 9027
rect 11655 8993 11664 9027
rect 11612 8984 11664 8993
rect 11796 9027 11848 9036
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 14372 8984 14424 9036
rect 15476 8984 15528 9036
rect 17040 9027 17092 9036
rect 17040 8993 17049 9027
rect 17049 8993 17083 9027
rect 17083 8993 17092 9027
rect 17040 8984 17092 8993
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 12072 8959 12124 8968
rect 12072 8925 12081 8959
rect 12081 8925 12115 8959
rect 12115 8925 12124 8959
rect 12072 8916 12124 8925
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 13360 8959 13412 8968
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 18604 8916 18656 8968
rect 20996 8959 21048 8968
rect 20996 8925 21005 8959
rect 21005 8925 21039 8959
rect 21039 8925 21048 8959
rect 20996 8916 21048 8925
rect 5356 8848 5408 8900
rect 7472 8848 7524 8900
rect 13912 8848 13964 8900
rect 14096 8891 14148 8900
rect 14096 8857 14105 8891
rect 14105 8857 14139 8891
rect 14139 8857 14148 8891
rect 14096 8848 14148 8857
rect 6920 8780 6972 8832
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 9496 8823 9548 8832
rect 9496 8789 9505 8823
rect 9505 8789 9539 8823
rect 9539 8789 9548 8823
rect 9496 8780 9548 8789
rect 9588 8780 9640 8832
rect 10784 8780 10836 8832
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 16304 8780 16356 8832
rect 18144 8780 18196 8832
rect 19340 8823 19392 8832
rect 19340 8789 19349 8823
rect 19349 8789 19383 8823
rect 19383 8789 19392 8823
rect 19340 8780 19392 8789
rect 19616 8823 19668 8832
rect 19616 8789 19625 8823
rect 19625 8789 19659 8823
rect 19659 8789 19668 8823
rect 19616 8780 19668 8789
rect 21180 8848 21232 8900
rect 23388 8780 23440 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 9496 8576 9548 8628
rect 11612 8576 11664 8628
rect 12808 8576 12860 8628
rect 15568 8576 15620 8628
rect 20812 8576 20864 8628
rect 20996 8619 21048 8628
rect 20996 8585 21005 8619
rect 21005 8585 21039 8619
rect 21039 8585 21048 8619
rect 20996 8576 21048 8585
rect 24768 8619 24820 8628
rect 24768 8585 24777 8619
rect 24777 8585 24811 8619
rect 24811 8585 24820 8619
rect 24768 8576 24820 8585
rect 848 8508 900 8560
rect 7104 8508 7156 8560
rect 9036 8508 9088 8560
rect 4528 8440 4580 8492
rect 5264 8483 5316 8492
rect 5264 8449 5273 8483
rect 5273 8449 5307 8483
rect 5307 8449 5316 8483
rect 5264 8440 5316 8449
rect 6000 8440 6052 8492
rect 6276 8440 6328 8492
rect 7012 8440 7064 8492
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 8852 8372 8904 8424
rect 9956 8440 10008 8492
rect 12072 8440 12124 8492
rect 14096 8440 14148 8492
rect 17040 8440 17092 8492
rect 6920 8347 6972 8356
rect 6184 8279 6236 8288
rect 6184 8245 6193 8279
rect 6193 8245 6227 8279
rect 6227 8245 6236 8279
rect 6184 8236 6236 8245
rect 6920 8313 6929 8347
rect 6929 8313 6963 8347
rect 6963 8313 6972 8347
rect 6920 8304 6972 8313
rect 7288 8304 7340 8356
rect 8024 8304 8076 8356
rect 8484 8304 8536 8356
rect 13084 8372 13136 8424
rect 14832 8372 14884 8424
rect 16764 8415 16816 8424
rect 16764 8381 16782 8415
rect 16782 8381 16816 8415
rect 19432 8440 19484 8492
rect 19984 8440 20036 8492
rect 16764 8372 16816 8381
rect 18788 8415 18840 8424
rect 18788 8381 18797 8415
rect 18797 8381 18831 8415
rect 18831 8381 18840 8415
rect 18788 8372 18840 8381
rect 23848 8372 23900 8424
rect 8668 8279 8720 8288
rect 8668 8245 8677 8279
rect 8677 8245 8711 8279
rect 8711 8245 8720 8279
rect 8668 8236 8720 8245
rect 10784 8236 10836 8288
rect 11244 8236 11296 8288
rect 11796 8279 11848 8288
rect 11796 8245 11805 8279
rect 11805 8245 11839 8279
rect 11839 8245 11848 8279
rect 11796 8236 11848 8245
rect 12072 8236 12124 8288
rect 15844 8236 15896 8288
rect 17776 8304 17828 8356
rect 18696 8304 18748 8356
rect 19616 8304 19668 8356
rect 21180 8347 21232 8356
rect 21180 8313 21189 8347
rect 21189 8313 21223 8347
rect 21223 8313 21232 8347
rect 21180 8304 21232 8313
rect 21272 8347 21324 8356
rect 21272 8313 21281 8347
rect 21281 8313 21315 8347
rect 21315 8313 21324 8347
rect 21272 8304 21324 8313
rect 16396 8236 16448 8288
rect 20628 8279 20680 8288
rect 20628 8245 20637 8279
rect 20637 8245 20671 8279
rect 20671 8245 20680 8279
rect 20628 8236 20680 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 5264 8075 5316 8084
rect 5264 8041 5273 8075
rect 5273 8041 5307 8075
rect 5307 8041 5316 8075
rect 5264 8032 5316 8041
rect 6920 8032 6972 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 10140 8032 10192 8084
rect 13176 8032 13228 8084
rect 15476 8075 15528 8084
rect 15476 8041 15485 8075
rect 15485 8041 15519 8075
rect 15519 8041 15528 8075
rect 15476 8032 15528 8041
rect 18788 8032 18840 8084
rect 22376 8032 22428 8084
rect 6276 8007 6328 8016
rect 6276 7973 6285 8007
rect 6285 7973 6319 8007
rect 6319 7973 6328 8007
rect 6276 7964 6328 7973
rect 6644 8007 6696 8016
rect 6644 7973 6653 8007
rect 6653 7973 6687 8007
rect 6687 7973 6696 8007
rect 6644 7964 6696 7973
rect 6092 7896 6144 7948
rect 8576 7896 8628 7948
rect 10048 7964 10100 8016
rect 10140 7896 10192 7948
rect 10692 7896 10744 7948
rect 12072 7964 12124 8016
rect 15844 7964 15896 8016
rect 19340 7964 19392 8016
rect 19984 8007 20036 8016
rect 19984 7973 19993 8007
rect 19993 7973 20027 8007
rect 20027 7973 20036 8007
rect 19984 7964 20036 7973
rect 20628 7964 20680 8016
rect 21364 7964 21416 8016
rect 10876 7896 10928 7948
rect 14096 7939 14148 7948
rect 14096 7905 14105 7939
rect 14105 7905 14139 7939
rect 14139 7905 14148 7939
rect 14096 7896 14148 7905
rect 16212 7939 16264 7948
rect 16212 7905 16221 7939
rect 16221 7905 16255 7939
rect 16255 7905 16264 7939
rect 16212 7896 16264 7905
rect 16948 7896 17000 7948
rect 17776 7896 17828 7948
rect 22468 7939 22520 7948
rect 22468 7905 22477 7939
rect 22477 7905 22511 7939
rect 22511 7905 22520 7939
rect 22468 7896 22520 7905
rect 6000 7828 6052 7880
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 11244 7871 11296 7880
rect 11244 7837 11253 7871
rect 11253 7837 11287 7871
rect 11287 7837 11296 7871
rect 11244 7828 11296 7837
rect 12348 7871 12400 7880
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 19984 7828 20036 7880
rect 20996 7871 21048 7880
rect 20996 7837 21005 7871
rect 21005 7837 21039 7871
rect 21039 7837 21048 7871
rect 20996 7828 21048 7837
rect 5540 7760 5592 7812
rect 8668 7760 8720 7812
rect 10600 7803 10652 7812
rect 10600 7769 10609 7803
rect 10609 7769 10643 7803
rect 10643 7769 10652 7803
rect 10600 7760 10652 7769
rect 17408 7760 17460 7812
rect 8208 7692 8260 7744
rect 8852 7692 8904 7744
rect 12440 7692 12492 7744
rect 14740 7692 14792 7744
rect 14832 7692 14884 7744
rect 16028 7735 16080 7744
rect 16028 7701 16037 7735
rect 16037 7701 16071 7735
rect 16071 7701 16080 7735
rect 16028 7692 16080 7701
rect 17132 7735 17184 7744
rect 17132 7701 17141 7735
rect 17141 7701 17175 7735
rect 17175 7701 17184 7735
rect 17132 7692 17184 7701
rect 17500 7692 17552 7744
rect 18604 7692 18656 7744
rect 21272 7692 21324 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 6092 7488 6144 7540
rect 6276 7488 6328 7540
rect 8576 7488 8628 7540
rect 13728 7531 13780 7540
rect 13728 7497 13737 7531
rect 13737 7497 13771 7531
rect 13771 7497 13780 7531
rect 13728 7488 13780 7497
rect 1584 7463 1636 7472
rect 1584 7429 1593 7463
rect 1593 7429 1627 7463
rect 1627 7429 1636 7463
rect 1584 7420 1636 7429
rect 14096 7463 14148 7472
rect 14096 7429 14105 7463
rect 14105 7429 14139 7463
rect 14139 7429 14148 7463
rect 14096 7420 14148 7429
rect 6644 7352 6696 7404
rect 7012 7352 7064 7404
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 7564 7216 7616 7268
rect 8852 7216 8904 7268
rect 10968 7284 11020 7336
rect 12164 7352 12216 7404
rect 11244 7284 11296 7336
rect 12440 7327 12492 7336
rect 8392 7191 8444 7200
rect 8392 7157 8401 7191
rect 8401 7157 8435 7191
rect 8435 7157 8444 7191
rect 8392 7148 8444 7157
rect 8760 7191 8812 7200
rect 8760 7157 8769 7191
rect 8769 7157 8803 7191
rect 8803 7157 8812 7191
rect 10600 7216 10652 7268
rect 11520 7259 11572 7268
rect 11520 7225 11529 7259
rect 11529 7225 11563 7259
rect 11563 7225 11572 7259
rect 11520 7216 11572 7225
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 14556 7327 14608 7336
rect 14556 7293 14565 7327
rect 14565 7293 14599 7327
rect 14599 7293 14608 7327
rect 14556 7284 14608 7293
rect 16304 7488 16356 7540
rect 19340 7488 19392 7540
rect 22468 7531 22520 7540
rect 22468 7497 22477 7531
rect 22477 7497 22511 7531
rect 22511 7497 22520 7531
rect 22468 7488 22520 7497
rect 16764 7463 16816 7472
rect 16764 7429 16773 7463
rect 16773 7429 16807 7463
rect 16807 7429 16816 7463
rect 16764 7420 16816 7429
rect 21180 7420 21232 7472
rect 14832 7395 14884 7404
rect 14832 7361 14841 7395
rect 14841 7361 14875 7395
rect 14875 7361 14884 7395
rect 14832 7352 14884 7361
rect 16028 7352 16080 7404
rect 17408 7352 17460 7404
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 20352 7352 20404 7404
rect 21272 7395 21324 7404
rect 21272 7361 21281 7395
rect 21281 7361 21315 7395
rect 21315 7361 21324 7395
rect 21272 7352 21324 7361
rect 21548 7395 21600 7404
rect 21548 7361 21557 7395
rect 21557 7361 21591 7395
rect 21591 7361 21600 7395
rect 21548 7352 21600 7361
rect 17316 7284 17368 7336
rect 16304 7259 16356 7268
rect 16304 7225 16313 7259
rect 16313 7225 16347 7259
rect 16347 7225 16356 7259
rect 16304 7216 16356 7225
rect 8760 7148 8812 7157
rect 10692 7148 10744 7200
rect 11704 7148 11756 7200
rect 12164 7191 12216 7200
rect 12164 7157 12173 7191
rect 12173 7157 12207 7191
rect 12207 7157 12216 7191
rect 12164 7148 12216 7157
rect 12348 7148 12400 7200
rect 15844 7148 15896 7200
rect 16764 7148 16816 7200
rect 18144 7284 18196 7336
rect 21364 7259 21416 7268
rect 17776 7191 17828 7200
rect 17776 7157 17785 7191
rect 17785 7157 17819 7191
rect 17819 7157 17828 7191
rect 17776 7148 17828 7157
rect 19432 7191 19484 7200
rect 19432 7157 19441 7191
rect 19441 7157 19475 7191
rect 19475 7157 19484 7191
rect 21364 7225 21373 7259
rect 21373 7225 21407 7259
rect 21407 7225 21416 7259
rect 21364 7216 21416 7225
rect 19432 7148 19484 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 6000 6944 6052 6996
rect 7564 6987 7616 6996
rect 7564 6953 7573 6987
rect 7573 6953 7607 6987
rect 7607 6953 7616 6987
rect 7564 6944 7616 6953
rect 8392 6944 8444 6996
rect 8484 6987 8536 6996
rect 8484 6953 8493 6987
rect 8493 6953 8527 6987
rect 8527 6953 8536 6987
rect 8484 6944 8536 6953
rect 9220 6944 9272 6996
rect 5540 6851 5592 6860
rect 5540 6817 5549 6851
rect 5549 6817 5583 6851
rect 5583 6817 5592 6851
rect 5540 6808 5592 6817
rect 6092 6808 6144 6860
rect 7288 6876 7340 6928
rect 10968 6944 11020 6996
rect 16212 6987 16264 6996
rect 16212 6953 16221 6987
rect 16221 6953 16255 6987
rect 16255 6953 16264 6987
rect 16212 6944 16264 6953
rect 17316 6944 17368 6996
rect 21364 6944 21416 6996
rect 27620 6944 27672 6996
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 11704 6851 11756 6860
rect 11704 6817 11713 6851
rect 11713 6817 11747 6851
rect 11747 6817 11756 6851
rect 11704 6808 11756 6817
rect 12072 6808 12124 6860
rect 6368 6740 6420 6792
rect 8484 6740 8536 6792
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 16764 6876 16816 6928
rect 17132 6876 17184 6928
rect 19432 6919 19484 6928
rect 19432 6885 19441 6919
rect 19441 6885 19475 6919
rect 19475 6885 19484 6919
rect 19432 6876 19484 6885
rect 19984 6919 20036 6928
rect 19984 6885 19993 6919
rect 19993 6885 20027 6919
rect 20027 6885 20036 6919
rect 19984 6876 20036 6885
rect 21548 6876 21600 6928
rect 23664 6876 23716 6928
rect 16028 6808 16080 6860
rect 17408 6851 17460 6860
rect 17408 6817 17417 6851
rect 17417 6817 17451 6851
rect 17451 6817 17460 6851
rect 18144 6851 18196 6860
rect 17408 6808 17460 6817
rect 18144 6817 18153 6851
rect 18153 6817 18187 6851
rect 18187 6817 18196 6851
rect 18144 6808 18196 6817
rect 20904 6851 20956 6860
rect 15292 6740 15344 6792
rect 17500 6740 17552 6792
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 10140 6672 10192 6724
rect 14556 6672 14608 6724
rect 15384 6672 15436 6724
rect 15476 6672 15528 6724
rect 18972 6740 19024 6792
rect 20812 6740 20864 6792
rect 22376 6808 22428 6860
rect 24032 6808 24084 6860
rect 25504 6808 25556 6860
rect 22652 6783 22704 6792
rect 22652 6749 22661 6783
rect 22661 6749 22695 6783
rect 22695 6749 22704 6783
rect 22652 6740 22704 6749
rect 20996 6672 21048 6724
rect 5448 6604 5500 6656
rect 6000 6604 6052 6656
rect 6828 6604 6880 6656
rect 8852 6647 8904 6656
rect 8852 6613 8861 6647
rect 8861 6613 8895 6647
rect 8895 6613 8904 6647
rect 8852 6604 8904 6613
rect 17408 6604 17460 6656
rect 18788 6647 18840 6656
rect 18788 6613 18797 6647
rect 18797 6613 18831 6647
rect 18831 6613 18840 6647
rect 18788 6604 18840 6613
rect 20352 6647 20404 6656
rect 20352 6613 20361 6647
rect 20361 6613 20395 6647
rect 20395 6613 20404 6647
rect 20352 6604 20404 6613
rect 22100 6672 22152 6724
rect 23756 6604 23808 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 20 6400 72 6452
rect 16028 6443 16080 6452
rect 16028 6409 16037 6443
rect 16037 6409 16071 6443
rect 16071 6409 16080 6443
rect 16028 6400 16080 6409
rect 17132 6443 17184 6452
rect 17132 6409 17141 6443
rect 17141 6409 17175 6443
rect 17175 6409 17184 6443
rect 17132 6400 17184 6409
rect 17500 6443 17552 6452
rect 17500 6409 17509 6443
rect 17509 6409 17543 6443
rect 17543 6409 17552 6443
rect 17500 6400 17552 6409
rect 18972 6400 19024 6452
rect 19432 6443 19484 6452
rect 19432 6409 19441 6443
rect 19441 6409 19475 6443
rect 19475 6409 19484 6443
rect 19432 6400 19484 6409
rect 20904 6443 20956 6452
rect 20904 6409 20913 6443
rect 20913 6409 20947 6443
rect 20947 6409 20956 6443
rect 20904 6400 20956 6409
rect 22376 6400 22428 6452
rect 25504 6443 25556 6452
rect 25504 6409 25513 6443
rect 25513 6409 25547 6443
rect 25547 6409 25556 6443
rect 25504 6400 25556 6409
rect 6552 6264 6604 6316
rect 8760 6264 8812 6316
rect 8852 6264 8904 6316
rect 5264 6239 5316 6248
rect 5264 6205 5273 6239
rect 5273 6205 5307 6239
rect 5307 6205 5316 6239
rect 5448 6239 5500 6248
rect 5264 6196 5316 6205
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 5448 6196 5500 6205
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 6920 6239 6972 6248
rect 6920 6205 6929 6239
rect 6929 6205 6963 6239
rect 6963 6205 6972 6239
rect 7104 6239 7156 6248
rect 6920 6196 6972 6205
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 8576 6239 8628 6248
rect 8576 6205 8585 6239
rect 8585 6205 8619 6239
rect 8619 6205 8628 6239
rect 8576 6196 8628 6205
rect 9956 6264 10008 6316
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 11152 6332 11204 6384
rect 17592 6332 17644 6384
rect 18788 6332 18840 6384
rect 10784 6239 10836 6248
rect 7564 6171 7616 6180
rect 7564 6137 7573 6171
rect 7573 6137 7607 6171
rect 7607 6137 7616 6171
rect 7564 6128 7616 6137
rect 6092 6060 6144 6112
rect 7932 6103 7984 6112
rect 7932 6069 7941 6103
rect 7941 6069 7975 6103
rect 7975 6069 7984 6103
rect 7932 6060 7984 6069
rect 8484 6103 8536 6112
rect 8484 6069 8493 6103
rect 8493 6069 8527 6103
rect 8527 6069 8536 6103
rect 8484 6060 8536 6069
rect 9588 6060 9640 6112
rect 10784 6205 10793 6239
rect 10793 6205 10827 6239
rect 10827 6205 10836 6239
rect 10784 6196 10836 6205
rect 11520 6264 11572 6316
rect 13268 6307 13320 6316
rect 13268 6273 13277 6307
rect 13277 6273 13311 6307
rect 13311 6273 13320 6307
rect 13268 6264 13320 6273
rect 14740 6264 14792 6316
rect 15476 6307 15528 6316
rect 15476 6273 15485 6307
rect 15485 6273 15519 6307
rect 15519 6273 15528 6307
rect 15476 6264 15528 6273
rect 22100 6332 22152 6384
rect 22652 6264 22704 6316
rect 24216 6264 24268 6316
rect 11704 6196 11756 6248
rect 11520 6171 11572 6180
rect 11520 6137 11529 6171
rect 11529 6137 11563 6171
rect 11563 6137 11572 6171
rect 11520 6128 11572 6137
rect 15108 6128 15160 6180
rect 12072 6060 12124 6112
rect 13176 6103 13228 6112
rect 13176 6069 13185 6103
rect 13185 6069 13219 6103
rect 13219 6069 13228 6103
rect 13176 6060 13228 6069
rect 16120 6060 16172 6112
rect 16856 6196 16908 6248
rect 22468 6196 22520 6248
rect 16764 6128 16816 6180
rect 20260 6128 20312 6180
rect 20444 6171 20496 6180
rect 20444 6137 20453 6171
rect 20453 6137 20487 6171
rect 20487 6137 20496 6171
rect 20444 6128 20496 6137
rect 21364 6128 21416 6180
rect 21640 6128 21692 6180
rect 22100 6128 22152 6180
rect 22560 6060 22612 6112
rect 24032 6060 24084 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 6368 5899 6420 5908
rect 6368 5865 6377 5899
rect 6377 5865 6411 5899
rect 6411 5865 6420 5899
rect 6368 5856 6420 5865
rect 12440 5856 12492 5908
rect 13268 5899 13320 5908
rect 13268 5865 13277 5899
rect 13277 5865 13311 5899
rect 13311 5865 13320 5899
rect 13268 5856 13320 5865
rect 7104 5788 7156 5840
rect 8208 5788 8260 5840
rect 9312 5788 9364 5840
rect 12072 5788 12124 5840
rect 12256 5831 12308 5840
rect 12256 5797 12259 5831
rect 12259 5797 12293 5831
rect 12293 5797 12308 5831
rect 12256 5788 12308 5797
rect 13176 5788 13228 5840
rect 14280 5856 14332 5908
rect 14740 5856 14792 5908
rect 13820 5831 13872 5840
rect 13820 5797 13829 5831
rect 13829 5797 13863 5831
rect 13863 5797 13872 5831
rect 13820 5788 13872 5797
rect 15108 5788 15160 5840
rect 15844 5788 15896 5840
rect 17132 5788 17184 5840
rect 6552 5720 6604 5772
rect 6736 5763 6788 5772
rect 6736 5729 6745 5763
rect 6745 5729 6779 5763
rect 6779 5729 6788 5763
rect 6736 5720 6788 5729
rect 7288 5720 7340 5772
rect 7932 5720 7984 5772
rect 8300 5763 8352 5772
rect 8300 5729 8309 5763
rect 8309 5729 8343 5763
rect 8343 5729 8352 5763
rect 8300 5720 8352 5729
rect 9588 5720 9640 5772
rect 10784 5763 10836 5772
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 9220 5652 9272 5704
rect 10784 5729 10793 5763
rect 10793 5729 10827 5763
rect 10827 5729 10836 5763
rect 10784 5720 10836 5729
rect 11336 5720 11388 5772
rect 11888 5763 11940 5772
rect 11888 5729 11897 5763
rect 11897 5729 11931 5763
rect 11931 5729 11940 5763
rect 11888 5720 11940 5729
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 19524 5856 19576 5908
rect 24124 5899 24176 5908
rect 24124 5865 24133 5899
rect 24133 5865 24167 5899
rect 24167 5865 24176 5899
rect 24124 5856 24176 5865
rect 19432 5788 19484 5840
rect 21088 5831 21140 5840
rect 21088 5797 21097 5831
rect 21097 5797 21131 5831
rect 21131 5797 21140 5831
rect 21088 5788 21140 5797
rect 21640 5831 21692 5840
rect 21640 5797 21649 5831
rect 21649 5797 21683 5831
rect 21683 5797 21692 5831
rect 21640 5788 21692 5797
rect 22192 5720 22244 5772
rect 22928 5763 22980 5772
rect 22928 5729 22937 5763
rect 22937 5729 22971 5763
rect 22971 5729 22980 5763
rect 22928 5720 22980 5729
rect 23388 5720 23440 5772
rect 5264 5627 5316 5636
rect 5264 5593 5273 5627
rect 5273 5593 5307 5627
rect 5307 5593 5316 5627
rect 5264 5584 5316 5593
rect 6184 5584 6236 5636
rect 7380 5584 7432 5636
rect 8392 5584 8444 5636
rect 13912 5652 13964 5704
rect 14464 5652 14516 5704
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 20720 5652 20772 5704
rect 22560 5652 22612 5704
rect 24216 5652 24268 5704
rect 9772 5627 9824 5636
rect 9772 5593 9781 5627
rect 9781 5593 9815 5627
rect 9815 5593 9824 5627
rect 9772 5584 9824 5593
rect 18880 5584 18932 5636
rect 20260 5627 20312 5636
rect 20260 5593 20269 5627
rect 20269 5593 20303 5627
rect 20303 5593 20312 5627
rect 20260 5584 20312 5593
rect 21548 5584 21600 5636
rect 7932 5559 7984 5568
rect 7932 5525 7941 5559
rect 7941 5525 7975 5559
rect 7975 5525 7984 5559
rect 7932 5516 7984 5525
rect 12072 5516 12124 5568
rect 12808 5559 12860 5568
rect 12808 5525 12817 5559
rect 12817 5525 12851 5559
rect 12851 5525 12860 5559
rect 12808 5516 12860 5525
rect 14280 5516 14332 5568
rect 15476 5516 15528 5568
rect 16212 5559 16264 5568
rect 16212 5525 16221 5559
rect 16221 5525 16255 5559
rect 16255 5525 16264 5559
rect 16212 5516 16264 5525
rect 18696 5559 18748 5568
rect 18696 5525 18705 5559
rect 18705 5525 18739 5559
rect 18739 5525 18748 5559
rect 18696 5516 18748 5525
rect 19892 5559 19944 5568
rect 19892 5525 19901 5559
rect 19901 5525 19935 5559
rect 19935 5525 19944 5559
rect 19892 5516 19944 5525
rect 20812 5516 20864 5568
rect 21364 5516 21416 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 6184 5355 6236 5364
rect 6184 5321 6193 5355
rect 6193 5321 6227 5355
rect 6227 5321 6236 5355
rect 6184 5312 6236 5321
rect 6736 5312 6788 5364
rect 9036 5355 9088 5364
rect 9036 5321 9045 5355
rect 9045 5321 9079 5355
rect 9079 5321 9088 5355
rect 9036 5312 9088 5321
rect 13820 5312 13872 5364
rect 16212 5312 16264 5364
rect 19892 5312 19944 5364
rect 20536 5312 20588 5364
rect 23388 5355 23440 5364
rect 23388 5321 23397 5355
rect 23397 5321 23431 5355
rect 23431 5321 23440 5355
rect 23388 5312 23440 5321
rect 24216 5312 24268 5364
rect 9220 5287 9272 5296
rect 9220 5253 9229 5287
rect 9229 5253 9263 5287
rect 9263 5253 9272 5287
rect 15476 5287 15528 5296
rect 9220 5244 9272 5253
rect 15476 5253 15485 5287
rect 15485 5253 15519 5287
rect 15519 5253 15528 5287
rect 15476 5244 15528 5253
rect 15844 5287 15896 5296
rect 15844 5253 15853 5287
rect 15853 5253 15887 5287
rect 15887 5253 15896 5287
rect 15844 5244 15896 5253
rect 11520 5176 11572 5228
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 16672 5176 16724 5228
rect 18696 5244 18748 5296
rect 20444 5219 20496 5228
rect 20444 5185 20453 5219
rect 20453 5185 20487 5219
rect 20487 5185 20496 5219
rect 20444 5176 20496 5185
rect 20628 5176 20680 5228
rect 23848 5176 23900 5228
rect 8300 5108 8352 5160
rect 5448 5040 5500 5092
rect 8392 5040 8444 5092
rect 9036 5108 9088 5160
rect 9772 5108 9824 5160
rect 11336 5151 11388 5160
rect 11336 5117 11345 5151
rect 11345 5117 11379 5151
rect 11379 5117 11388 5151
rect 11336 5108 11388 5117
rect 11612 5040 11664 5092
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 7748 4972 7800 5024
rect 11796 4972 11848 5024
rect 13176 5040 13228 5092
rect 18696 5108 18748 5160
rect 14924 5083 14976 5092
rect 14924 5049 14933 5083
rect 14933 5049 14967 5083
rect 14967 5049 14976 5083
rect 14924 5040 14976 5049
rect 16488 5083 16540 5092
rect 16488 5049 16497 5083
rect 16497 5049 16531 5083
rect 16531 5049 16540 5083
rect 16488 5040 16540 5049
rect 16764 5040 16816 5092
rect 17224 5040 17276 5092
rect 18788 5040 18840 5092
rect 21916 5151 21968 5160
rect 19156 5040 19208 5092
rect 21916 5117 21925 5151
rect 21925 5117 21959 5151
rect 21959 5117 21968 5151
rect 21916 5108 21968 5117
rect 22376 5151 22428 5160
rect 22376 5117 22385 5151
rect 22385 5117 22419 5151
rect 22419 5117 22428 5151
rect 22376 5108 22428 5117
rect 23940 5108 23992 5160
rect 17132 4972 17184 5024
rect 18696 4972 18748 5024
rect 19432 4972 19484 5024
rect 20536 5083 20588 5092
rect 20536 5049 20545 5083
rect 20545 5049 20579 5083
rect 20579 5049 20588 5083
rect 20536 5040 20588 5049
rect 21272 5040 21324 5092
rect 21088 4972 21140 5024
rect 21732 5015 21784 5024
rect 21732 4981 21741 5015
rect 21741 4981 21775 5015
rect 21775 4981 21784 5015
rect 21732 4972 21784 4981
rect 22376 4972 22428 5024
rect 22928 5015 22980 5024
rect 22928 4981 22937 5015
rect 22937 4981 22971 5015
rect 22971 4981 22980 5015
rect 22928 4972 22980 4981
rect 23480 4972 23532 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 8116 4768 8168 4820
rect 11244 4768 11296 4820
rect 11888 4811 11940 4820
rect 11888 4777 11897 4811
rect 11897 4777 11931 4811
rect 11931 4777 11940 4811
rect 11888 4768 11940 4777
rect 13084 4811 13136 4820
rect 13084 4777 13093 4811
rect 13093 4777 13127 4811
rect 13127 4777 13136 4811
rect 13084 4768 13136 4777
rect 15292 4768 15344 4820
rect 16488 4811 16540 4820
rect 16488 4777 16497 4811
rect 16497 4777 16531 4811
rect 16531 4777 16540 4811
rect 16488 4768 16540 4777
rect 18512 4768 18564 4820
rect 10416 4700 10468 4752
rect 12256 4700 12308 4752
rect 12808 4700 12860 4752
rect 13452 4700 13504 4752
rect 14280 4743 14332 4752
rect 14280 4709 14289 4743
rect 14289 4709 14323 4743
rect 14323 4709 14332 4743
rect 14280 4700 14332 4709
rect 15844 4700 15896 4752
rect 17132 4700 17184 4752
rect 18880 4768 18932 4820
rect 19524 4811 19576 4820
rect 19524 4777 19533 4811
rect 19533 4777 19567 4811
rect 19567 4777 19576 4811
rect 19524 4768 19576 4777
rect 20444 4768 20496 4820
rect 20720 4811 20772 4820
rect 20720 4777 20729 4811
rect 20729 4777 20763 4811
rect 20763 4777 20772 4811
rect 20720 4768 20772 4777
rect 21916 4811 21968 4820
rect 18788 4700 18840 4752
rect 21916 4777 21925 4811
rect 21925 4777 21959 4811
rect 21959 4777 21968 4811
rect 21916 4768 21968 4777
rect 22192 4768 22244 4820
rect 22560 4811 22612 4820
rect 22560 4777 22569 4811
rect 22569 4777 22603 4811
rect 22603 4777 22612 4811
rect 22560 4768 22612 4777
rect 6552 4632 6604 4684
rect 7932 4632 7984 4684
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 9680 4675 9732 4684
rect 9680 4641 9689 4675
rect 9689 4641 9723 4675
rect 9723 4641 9732 4675
rect 9680 4632 9732 4641
rect 10140 4675 10192 4684
rect 10140 4641 10149 4675
rect 10149 4641 10183 4675
rect 10183 4641 10192 4675
rect 10140 4632 10192 4641
rect 10508 4675 10560 4684
rect 10508 4641 10517 4675
rect 10517 4641 10551 4675
rect 10551 4641 10560 4675
rect 10508 4632 10560 4641
rect 9588 4564 9640 4616
rect 11428 4632 11480 4684
rect 14924 4675 14976 4684
rect 14924 4641 14933 4675
rect 14933 4641 14967 4675
rect 14967 4641 14976 4675
rect 14924 4632 14976 4641
rect 15292 4632 15344 4684
rect 17316 4632 17368 4684
rect 20904 4675 20956 4684
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 23296 4700 23348 4752
rect 20904 4632 20956 4641
rect 11244 4564 11296 4616
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 12808 4564 12860 4616
rect 14648 4564 14700 4616
rect 18696 4564 18748 4616
rect 18880 4607 18932 4616
rect 18880 4573 18889 4607
rect 18889 4573 18923 4607
rect 18923 4573 18932 4607
rect 18880 4564 18932 4573
rect 18972 4564 19024 4616
rect 20812 4564 20864 4616
rect 21456 4632 21508 4684
rect 22836 4632 22888 4684
rect 22928 4675 22980 4684
rect 22928 4641 22937 4675
rect 22937 4641 22971 4675
rect 22971 4641 22980 4675
rect 24032 4675 24084 4684
rect 22928 4632 22980 4641
rect 24032 4641 24041 4675
rect 24041 4641 24075 4675
rect 24075 4641 24084 4675
rect 24032 4632 24084 4641
rect 25504 4632 25556 4684
rect 21732 4564 21784 4616
rect 24124 4564 24176 4616
rect 24860 4564 24912 4616
rect 7472 4496 7524 4548
rect 9772 4496 9824 4548
rect 20996 4496 21048 4548
rect 9312 4428 9364 4480
rect 9680 4428 9732 4480
rect 11520 4471 11572 4480
rect 11520 4437 11529 4471
rect 11529 4437 11563 4471
rect 11563 4437 11572 4471
rect 11520 4428 11572 4437
rect 14556 4471 14608 4480
rect 14556 4437 14565 4471
rect 14565 4437 14599 4471
rect 14599 4437 14608 4471
rect 14556 4428 14608 4437
rect 15936 4428 15988 4480
rect 17776 4428 17828 4480
rect 18604 4428 18656 4480
rect 22376 4428 22428 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 12072 4224 12124 4276
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 15752 4224 15804 4276
rect 16396 4224 16448 4276
rect 17040 4224 17092 4276
rect 17316 4224 17368 4276
rect 18512 4267 18564 4276
rect 18512 4233 18521 4267
rect 18521 4233 18555 4267
rect 18555 4233 18564 4267
rect 18512 4224 18564 4233
rect 18788 4224 18840 4276
rect 19248 4224 19300 4276
rect 20904 4224 20956 4276
rect 21732 4267 21784 4276
rect 21732 4233 21741 4267
rect 21741 4233 21775 4267
rect 21775 4233 21784 4267
rect 21732 4224 21784 4233
rect 22836 4224 22888 4276
rect 24032 4267 24084 4276
rect 24032 4233 24041 4267
rect 24041 4233 24075 4267
rect 24075 4233 24084 4267
rect 24032 4224 24084 4233
rect 25136 4267 25188 4276
rect 25136 4233 25145 4267
rect 25145 4233 25179 4267
rect 25179 4233 25188 4267
rect 25136 4224 25188 4233
rect 7472 4199 7524 4208
rect 7472 4165 7481 4199
rect 7481 4165 7515 4199
rect 7515 4165 7524 4199
rect 7472 4156 7524 4165
rect 7748 4156 7800 4208
rect 9036 4156 9088 4208
rect 16672 4156 16724 4208
rect 19524 4156 19576 4208
rect 6920 4088 6972 4140
rect 7932 4088 7984 4140
rect 9588 4088 9640 4140
rect 9680 4088 9732 4140
rect 12532 4088 12584 4140
rect 12808 4131 12860 4140
rect 12808 4097 12817 4131
rect 12817 4097 12851 4131
rect 12851 4097 12860 4131
rect 12808 4088 12860 4097
rect 13912 4088 13964 4140
rect 14556 4088 14608 4140
rect 15844 4088 15896 4140
rect 16764 4131 16816 4140
rect 16764 4097 16773 4131
rect 16773 4097 16807 4131
rect 16807 4097 16816 4131
rect 16764 4088 16816 4097
rect 18696 4088 18748 4140
rect 19064 4088 19116 4140
rect 19248 4088 19300 4140
rect 3516 3952 3568 4004
rect 6552 3995 6604 4004
rect 6552 3961 6561 3995
rect 6561 3961 6595 3995
rect 6595 3961 6604 3995
rect 6552 3952 6604 3961
rect 6828 3952 6880 4004
rect 9128 3952 9180 4004
rect 9496 4063 9548 4072
rect 9496 4029 9505 4063
rect 9505 4029 9539 4063
rect 9539 4029 9548 4063
rect 10140 4063 10192 4072
rect 9496 4020 9548 4029
rect 10140 4029 10149 4063
rect 10149 4029 10183 4063
rect 10183 4029 10192 4063
rect 10140 4020 10192 4029
rect 10508 4063 10560 4072
rect 10508 4029 10517 4063
rect 10517 4029 10551 4063
rect 10551 4029 10560 4063
rect 10508 4020 10560 4029
rect 10876 4063 10928 4072
rect 10876 4029 10885 4063
rect 10885 4029 10919 4063
rect 10919 4029 10928 4063
rect 10876 4020 10928 4029
rect 16396 4020 16448 4072
rect 21456 4088 21508 4140
rect 22560 4088 22612 4140
rect 25504 4131 25556 4140
rect 25504 4097 25513 4131
rect 25513 4097 25547 4131
rect 25547 4097 25556 4131
rect 25504 4088 25556 4097
rect 27068 4088 27120 4140
rect 25136 4020 25188 4072
rect 25872 4020 25924 4072
rect 9864 3884 9916 3936
rect 12348 3952 12400 4004
rect 10692 3884 10744 3936
rect 11428 3884 11480 3936
rect 12440 3884 12492 3936
rect 12624 3995 12676 4004
rect 12624 3961 12633 3995
rect 12633 3961 12667 3995
rect 12667 3961 12676 3995
rect 12624 3952 12676 3961
rect 14372 3952 14424 4004
rect 15660 3995 15712 4004
rect 15660 3961 15669 3995
rect 15669 3961 15703 3995
rect 15703 3961 15712 3995
rect 15660 3952 15712 3961
rect 15752 3995 15804 4004
rect 15752 3961 15761 3995
rect 15761 3961 15795 3995
rect 15795 3961 15804 3995
rect 15752 3952 15804 3961
rect 15936 3952 15988 4004
rect 18420 3952 18472 4004
rect 18880 3952 18932 4004
rect 19156 3952 19208 4004
rect 17960 3884 18012 3936
rect 19984 3884 20036 3936
rect 20628 3884 20680 3936
rect 22192 3884 22244 3936
rect 25504 3884 25556 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 7932 3680 7984 3732
rect 9864 3680 9916 3732
rect 10876 3680 10928 3732
rect 12440 3680 12492 3732
rect 17960 3723 18012 3732
rect 17960 3689 17969 3723
rect 17969 3689 18003 3723
rect 18003 3689 18012 3723
rect 17960 3680 18012 3689
rect 19064 3723 19116 3732
rect 19064 3689 19073 3723
rect 19073 3689 19107 3723
rect 19107 3689 19116 3723
rect 19064 3680 19116 3689
rect 9404 3655 9456 3664
rect 9404 3621 9413 3655
rect 9413 3621 9447 3655
rect 9447 3621 9456 3655
rect 13728 3655 13780 3664
rect 9404 3612 9456 3621
rect 13728 3621 13737 3655
rect 13737 3621 13771 3655
rect 13771 3621 13780 3655
rect 13728 3612 13780 3621
rect 15476 3655 15528 3664
rect 6276 3544 6328 3596
rect 7012 3544 7064 3596
rect 8944 3544 8996 3596
rect 9312 3544 9364 3596
rect 9496 3544 9548 3596
rect 10140 3544 10192 3596
rect 10600 3587 10652 3596
rect 10048 3476 10100 3528
rect 10600 3553 10609 3587
rect 10609 3553 10643 3587
rect 10643 3553 10652 3587
rect 10600 3544 10652 3553
rect 11428 3544 11480 3596
rect 11980 3587 12032 3596
rect 11980 3553 11989 3587
rect 11989 3553 12023 3587
rect 12023 3553 12032 3587
rect 11980 3544 12032 3553
rect 12348 3544 12400 3596
rect 14188 3544 14240 3596
rect 15476 3621 15485 3655
rect 15485 3621 15519 3655
rect 15519 3621 15528 3655
rect 15476 3612 15528 3621
rect 16028 3655 16080 3664
rect 16028 3621 16037 3655
rect 16037 3621 16071 3655
rect 16071 3621 16080 3655
rect 16028 3612 16080 3621
rect 11152 3519 11204 3528
rect 8208 3408 8260 3460
rect 11152 3485 11161 3519
rect 11161 3485 11195 3519
rect 11195 3485 11204 3519
rect 11152 3476 11204 3485
rect 12256 3476 12308 3528
rect 12716 3408 12768 3460
rect 15660 3476 15712 3528
rect 19524 3612 19576 3664
rect 22192 3680 22244 3732
rect 22284 3680 22336 3732
rect 20996 3655 21048 3664
rect 20996 3621 21005 3655
rect 21005 3621 21039 3655
rect 21039 3621 21048 3655
rect 20996 3612 21048 3621
rect 21180 3612 21232 3664
rect 21732 3612 21784 3664
rect 25504 3612 25556 3664
rect 22468 3587 22520 3596
rect 22468 3553 22477 3587
rect 22477 3553 22511 3587
rect 22511 3553 22520 3587
rect 22468 3544 22520 3553
rect 24124 3544 24176 3596
rect 24676 3544 24728 3596
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 21456 3476 21508 3528
rect 21824 3476 21876 3528
rect 15936 3408 15988 3460
rect 8024 3383 8076 3392
rect 8024 3349 8033 3383
rect 8033 3349 8067 3383
rect 8067 3349 8076 3383
rect 8024 3340 8076 3349
rect 8300 3340 8352 3392
rect 8852 3340 8904 3392
rect 9312 3340 9364 3392
rect 11520 3340 11572 3392
rect 11612 3340 11664 3392
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 12900 3383 12952 3392
rect 12900 3349 12909 3383
rect 12909 3349 12943 3383
rect 12943 3349 12952 3383
rect 12900 3340 12952 3349
rect 13268 3383 13320 3392
rect 13268 3349 13277 3383
rect 13277 3349 13311 3383
rect 13311 3349 13320 3383
rect 13268 3340 13320 3349
rect 14648 3383 14700 3392
rect 14648 3349 14657 3383
rect 14657 3349 14691 3383
rect 14691 3349 14700 3383
rect 14648 3340 14700 3349
rect 15292 3340 15344 3392
rect 16580 3340 16632 3392
rect 18512 3383 18564 3392
rect 18512 3349 18521 3383
rect 18521 3349 18555 3383
rect 18555 3349 18564 3383
rect 18512 3340 18564 3349
rect 19524 3383 19576 3392
rect 19524 3349 19533 3383
rect 19533 3349 19567 3383
rect 19567 3349 19576 3383
rect 19524 3340 19576 3349
rect 20352 3408 20404 3460
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 8944 3136 8996 3188
rect 9864 3136 9916 3188
rect 11428 3179 11480 3188
rect 11428 3145 11437 3179
rect 11437 3145 11471 3179
rect 11471 3145 11480 3179
rect 11428 3136 11480 3145
rect 11980 3179 12032 3188
rect 11980 3145 11989 3179
rect 11989 3145 12023 3179
rect 12023 3145 12032 3179
rect 11980 3136 12032 3145
rect 15476 3179 15528 3188
rect 15476 3145 15485 3179
rect 15485 3145 15519 3179
rect 15519 3145 15528 3179
rect 15476 3136 15528 3145
rect 15936 3179 15988 3188
rect 15936 3145 15945 3179
rect 15945 3145 15979 3179
rect 15979 3145 15988 3179
rect 15936 3136 15988 3145
rect 16764 3136 16816 3188
rect 17960 3136 18012 3188
rect 18512 3136 18564 3188
rect 19984 3179 20036 3188
rect 19984 3145 19993 3179
rect 19993 3145 20027 3179
rect 20027 3145 20036 3179
rect 19984 3136 20036 3145
rect 21548 3179 21600 3188
rect 21548 3145 21557 3179
rect 21557 3145 21591 3179
rect 21591 3145 21600 3179
rect 21548 3136 21600 3145
rect 23204 3136 23256 3188
rect 6184 3000 6236 3052
rect 7196 3068 7248 3120
rect 15200 3068 15252 3120
rect 9128 3000 9180 3052
rect 9312 2975 9364 2984
rect 9312 2941 9321 2975
rect 9321 2941 9355 2975
rect 9355 2941 9364 2975
rect 9312 2932 9364 2941
rect 8484 2907 8536 2916
rect 8484 2873 8493 2907
rect 8493 2873 8527 2907
rect 8527 2873 8536 2907
rect 8484 2864 8536 2873
rect 7472 2796 7524 2848
rect 7932 2796 7984 2848
rect 10600 3000 10652 3052
rect 11152 3000 11204 3052
rect 10876 2932 10928 2984
rect 11244 2932 11296 2984
rect 13268 2932 13320 2984
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 14372 2932 14424 2984
rect 16856 3068 16908 3120
rect 16580 3000 16632 3052
rect 18420 3000 18472 3052
rect 19248 3000 19300 3052
rect 20628 3068 20680 3120
rect 21088 3068 21140 3120
rect 22468 3068 22520 3120
rect 24124 3111 24176 3120
rect 24124 3077 24133 3111
rect 24133 3077 24167 3111
rect 24167 3077 24176 3111
rect 24124 3068 24176 3077
rect 21732 3043 21784 3052
rect 21732 3009 21741 3043
rect 21741 3009 21775 3043
rect 21775 3009 21784 3043
rect 21732 3000 21784 3009
rect 21824 3000 21876 3052
rect 22376 2932 22428 2984
rect 24860 2932 24912 2984
rect 10784 2907 10836 2916
rect 10784 2873 10793 2907
rect 10793 2873 10827 2907
rect 10827 2873 10836 2907
rect 10784 2864 10836 2873
rect 11428 2864 11480 2916
rect 11796 2864 11848 2916
rect 12624 2864 12676 2916
rect 13728 2864 13780 2916
rect 17776 2864 17828 2916
rect 20168 2907 20220 2916
rect 18512 2796 18564 2848
rect 20168 2873 20177 2907
rect 20177 2873 20211 2907
rect 20211 2873 20220 2907
rect 20168 2864 20220 2873
rect 19984 2796 20036 2848
rect 20536 2796 20588 2848
rect 21180 2796 21232 2848
rect 21548 2796 21600 2848
rect 23572 2796 23624 2848
rect 24676 2796 24728 2848
rect 26148 2796 26200 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 7748 2592 7800 2644
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 8484 2592 8536 2644
rect 14188 2635 14240 2644
rect 5540 2456 5592 2508
rect 9680 2524 9732 2576
rect 9036 2456 9088 2508
rect 9128 2456 9180 2508
rect 9404 2456 9456 2508
rect 11428 2524 11480 2576
rect 11612 2567 11664 2576
rect 11612 2533 11621 2567
rect 11621 2533 11655 2567
rect 11655 2533 11664 2567
rect 11612 2524 11664 2533
rect 14188 2601 14197 2635
rect 14197 2601 14231 2635
rect 14231 2601 14240 2635
rect 14188 2592 14240 2601
rect 14280 2592 14332 2644
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 17592 2635 17644 2644
rect 17592 2601 17601 2635
rect 17601 2601 17635 2635
rect 17635 2601 17644 2635
rect 17592 2592 17644 2601
rect 18788 2635 18840 2644
rect 18788 2601 18797 2635
rect 18797 2601 18831 2635
rect 18831 2601 18840 2635
rect 18788 2592 18840 2601
rect 20168 2635 20220 2644
rect 20168 2601 20177 2635
rect 20177 2601 20211 2635
rect 20211 2601 20220 2635
rect 20168 2592 20220 2601
rect 21824 2592 21876 2644
rect 20536 2524 20588 2576
rect 21272 2567 21324 2576
rect 21272 2533 21281 2567
rect 21281 2533 21315 2567
rect 21315 2533 21324 2567
rect 21272 2524 21324 2533
rect 21364 2567 21416 2576
rect 21364 2533 21373 2567
rect 21373 2533 21407 2567
rect 21407 2533 21416 2567
rect 21364 2524 21416 2533
rect 10784 2456 10836 2508
rect 16856 2456 16908 2508
rect 23572 2592 23624 2644
rect 23756 2592 23808 2644
rect 24032 2499 24084 2508
rect 24032 2465 24076 2499
rect 24076 2465 24084 2499
rect 24032 2456 24084 2465
rect 10692 2388 10744 2440
rect 5816 2320 5868 2372
rect 8576 2320 8628 2372
rect 9772 2320 9824 2372
rect 10048 2320 10100 2372
rect 13912 2388 13964 2440
rect 18788 2388 18840 2440
rect 19248 2431 19300 2440
rect 19248 2397 19257 2431
rect 19257 2397 19291 2431
rect 19291 2397 19300 2431
rect 19248 2388 19300 2397
rect 21364 2388 21416 2440
rect 21456 2388 21508 2440
rect 16120 2363 16172 2372
rect 16120 2329 16129 2363
rect 16129 2329 16163 2363
rect 16163 2329 16172 2363
rect 16120 2320 16172 2329
rect 16764 2320 16816 2372
rect 19984 2320 20036 2372
rect 21824 2363 21876 2372
rect 7288 2252 7340 2304
rect 9036 2252 9088 2304
rect 12900 2252 12952 2304
rect 16856 2295 16908 2304
rect 16856 2261 16865 2295
rect 16865 2261 16899 2295
rect 16899 2261 16908 2295
rect 16856 2252 16908 2261
rect 21824 2329 21833 2363
rect 21833 2329 21867 2363
rect 21867 2329 21876 2363
rect 21824 2320 21876 2329
rect 22836 2320 22888 2372
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 1676 2048 1728 2100
rect 6092 2048 6144 2100
rect 9404 2048 9456 2100
rect 2228 1980 2280 2032
rect 6828 1980 6880 2032
rect 15844 76 15896 128
rect 16488 76 16540 128
rect 13912 8 13964 60
rect 19524 8 19576 60
<< metal2 >>
rect 20 27532 72 27538
rect 662 27532 718 28000
rect 662 27520 664 27532
rect 20 27474 72 27480
rect 716 27520 718 27532
rect 2042 27520 2098 28000
rect 2780 27532 2832 27538
rect 664 27474 716 27480
rect 32 6458 60 27474
rect 676 27443 704 27474
rect 1214 24848 1270 24857
rect 1214 24783 1270 24792
rect 1228 23662 1256 24783
rect 1216 23656 1268 23662
rect 110 23624 166 23633
rect 1216 23598 1268 23604
rect 110 23559 166 23568
rect 124 23322 152 23559
rect 112 23316 164 23322
rect 112 23258 164 23264
rect 1400 23180 1452 23186
rect 1400 23122 1452 23128
rect 1412 22574 1440 23122
rect 1400 22568 1452 22574
rect 1400 22510 1452 22516
rect 110 21856 166 21865
rect 110 21791 166 21800
rect 124 19281 152 21791
rect 110 19272 166 19281
rect 110 19207 166 19216
rect 1582 16008 1638 16017
rect 1582 15943 1638 15952
rect 1596 15706 1624 15943
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1412 14822 1440 15506
rect 2056 15434 2084 27520
rect 3422 27532 3478 28000
rect 3422 27520 3424 27532
rect 2780 27474 2832 27480
rect 3476 27520 3478 27532
rect 4356 27526 4752 27554
rect 3424 27474 3476 27480
rect 1492 15428 1544 15434
rect 1492 15370 1544 15376
rect 2044 15428 2096 15434
rect 2044 15370 2096 15376
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 110 13152 166 13161
rect 110 13087 166 13096
rect 124 12986 152 13087
rect 112 12980 164 12986
rect 112 12922 164 12928
rect 1504 11694 1532 15370
rect 1582 14376 1638 14385
rect 1582 14311 1638 14320
rect 1596 14074 1624 14311
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1504 9382 1532 10066
rect 1964 9761 1992 13806
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 2056 11257 2084 12582
rect 2042 11248 2098 11257
rect 2042 11183 2098 11192
rect 2792 10810 2820 27474
rect 3436 27443 3464 27474
rect 4068 23520 4120 23526
rect 4356 23474 4384 27526
rect 4724 27520 4752 27526
rect 4802 27520 4858 28000
rect 6182 27520 6238 28000
rect 7654 27520 7710 28000
rect 9034 27520 9090 28000
rect 10414 27520 10470 28000
rect 10520 27526 10824 27554
rect 10520 27520 10548 27526
rect 4724 27492 4844 27520
rect 4710 26616 4766 26625
rect 4710 26551 4766 26560
rect 4724 23662 4752 26551
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6196 23866 6224 27520
rect 6184 23860 6236 23866
rect 6184 23802 6236 23808
rect 4712 23656 4764 23662
rect 4712 23598 4764 23604
rect 4068 23462 4120 23468
rect 3422 17776 3478 17785
rect 3422 17711 3478 17720
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 1950 9752 2006 9761
rect 1950 9687 2006 9696
rect 3436 9625 3464 17711
rect 3974 10840 4030 10849
rect 3974 10775 4030 10784
rect 3988 10130 4016 10775
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 3988 9722 4016 10066
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 3422 9616 3478 9625
rect 4080 9586 4108 23462
rect 4264 23446 4384 23474
rect 4158 9752 4214 9761
rect 4158 9687 4214 9696
rect 3422 9551 3478 9560
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1398 9072 1454 9081
rect 1398 9007 1454 9016
rect 848 8560 900 8566
rect 848 8502 900 8508
rect 20 6452 72 6458
rect 20 6394 72 6400
rect 478 82 534 480
rect 860 82 888 8502
rect 1412 7857 1440 9007
rect 1398 7848 1454 7857
rect 1398 7783 1454 7792
rect 1412 7342 1440 7783
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1504 6633 1532 9318
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 1596 7478 1624 7511
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1490 6624 1546 6633
rect 1490 6559 1546 6568
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 1676 2100 1728 2106
rect 1676 2042 1728 2048
rect 478 54 888 82
rect 1398 82 1454 480
rect 1688 82 1716 2042
rect 2228 2032 2280 2038
rect 2228 1974 2280 1980
rect 1398 54 1716 82
rect 2240 82 2268 1974
rect 2318 82 2374 480
rect 2240 54 2374 82
rect 478 0 534 54
rect 1398 0 1454 54
rect 2318 0 2374 54
rect 3330 82 3386 480
rect 3528 82 3556 3946
rect 3330 54 3556 82
rect 4172 82 4200 9687
rect 4264 9518 4292 23446
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 7472 17808 7524 17814
rect 7472 17750 7524 17756
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 7484 17338 7512 17750
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5276 13841 5304 14758
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5262 13832 5318 13841
rect 5262 13767 5318 13776
rect 5170 10704 5226 10713
rect 5170 10639 5226 10648
rect 5184 9761 5212 10639
rect 5170 9752 5226 9761
rect 5170 9687 5226 9696
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4540 8498 4568 8910
rect 5276 8786 5304 13767
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5368 9722 5396 9998
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5356 9444 5408 9450
rect 5460 9432 5488 10134
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5408 9404 5488 9432
rect 5356 9386 5408 9392
rect 5368 8906 5396 9386
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5276 8758 5396 8786
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5276 8090 5304 8434
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5276 5642 5304 6190
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5368 4154 5396 8758
rect 5552 7818 5580 8910
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6012 8498 6040 9998
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6012 7886 6040 8434
rect 6104 7954 6132 17070
rect 7208 16726 7236 17138
rect 7668 17134 7696 27520
rect 9048 24857 9076 27520
rect 10428 27492 10548 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 9034 24848 9090 24857
rect 9034 24783 9090 24792
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10796 24274 10824 27526
rect 11440 27526 11744 27554
rect 10784 24268 10836 24274
rect 10784 24210 10836 24216
rect 8024 23724 8076 23730
rect 8024 23666 8076 23672
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7760 18426 7788 23462
rect 7748 18420 7800 18426
rect 7748 18362 7800 18368
rect 8036 18290 8064 23666
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 8574 19816 8630 19825
rect 8574 19751 8630 19760
rect 8588 19242 8616 19751
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11348 19281 11376 19314
rect 11334 19272 11390 19281
rect 8576 19236 8628 19242
rect 11334 19207 11390 19216
rect 8576 19178 8628 19184
rect 8588 18834 8616 19178
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10888 18970 10916 19110
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8588 18426 8616 18770
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8220 17814 8248 18022
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8116 17672 8168 17678
rect 8116 17614 8168 17620
rect 8128 17338 8156 17614
rect 8772 17610 8800 18158
rect 9048 17882 9076 18226
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 8760 17604 8812 17610
rect 8760 17546 8812 17552
rect 9508 17338 9536 18022
rect 8116 17332 8168 17338
rect 8116 17274 8168 17280
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 8128 16794 8156 17274
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8680 16726 8708 17070
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 8668 16720 8720 16726
rect 8668 16662 8720 16668
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 6748 15978 6776 16594
rect 8128 16250 8156 16594
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 8128 15026 8156 16186
rect 8404 16046 8432 16594
rect 9600 16114 9628 18090
rect 9876 18086 9904 18838
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 10060 17678 10088 18634
rect 10244 18426 10272 18702
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10888 18290 10916 18906
rect 11348 18834 11376 19207
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10692 17808 10744 17814
rect 10692 17750 10744 17756
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 16250 9720 16526
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8312 15434 8340 15982
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8404 15366 8432 15982
rect 8944 15972 8996 15978
rect 8944 15914 8996 15920
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8404 14482 8432 15302
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 7944 13462 7972 13806
rect 7932 13456 7984 13462
rect 8128 13433 8156 13806
rect 8220 13734 8248 14418
rect 8392 13796 8444 13802
rect 8392 13738 8444 13744
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 7932 13398 7984 13404
rect 8114 13424 8170 13433
rect 8024 13388 8076 13394
rect 8114 13359 8116 13368
rect 8024 13330 8076 13336
rect 8168 13359 8170 13368
rect 8116 13330 8168 13336
rect 8036 12918 8064 13330
rect 8128 12986 8156 13330
rect 8220 13297 8248 13670
rect 8206 13288 8262 13297
rect 8206 13223 8262 13232
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8024 12912 8076 12918
rect 8404 12889 8432 13738
rect 8024 12854 8076 12860
rect 8390 12880 8446 12889
rect 8390 12815 8446 12824
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7300 10538 7328 10950
rect 7484 10606 7512 10950
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7288 10532 7340 10538
rect 7288 10474 7340 10480
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6276 9444 6328 9450
rect 6276 9386 6328 9392
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6196 8294 6224 9046
rect 6288 8498 6316 9386
rect 7116 9382 7144 9862
rect 7576 9722 7604 11494
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7760 10266 7788 11086
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7760 10130 7788 10202
rect 7944 10130 7972 11698
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5538 7304 5594 7313
rect 5538 7239 5594 7248
rect 5552 6866 5580 7239
rect 6012 7002 6040 7822
rect 6104 7546 6132 7890
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 6092 6860 6144 6866
rect 6196 6848 6224 8230
rect 6288 8022 6316 8434
rect 6932 8362 6960 8774
rect 7116 8566 7144 9318
rect 7760 9178 7788 10066
rect 7944 9722 7972 10066
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6932 8090 6960 8298
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6144 6820 6224 6848
rect 6092 6802 6144 6808
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5460 6254 5488 6598
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5460 5098 5488 6190
rect 5552 5914 5580 6802
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5368 4126 5580 4154
rect 5552 2514 5580 4126
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 4250 82 4306 480
rect 4172 54 4306 82
rect 3330 0 3386 54
rect 4250 0 4306 54
rect 5262 82 5318 480
rect 5552 82 5580 2450
rect 5906 2408 5962 2417
rect 5816 2372 5868 2378
rect 5868 2352 5906 2360
rect 5868 2343 5962 2352
rect 5868 2332 5948 2343
rect 5816 2314 5868 2320
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5262 54 5580 82
rect 6012 82 6040 6598
rect 6104 6118 6132 6802
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6104 2106 6132 6054
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 6196 5370 6224 5578
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6288 3602 6316 7482
rect 6656 7410 6684 7958
rect 7024 7410 7052 8434
rect 7300 8362 7328 8910
rect 7484 8906 7512 8978
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7484 8090 7512 8842
rect 8036 8634 8064 10610
rect 8220 10538 8248 11562
rect 8588 10792 8616 14758
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8772 13161 8800 13262
rect 8758 13152 8814 13161
rect 8758 13087 8814 13096
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8852 12164 8904 12170
rect 8852 12106 8904 12112
rect 8772 11665 8800 12106
rect 8864 11694 8892 12106
rect 8852 11688 8904 11694
rect 8758 11656 8814 11665
rect 8852 11630 8904 11636
rect 8758 11591 8814 11600
rect 8772 11558 8800 11591
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8588 10764 8708 10792
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8496 10470 8524 10678
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8036 8362 8064 8570
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7208 7410 7236 7822
rect 8220 7750 8248 9522
rect 8496 9382 8524 10406
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8588 8838 8616 10610
rect 8680 8945 8708 10764
rect 8666 8936 8722 8945
rect 8666 8871 8722 8880
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8430 8616 8774
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6380 5914 6408 6734
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6564 5778 6592 6258
rect 6840 6254 6868 6598
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 6932 6100 6960 6190
rect 6840 6072 6960 6100
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6564 5030 6592 5714
rect 6748 5370 6776 5714
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6564 4010 6592 4626
rect 6840 4185 6868 6072
rect 7116 5846 7144 6190
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 6826 4176 6882 4185
rect 6826 4111 6882 4120
rect 6920 4140 6972 4146
rect 6840 4010 6868 4111
rect 6920 4082 6972 4088
rect 6932 4049 6960 4082
rect 6918 4040 6974 4049
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6828 4004 6880 4010
rect 6918 3975 6974 3984
rect 6828 3946 6880 3952
rect 6564 3641 6592 3946
rect 6550 3632 6606 3641
rect 6276 3596 6328 3602
rect 6550 3567 6606 3576
rect 6276 3538 6328 3544
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6196 2961 6224 2994
rect 6182 2952 6238 2961
rect 6182 2887 6238 2896
rect 6092 2100 6144 2106
rect 6092 2042 6144 2048
rect 6840 2038 6868 3946
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7024 3194 7052 3538
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7208 3126 7236 7346
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7576 7002 7604 7210
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 7300 5778 7328 6870
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7380 5636 7432 5642
rect 7432 5596 7512 5624
rect 7380 5578 7432 5584
rect 7484 4554 7512 5596
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7484 4214 7512 4490
rect 7576 4457 7604 6122
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7944 5778 7972 6054
rect 8220 5846 8248 7686
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8404 7002 8432 7142
rect 8496 7002 8524 8298
rect 8588 7954 8616 8366
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8588 7546 8616 7890
rect 8680 7818 8708 8230
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8772 7698 8800 11494
rect 8864 10062 8892 11630
rect 8956 11218 8984 15914
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9048 13734 9076 14418
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 12714 9076 13670
rect 9140 13530 9168 15030
rect 9324 14958 9352 15302
rect 9784 15162 9812 16186
rect 9876 15502 9904 17478
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 10060 16794 10088 17002
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16794 10732 17750
rect 10784 17604 10836 17610
rect 10784 17546 10836 17552
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10060 16250 10088 16730
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10796 16182 10824 17546
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9772 15156 9824 15162
rect 9692 15116 9772 15144
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9232 13938 9260 14214
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9232 13326 9260 13874
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9232 12918 9260 13126
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 9324 12646 9352 14894
rect 9692 14822 9720 15116
rect 9772 15098 9824 15104
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14550 9720 14758
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9692 14074 9720 14486
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9632 13828 9688 13837
rect 9784 13814 9812 14894
rect 9876 14618 9904 15438
rect 9968 15366 9996 15914
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10048 15632 10100 15638
rect 10048 15574 10100 15580
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9688 13786 9812 13814
rect 9632 13763 9688 13772
rect 9634 13728 9686 13734
rect 9600 13676 9634 13682
rect 9600 13670 9686 13676
rect 9600 13654 9674 13670
rect 9600 13530 9628 13654
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9494 13424 9550 13433
rect 9494 13359 9550 13368
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9312 12096 9364 12102
rect 9364 12056 9444 12084
rect 9312 12038 9364 12044
rect 9416 11694 9444 12056
rect 9508 11762 9536 13359
rect 9876 13258 9904 14554
rect 10060 14074 10088 15574
rect 10152 15162 10180 15846
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10508 15632 10560 15638
rect 10508 15574 10560 15580
rect 10520 15162 10548 15574
rect 10796 15570 10824 16118
rect 10980 15638 11008 18090
rect 11256 17814 11284 18702
rect 11244 17808 11296 17814
rect 11244 17750 11296 17756
rect 10968 15632 11020 15638
rect 10968 15574 11020 15580
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10980 15162 11008 15574
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10980 14618 11008 15098
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13530 10732 14350
rect 11440 14074 11468 27526
rect 11716 27520 11744 27526
rect 11794 27520 11850 28000
rect 13174 27520 13230 28000
rect 14646 27520 14702 28000
rect 16026 27520 16082 28000
rect 17406 27520 17462 28000
rect 18786 27520 18842 28000
rect 19524 27532 19576 27538
rect 11716 27492 11836 27520
rect 13188 23866 13216 27520
rect 14660 23866 14688 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15934 24848 15990 24857
rect 15934 24783 15990 24792
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 13176 23860 13228 23866
rect 13176 23802 13228 23808
rect 14648 23860 14700 23866
rect 14648 23802 14700 23808
rect 15948 23662 15976 24783
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 15936 23656 15988 23662
rect 15936 23598 15988 23604
rect 12452 22710 12480 23598
rect 14832 23520 14884 23526
rect 14832 23462 14884 23468
rect 11980 22704 12032 22710
rect 11980 22646 12032 22652
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 11992 22574 12020 22646
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11624 16726 11652 19654
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11716 16998 11744 17818
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11808 17338 11836 17750
rect 11900 17678 11928 18090
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11716 16726 11744 16934
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11624 16250 11652 16662
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11716 16114 11744 16662
rect 11900 16590 11928 17614
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11716 14618 11744 15438
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 10876 14000 10928 14006
rect 10876 13942 10928 13948
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 9140 11014 9168 11630
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 9048 10130 9076 10474
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8944 9988 8996 9994
rect 8944 9930 8996 9936
rect 8956 9654 8984 9930
rect 9048 9926 9076 10066
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 9048 9450 9076 9862
rect 9324 9518 9352 9862
rect 9416 9586 9444 11630
rect 9692 9722 9720 12718
rect 9968 12374 9996 13330
rect 10152 12714 10180 13330
rect 10782 13288 10838 13297
rect 10782 13223 10838 13232
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10060 11354 10088 12038
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10796 11354 10824 13223
rect 10888 12442 10916 13942
rect 11440 13870 11468 14010
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 10980 13530 11008 13670
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10980 12850 11008 13466
rect 11348 13462 11376 13738
rect 11532 13462 11560 14554
rect 11336 13456 11388 13462
rect 11336 13398 11388 13404
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11348 12918 11376 13398
rect 11808 12986 11836 13398
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 11992 12753 12020 22510
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 12084 19174 12112 19858
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13924 19378 13952 19654
rect 14844 19514 14872 23462
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 13544 19236 13596 19242
rect 13544 19178 13596 19184
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12084 18970 12112 19110
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12176 18426 12204 18770
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12820 18222 12848 18566
rect 12912 18222 12940 19110
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 12084 15570 12112 17614
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12636 16454 12664 17070
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12084 15366 12112 15506
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12176 14074 12204 14962
rect 12532 14952 12584 14958
rect 12452 14912 12532 14940
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12176 13870 12204 14010
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 11978 12744 12034 12753
rect 10968 12708 11020 12714
rect 11978 12679 12034 12688
rect 10968 12650 11020 12656
rect 10980 12442 11008 12650
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10888 11898 10916 12378
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9968 9926 9996 10950
rect 10336 10674 10364 11154
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10796 10538 10824 11290
rect 10888 11014 10916 11698
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10888 10674 10916 10950
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10784 10532 10836 10538
rect 10784 10474 10836 10480
rect 11164 10470 11192 11086
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 9048 9042 9076 9386
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9324 8974 9352 9454
rect 9600 9382 9628 9590
rect 9968 9586 9996 9862
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9508 8838 9536 8978
rect 9600 8838 9628 9318
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9508 8634 9536 8774
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8864 7750 8892 8366
rect 8680 7670 8800 7698
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8496 6118 8524 6734
rect 8588 6254 8616 7482
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 7944 5574 7972 5714
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7562 4448 7618 4457
rect 7562 4383 7618 4392
rect 7760 4214 7788 4966
rect 7944 4690 7972 5510
rect 8128 4826 8156 5646
rect 8312 5166 8340 5714
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8312 4690 8340 5102
rect 8404 5098 8432 5578
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7748 4208 7800 4214
rect 7748 4150 7800 4156
rect 7944 4146 7972 4626
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7944 3738 7972 4082
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7746 3496 7802 3505
rect 7746 3431 7802 3440
rect 8208 3460 8260 3466
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 6828 2032 6880 2038
rect 6828 1974 6880 1980
rect 6182 82 6238 480
rect 6012 54 6238 82
rect 5262 0 5318 54
rect 6182 0 6238 54
rect 7194 82 7250 480
rect 7300 82 7328 2246
rect 7484 1737 7512 2790
rect 7760 2650 7788 3431
rect 8208 3402 8260 3408
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 7944 2650 7972 2790
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 7470 1728 7526 1737
rect 7470 1663 7526 1672
rect 8036 1465 8064 3334
rect 8022 1456 8078 1465
rect 8022 1391 8078 1400
rect 7194 54 7328 82
rect 8114 82 8170 480
rect 8220 82 8248 3402
rect 8312 3398 8340 4626
rect 8680 4154 8708 7670
rect 8864 7274 8892 7686
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8772 6322 8800 7142
rect 8864 6662 8892 7210
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8864 6322 8892 6598
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8942 5808 8998 5817
rect 8942 5743 8998 5752
rect 8588 4126 8708 4154
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 8496 2650 8524 2858
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8588 2378 8616 4126
rect 8956 3602 8984 5743
rect 9048 5370 9076 8502
rect 9968 8498 9996 9522
rect 10060 9382 10088 9998
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10612 9654 10640 9862
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10704 9518 10732 10066
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 9586 11100 9862
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 8974 10088 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 10060 8022 10088 8910
rect 10152 8090 10180 8978
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10704 7954 10732 9454
rect 10980 9382 11008 9454
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 11072 9178 11100 9522
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8294 10824 8774
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9232 6254 9260 6938
rect 10152 6730 10180 7890
rect 10600 7812 10652 7818
rect 10796 7800 10824 8230
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10652 7772 10824 7800
rect 10600 7754 10652 7760
rect 10612 7274 10640 7754
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10692 7200 10744 7206
rect 10888 7188 10916 7890
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10744 7160 10916 7188
rect 10692 7142 10744 7148
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9220 6248 9272 6254
rect 9272 6208 9444 6236
rect 9220 6190 9272 6196
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9048 5166 9076 5306
rect 9232 5302 9260 5646
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 9048 4214 9076 5102
rect 9324 4486 9352 5782
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 8114 54 8248 82
rect 8864 82 8892 3334
rect 8956 3194 8984 3538
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9140 3058 9168 3946
rect 9324 3602 9352 4422
rect 9416 3670 9444 6208
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9600 5778 9628 6054
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9600 4622 9628 5714
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9784 5166 9812 5578
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9600 4146 9628 4558
rect 9692 4486 9720 4626
rect 9784 4554 9812 5102
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9600 4017 9628 4082
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9508 3602 9536 4014
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9324 3398 9352 3538
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9140 2514 9168 2994
rect 9324 2990 9352 3334
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9692 2582 9720 4082
rect 9968 4060 9996 6258
rect 10704 6225 10732 7142
rect 10980 7002 11008 7278
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11164 6390 11192 10406
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 7886 11284 8230
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11256 7342 11284 7822
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11348 6866 11376 10474
rect 11440 9586 11468 12106
rect 11900 11898 11928 12310
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11532 11286 11560 11834
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11532 10810 11560 11222
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11900 10470 11928 11086
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11900 10198 11928 10406
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 12084 9178 12112 9998
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 11624 9042 11652 9114
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11624 8634 11652 8978
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11152 6384 11204 6390
rect 11152 6326 11204 6332
rect 10784 6248 10836 6254
rect 10690 6216 10746 6225
rect 10784 6190 10836 6196
rect 10690 6151 10746 6160
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10796 5778 10824 6190
rect 11348 5778 11376 6802
rect 11532 6322 11560 7210
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 10784 5772 10836 5778
rect 11336 5772 11388 5778
rect 10784 5714 10836 5720
rect 11256 5732 11336 5760
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 11256 4826 11284 5732
rect 11336 5714 11388 5720
rect 11532 5234 11560 6122
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10152 4185 10180 4626
rect 10428 4593 10456 4694
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10414 4584 10470 4593
rect 10414 4519 10470 4528
rect 10138 4176 10194 4185
rect 10138 4111 10194 4120
rect 10520 4078 10548 4626
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 10140 4072 10192 4078
rect 9968 4032 10140 4060
rect 10140 4014 10192 4020
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9876 3738 9904 3878
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9876 3194 9904 3674
rect 10152 3602 10180 4014
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10600 3596 10652 3602
rect 10704 3584 10732 3878
rect 10888 3738 10916 4014
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10652 3556 10732 3584
rect 10600 3538 10652 3544
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 9048 2310 9076 2450
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9416 2106 9444 2450
rect 10060 2378 10088 3470
rect 10612 3058 10640 3538
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10888 2990 10916 3674
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11164 3058 11192 3470
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11256 2990 11284 4558
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10796 2514 10824 2858
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 9772 2372 9824 2378
rect 9772 2314 9824 2320
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 9404 2100 9456 2106
rect 9404 2042 9456 2048
rect 9126 82 9182 480
rect 8864 54 9182 82
rect 9784 82 9812 2314
rect 10046 82 10102 480
rect 9784 54 10102 82
rect 10704 82 10732 2382
rect 11348 649 11376 5102
rect 11624 5098 11652 8570
rect 11808 8294 11836 8978
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12084 8498 12112 8910
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 12084 8022 12112 8230
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 11704 7200 11756 7206
rect 12084 7188 12112 7958
rect 12176 7410 12204 13806
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12164 7200 12216 7206
rect 12084 7160 12164 7188
rect 11704 7142 11756 7148
rect 12164 7142 12216 7148
rect 11716 6866 11744 7142
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 11716 6254 11744 6802
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11900 5778 11928 6734
rect 12084 6118 12112 6802
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12084 5846 12112 6054
rect 12072 5840 12124 5846
rect 12176 5828 12204 7142
rect 12268 6769 12296 14554
rect 12452 14278 12480 14912
rect 12532 14894 12584 14900
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12452 13433 12480 14214
rect 12438 13424 12494 13433
rect 12438 13359 12494 13368
rect 12636 13297 12664 16390
rect 12820 15434 12848 18158
rect 12912 17542 12940 18158
rect 13360 18148 13412 18154
rect 13360 18090 13412 18096
rect 13372 17882 13400 18090
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13358 17776 13414 17785
rect 13358 17711 13414 17720
rect 13372 17678 13400 17711
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12912 17134 12940 17478
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12820 13394 12848 15370
rect 12912 14958 12940 17070
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 13188 16114 13216 17002
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 16726 13492 16934
rect 13556 16726 13584 19178
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13740 18358 13768 18838
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13740 18086 13768 18294
rect 14568 18290 14596 18702
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13188 15706 13216 16050
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 13004 14890 13032 15438
rect 12992 14884 13044 14890
rect 12992 14826 13044 14832
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13004 14618 13032 14826
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 13188 14414 13216 14826
rect 13464 14618 13492 15914
rect 13556 15706 13584 16662
rect 13740 15910 13768 18022
rect 14096 17876 14148 17882
rect 14096 17818 14148 17824
rect 14108 17202 14136 17818
rect 14292 17542 14320 18090
rect 14568 17678 14596 18226
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 13832 16250 13860 16662
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13740 15638 13768 15846
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13740 15162 13768 15574
rect 13832 15162 13860 16186
rect 13924 15978 13952 16934
rect 14568 16794 14596 17614
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14844 16590 14872 19178
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15580 18358 15608 18838
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15672 18358 15700 18702
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 15660 18352 15712 18358
rect 15660 18294 15712 18300
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15396 17338 15424 18022
rect 15476 17808 15528 17814
rect 15476 17750 15528 17756
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15396 16998 15424 17274
rect 15488 17270 15516 17750
rect 15856 17678 15884 19246
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15580 17338 15608 17478
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15476 17264 15528 17270
rect 15476 17206 15528 17212
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15292 16720 15344 16726
rect 15292 16662 15344 16668
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14844 16250 14872 16526
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 15304 15978 15332 16662
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15488 15162 15516 15574
rect 15580 15502 15608 17138
rect 15856 16114 15884 17614
rect 15948 17610 15976 18226
rect 15936 17604 15988 17610
rect 15936 17546 15988 17552
rect 15936 17060 15988 17066
rect 15936 17002 15988 17008
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15856 15502 15884 16050
rect 15948 15706 15976 17002
rect 16040 16250 16068 27520
rect 17420 23866 17448 27520
rect 18800 24410 18828 27520
rect 20166 27520 20222 28000
rect 21638 27532 21694 28000
rect 21638 27520 21640 27532
rect 19524 27474 19576 27480
rect 18788 24404 18840 24410
rect 18788 24346 18840 24352
rect 17592 24268 17644 24274
rect 17592 24210 17644 24216
rect 17604 23866 17632 24210
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 16948 23656 17000 23662
rect 16948 23598 17000 23604
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16132 18290 16160 18702
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 16132 16182 16160 18226
rect 16776 17134 16804 18906
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 16794 16252 16934
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16120 16176 16172 16182
rect 16172 16136 16252 16164
rect 16120 16118 16172 16124
rect 16028 15972 16080 15978
rect 16028 15914 16080 15920
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15580 15162 15608 15438
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 13832 14822 13860 15098
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13832 14618 13860 14758
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 13084 13932 13136 13938
rect 12912 13892 13084 13920
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12622 13288 12678 13297
rect 12622 13223 12678 13232
rect 12820 12986 12848 13330
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12636 12238 12664 12650
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12360 11354 12388 12174
rect 12728 11694 12756 12854
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12452 11132 12480 11222
rect 12360 11104 12480 11132
rect 12360 9602 12388 11104
rect 12544 10606 12572 11562
rect 12728 11286 12756 11630
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12544 10130 12572 10542
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12532 10124 12584 10130
rect 12452 10084 12532 10112
rect 12452 9722 12480 10084
rect 12532 10066 12584 10072
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12360 9574 12480 9602
rect 12544 9586 12572 9930
rect 12636 9722 12664 10474
rect 12912 10266 12940 13892
rect 13084 13874 13136 13880
rect 13084 13796 13136 13802
rect 13084 13738 13136 13744
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 13004 11694 13032 12922
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 13096 11150 13124 13738
rect 13188 13530 13216 14350
rect 13464 14074 13492 14554
rect 14200 14278 14228 14826
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13464 13814 13492 14010
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13464 13786 13584 13814
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13452 12708 13504 12714
rect 13372 12668 13452 12696
rect 13372 12102 13400 12668
rect 13452 12650 13504 12656
rect 13556 12442 13584 13786
rect 13648 13394 13676 13942
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13648 12986 13676 13330
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13096 10266 13124 11086
rect 13372 11014 13400 12038
rect 13556 11626 13584 12378
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13556 11286 13584 11562
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13556 10810 13584 11222
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13556 10538 13584 10746
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12360 7206 12388 7822
rect 12452 7750 12480 9574
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 12820 8838 12848 9386
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 9110 12940 9318
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12820 8634 12848 8774
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 13096 8430 13124 8910
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 13188 8090 13216 9046
rect 13372 8974 13400 9386
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13464 8786 13492 10406
rect 13648 10130 13676 12310
rect 13740 11898 13768 13262
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 12306 13952 12582
rect 14200 12442 14228 14214
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 14292 13258 14320 13806
rect 15396 13326 15424 14350
rect 15488 14074 15516 15098
rect 16040 15026 16068 15914
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 15764 14890 15976 14906
rect 15752 14884 15976 14890
rect 15804 14878 15976 14884
rect 15752 14826 15804 14832
rect 15948 14822 15976 14878
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 16132 14618 16160 15846
rect 16224 15638 16252 16136
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16224 15026 16252 15574
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15672 13802 15700 14554
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 15660 13796 15712 13802
rect 15660 13738 15712 13744
rect 16040 13394 16068 14010
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16028 13388 16080 13394
rect 15948 13348 16028 13376
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14292 13161 14320 13194
rect 14278 13152 14334 13161
rect 14278 13087 14334 13096
rect 14660 12646 14688 13194
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15396 12889 15424 13262
rect 15948 12986 15976 13348
rect 16028 13330 16080 13336
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 16028 12912 16080 12918
rect 15382 12880 15438 12889
rect 14924 12844 14976 12850
rect 16592 12889 16620 13330
rect 16684 12968 16712 13806
rect 16684 12940 16804 12968
rect 16028 12854 16080 12860
rect 16578 12880 16634 12889
rect 15382 12815 15438 12824
rect 14924 12786 14976 12792
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13740 11218 13768 11630
rect 13832 11558 13860 12174
rect 14844 11898 14872 12582
rect 14936 12442 14964 12786
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 16040 12374 16068 12854
rect 16578 12815 16634 12824
rect 16672 12844 16724 12850
rect 16592 12782 16620 12815
rect 16672 12786 16724 12792
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16592 12374 16620 12718
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 16028 12368 16080 12374
rect 16028 12310 16080 12316
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13740 9382 13768 10066
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13542 8800 13598 8809
rect 13464 8758 13542 8786
rect 13542 8735 13598 8744
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12452 7342 12480 7686
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12254 6760 12310 6769
rect 12254 6695 12310 6704
rect 12452 5914 12480 7278
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 13188 5846 13216 6054
rect 13280 5914 13308 6258
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 12256 5840 12308 5846
rect 12176 5800 12256 5828
rect 12072 5782 12124 5788
rect 12256 5782 12308 5788
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11440 3942 11468 4626
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3602 11468 3878
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11440 3194 11468 3538
rect 11532 3398 11560 4422
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11428 2916 11480 2922
rect 11428 2858 11480 2864
rect 11440 2582 11468 2858
rect 11624 2582 11652 3334
rect 11808 2922 11836 4966
rect 11900 4826 11928 5714
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 12084 4622 12112 5510
rect 12820 4758 12848 5510
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13096 4826 13124 5170
rect 13188 5098 13216 5782
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12084 4282 12112 4558
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11978 4176 12034 4185
rect 11978 4111 12034 4120
rect 11992 3641 12020 4111
rect 11978 3632 12034 3641
rect 11978 3567 11980 3576
rect 12032 3567 12034 3576
rect 11980 3538 12032 3544
rect 11992 3194 12020 3538
rect 12268 3534 12296 4694
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12820 4146 12848 4558
rect 13464 4282 13492 4694
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13556 4154 13584 8735
rect 13648 6361 13676 9114
rect 13740 7546 13768 9318
rect 13832 9178 13860 11494
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10674 14320 10950
rect 14844 10810 14872 11494
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14292 10198 14320 10610
rect 15304 10266 15332 11154
rect 15396 11150 15424 12174
rect 15488 11558 15516 12310
rect 16040 11830 16068 12310
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 11354 16252 11494
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15384 10464 15436 10470
rect 15488 10452 15516 11222
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15764 10674 15792 10950
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15856 10538 15884 11018
rect 16040 10674 16068 11086
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 15436 10424 15516 10452
rect 15384 10406 15436 10412
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 14016 8945 14044 9454
rect 14002 8936 14058 8945
rect 13912 8900 13964 8906
rect 14108 8906 14136 9998
rect 14186 9480 14242 9489
rect 14186 9415 14242 9424
rect 14200 9382 14228 9415
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14384 9042 14412 9998
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15396 9110 15424 10406
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 15948 10033 15976 10066
rect 16212 10056 16264 10062
rect 15934 10024 15990 10033
rect 16212 9998 16264 10004
rect 15934 9959 15990 9968
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15580 9722 15608 9862
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15580 9450 15608 9658
rect 15948 9654 15976 9959
rect 15936 9648 15988 9654
rect 15936 9590 15988 9596
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 14002 8871 14058 8880
rect 14096 8900 14148 8906
rect 13912 8842 13964 8848
rect 14096 8842 14148 8848
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13634 6352 13690 6361
rect 13634 6287 13690 6296
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13832 5370 13860 5782
rect 13924 5710 13952 8842
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14108 7954 14136 8434
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14108 7857 14136 7890
rect 14094 7848 14150 7857
rect 14094 7783 14150 7792
rect 14108 7478 14136 7783
rect 14844 7750 14872 8366
rect 15488 8090 15516 8978
rect 15580 8634 15608 9386
rect 15764 9178 15792 9522
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15856 8294 15884 9046
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15856 8022 15884 8230
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14096 7472 14148 7478
rect 14096 7414 14148 7420
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14568 6730 14596 7278
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 14752 6322 14780 7686
rect 14844 7410 14872 7686
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 15856 7206 15884 7958
rect 16040 7750 16068 9522
rect 16224 7954 16252 9998
rect 16592 9450 16620 10066
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 16684 9330 16712 12786
rect 16776 12782 16804 12940
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16776 12442 16804 12718
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 16776 11257 16804 12106
rect 16762 11248 16818 11257
rect 16762 11183 16818 11192
rect 16868 9926 16896 14758
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16592 9302 16712 9330
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 16040 7410 16068 7686
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14752 5914 14780 6258
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 14292 5574 14320 5850
rect 15120 5846 15148 6122
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 15304 5778 15332 6734
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15396 6633 15424 6666
rect 15382 6624 15438 6633
rect 15382 6559 15438 6568
rect 15488 6474 15516 6666
rect 15396 6446 15516 6474
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 14292 4758 14320 5510
rect 14280 4752 14332 4758
rect 14280 4694 14332 4700
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 13464 4126 13584 4154
rect 13912 4140 13964 4146
rect 12348 4004 12400 4010
rect 12544 3992 12572 4082
rect 12624 4004 12676 4010
rect 12544 3964 12624 3992
rect 12348 3946 12400 3952
rect 12624 3946 12676 3952
rect 12360 3602 12388 3946
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 3738 12480 3878
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12256 3528 12308 3534
rect 12452 3505 12480 3674
rect 12256 3470 12308 3476
rect 12438 3496 12494 3505
rect 12438 3431 12494 3440
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12636 2922 12664 3334
rect 11796 2916 11848 2922
rect 11796 2858 11848 2864
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 11428 2576 11480 2582
rect 11428 2518 11480 2524
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 11334 640 11390 649
rect 11334 575 11390 584
rect 11058 82 11114 480
rect 10704 54 11114 82
rect 7194 0 7250 54
rect 8114 0 8170 54
rect 9126 0 9182 54
rect 10046 0 10102 54
rect 11058 0 11114 54
rect 11978 96 12034 480
rect 12728 82 12756 3402
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 12912 2310 12940 3334
rect 13280 2990 13308 3334
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 13464 2009 13492 4126
rect 13912 4082 13964 4088
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13740 2922 13768 3606
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13924 2446 13952 4082
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14200 2650 14228 3538
rect 14384 2990 14412 3946
rect 14476 3097 14504 5646
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14924 5092 14976 5098
rect 14924 5034 14976 5040
rect 14738 4720 14794 4729
rect 14936 4690 14964 5034
rect 15304 4826 15332 5714
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 14738 4655 14794 4664
rect 14924 4684 14976 4690
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14568 4146 14596 4422
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14660 3398 14688 4558
rect 14752 4457 14780 4655
rect 14924 4626 14976 4632
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 14936 4593 14964 4626
rect 14922 4584 14978 4593
rect 14922 4519 14978 4528
rect 14738 4448 14794 4457
rect 14738 4383 14794 4392
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15304 3398 15332 4626
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 14462 3088 14518 3097
rect 14462 3023 14518 3032
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14292 2650 14320 2926
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 13912 2440 13964 2446
rect 14660 2417 14688 3334
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15212 2650 15240 3062
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15304 2553 15332 3334
rect 15290 2544 15346 2553
rect 15290 2479 15346 2488
rect 13912 2382 13964 2388
rect 14646 2408 14702 2417
rect 14646 2343 14702 2352
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 13450 2000 13506 2009
rect 13450 1935 13506 1944
rect 12990 82 13046 480
rect 12728 54 13046 82
rect 11978 0 12034 40
rect 12990 0 13046 54
rect 13910 60 13966 480
rect 13910 8 13912 60
rect 13964 8 13966 60
rect 13910 0 13966 8
rect 14922 82 14978 480
rect 15396 116 15424 6446
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15488 5574 15516 6258
rect 15856 5846 15884 7142
rect 16224 7002 16252 7890
rect 16316 7546 16344 8774
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16316 7274 16344 7482
rect 16408 7313 16436 8230
rect 16394 7304 16450 7313
rect 16304 7268 16356 7274
rect 16394 7239 16450 7248
rect 16304 7210 16356 7216
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16040 6458 16068 6802
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 15844 5840 15896 5846
rect 15844 5782 15896 5788
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 5302 15516 5510
rect 15856 5302 15884 5782
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 15856 4758 15884 5238
rect 15844 4752 15896 4758
rect 15844 4694 15896 4700
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15764 4010 15792 4218
rect 15856 4146 15884 4694
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15948 4010 15976 4422
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15752 4004 15804 4010
rect 15752 3946 15804 3952
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15474 3768 15530 3777
rect 15474 3703 15530 3712
rect 15488 3670 15516 3703
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15488 3194 15516 3606
rect 15672 3534 15700 3946
rect 15948 3652 15976 3946
rect 16028 3664 16080 3670
rect 15948 3624 16028 3652
rect 16028 3606 16080 3612
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15948 3194 15976 3402
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 16132 2378 16160 6054
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 16224 5370 16252 5510
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16500 4826 16528 5034
rect 16488 4820 16540 4826
rect 16316 4780 16488 4808
rect 16316 2961 16344 4780
rect 16488 4762 16540 4768
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16408 4078 16436 4218
rect 16592 4154 16620 9302
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16776 7478 16804 8366
rect 16960 7954 16988 23598
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 17052 15978 17080 16594
rect 17236 16046 17264 23598
rect 17604 17542 17632 23802
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17696 17746 17724 19314
rect 18616 17785 18644 20742
rect 19536 18222 19564 27474
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20180 23866 20208 27520
rect 21692 27520 21694 27532
rect 22468 27532 22520 27538
rect 21640 27474 21692 27480
rect 23018 27532 23074 28000
rect 24398 27554 24454 28000
rect 23018 27520 23020 27532
rect 22468 27474 22520 27480
rect 23072 27520 23074 27532
rect 24228 27526 24454 27554
rect 23020 27474 23072 27480
rect 21652 27443 21680 27474
rect 20168 23860 20220 23866
rect 20168 23802 20220 23808
rect 21456 23588 21508 23594
rect 21456 23530 21508 23536
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 21468 18358 21496 23530
rect 22008 22432 22060 22438
rect 22008 22374 22060 22380
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21560 18426 21588 18770
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 20536 18148 20588 18154
rect 20536 18090 20588 18096
rect 21456 18148 21508 18154
rect 21456 18090 21508 18096
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19444 17814 19472 18022
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 20548 17882 20576 18090
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 20536 17876 20588 17882
rect 20536 17818 20588 17824
rect 21100 17814 21128 18022
rect 19432 17808 19484 17814
rect 18602 17776 18658 17785
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17960 17740 18012 17746
rect 19432 17750 19484 17756
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 18602 17711 18658 17720
rect 17960 17682 18012 17688
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17420 16658 17448 17138
rect 17592 16992 17644 16998
rect 17696 16980 17724 17682
rect 17972 17202 18000 17682
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 17644 16952 17724 16980
rect 17592 16934 17644 16940
rect 17408 16652 17460 16658
rect 17408 16594 17460 16600
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17040 15972 17092 15978
rect 17040 15914 17092 15920
rect 17420 15910 17448 16594
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17420 14482 17448 15846
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17328 14074 17356 14418
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17328 13814 17356 14010
rect 17420 13870 17448 14418
rect 17500 14000 17552 14006
rect 17500 13942 17552 13948
rect 17236 13786 17356 13814
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17236 10033 17264 13786
rect 17420 13394 17448 13806
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17328 12442 17356 13330
rect 17420 12986 17448 13330
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17222 10024 17278 10033
rect 17222 9959 17278 9968
rect 17328 9761 17356 12378
rect 17512 11218 17540 13942
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17512 10810 17540 11154
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17500 10124 17552 10130
rect 17604 10112 17632 16934
rect 18432 16658 18460 17614
rect 18788 17060 18840 17066
rect 18788 17002 18840 17008
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 18064 16114 18092 16526
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18234 16008 18290 16017
rect 18234 15943 18290 15952
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17788 15638 17816 15846
rect 17776 15632 17828 15638
rect 17776 15574 17828 15580
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17696 11665 17724 14894
rect 17788 14822 17816 15574
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17972 15162 18000 15438
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17788 12628 17816 14758
rect 17972 14550 18000 15098
rect 17960 14544 18012 14550
rect 17960 14486 18012 14492
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 18064 13870 18092 14214
rect 18248 14074 18276 15943
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 12918 18092 13806
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 17868 12640 17920 12646
rect 17788 12600 17868 12628
rect 17868 12582 17920 12588
rect 17880 12374 17908 12582
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17682 11656 17738 11665
rect 17682 11591 17738 11600
rect 17880 11558 17908 12310
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17972 10470 18000 11154
rect 18064 10674 18092 11698
rect 18156 10674 18184 12650
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 18340 11626 18368 12174
rect 18328 11620 18380 11626
rect 18328 11562 18380 11568
rect 18524 11218 18552 13262
rect 18616 11694 18644 16050
rect 18708 15473 18736 16934
rect 18800 16454 18828 17002
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18694 15464 18750 15473
rect 18694 15399 18750 15408
rect 18800 15162 18828 16390
rect 18984 16250 19012 16934
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18892 13938 18920 14214
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18708 12782 18736 13126
rect 18892 12850 18920 13262
rect 18984 13138 19012 15982
rect 19260 15892 19288 16730
rect 19352 16250 19380 17614
rect 19444 17066 19472 17750
rect 20904 17264 20956 17270
rect 20904 17206 20956 17212
rect 20916 17066 20944 17206
rect 19432 17060 19484 17066
rect 19432 17002 19484 17008
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20904 17060 20956 17066
rect 20904 17002 20956 17008
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19628 16182 19656 16594
rect 19616 16176 19668 16182
rect 19616 16118 19668 16124
rect 19340 15904 19392 15910
rect 19260 15864 19340 15892
rect 19340 15846 19392 15852
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19168 15026 19196 15302
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19168 13814 19196 14962
rect 19352 14958 19380 15846
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19352 14618 19380 14894
rect 20168 14884 20220 14890
rect 20168 14826 20220 14832
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19076 13786 19196 13814
rect 19076 13462 19104 13786
rect 19352 13734 19380 14554
rect 20180 14074 20208 14826
rect 20272 14822 20300 15506
rect 20640 15502 20668 17002
rect 20812 16720 20864 16726
rect 20916 16708 20944 17002
rect 20996 16788 21048 16794
rect 21100 16776 21128 17750
rect 21468 17678 21496 18090
rect 21548 17808 21600 17814
rect 21548 17750 21600 17756
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21048 16748 21128 16776
rect 20996 16730 21048 16736
rect 21192 16726 21220 17614
rect 21468 17066 21496 17614
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 20864 16680 20944 16708
rect 21180 16720 21232 16726
rect 20812 16662 20864 16668
rect 21180 16662 21232 16668
rect 20824 16250 20852 16662
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 21192 16114 21220 16662
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 20996 15972 21048 15978
rect 20996 15914 21048 15920
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 19352 13462 19380 13670
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 20180 13530 20208 13670
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 19064 13456 19116 13462
rect 19064 13398 19116 13404
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 18984 13110 19104 13138
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 18144 10668 18196 10674
rect 18144 10610 18196 10616
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18156 10130 18184 10406
rect 18248 10266 18276 11086
rect 18708 10985 18736 12718
rect 18694 10976 18750 10985
rect 18694 10911 18750 10920
rect 19076 10713 19104 13110
rect 19352 12918 19380 13398
rect 20272 13002 20300 14758
rect 20364 14618 20392 14758
rect 20456 14618 20484 15302
rect 20824 14822 20852 15574
rect 21008 15162 21036 15914
rect 21192 15706 21220 16050
rect 21180 15700 21232 15706
rect 21232 15660 21312 15688
rect 21180 15642 21232 15648
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 21100 14550 21128 15370
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20824 13870 20852 14418
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20996 13524 21048 13530
rect 21100 13512 21128 14486
rect 21284 14414 21312 15660
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21376 15162 21404 15438
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21468 15026 21496 17002
rect 21560 16998 21588 17750
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21560 16794 21588 16934
rect 21548 16788 21600 16794
rect 21548 16730 21600 16736
rect 21560 15434 21588 16730
rect 21732 15972 21784 15978
rect 21732 15914 21784 15920
rect 21744 15502 21772 15914
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 21548 15428 21600 15434
rect 21548 15370 21600 15376
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21744 14890 21772 15438
rect 21732 14884 21784 14890
rect 21732 14826 21784 14832
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21048 13484 21128 13512
rect 20996 13466 21048 13472
rect 20812 13456 20864 13462
rect 20812 13398 20864 13404
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20180 12974 20300 13002
rect 20180 12918 20208 12974
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 19352 11830 19380 12854
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 20088 12442 20116 12718
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 20180 12374 20208 12582
rect 20168 12368 20220 12374
rect 20168 12310 20220 12316
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19628 11830 19656 12038
rect 19340 11824 19392 11830
rect 19340 11766 19392 11772
rect 19616 11824 19668 11830
rect 19616 11766 19668 11772
rect 19352 11694 19380 11766
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19352 11558 19380 11630
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19352 11354 19380 11494
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19996 11354 20024 12242
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19062 10704 19118 10713
rect 19062 10639 19118 10648
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 17552 10084 17632 10112
rect 18144 10124 18196 10130
rect 17500 10066 17552 10072
rect 18144 10066 18196 10072
rect 17314 9752 17370 9761
rect 17314 9687 17370 9696
rect 17040 9036 17092 9042
rect 17040 8978 17092 8984
rect 17052 8498 17080 8978
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16776 6934 16804 7142
rect 17144 6934 17172 7686
rect 17328 7342 17356 9687
rect 17512 9382 17540 10066
rect 18156 9450 18184 10066
rect 18248 9586 18276 10202
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17512 8537 17540 9318
rect 17498 8528 17554 8537
rect 17554 8486 17632 8514
rect 17498 8463 17554 8472
rect 17408 7812 17460 7818
rect 17408 7754 17460 7760
rect 17420 7410 17448 7754
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 16764 6928 16816 6934
rect 16764 6870 16816 6876
rect 17132 6928 17184 6934
rect 17132 6870 17184 6876
rect 17144 6458 17172 6870
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16684 4214 16712 5170
rect 16776 5098 16804 6122
rect 16764 5092 16816 5098
rect 16764 5034 16816 5040
rect 16500 4126 16620 4154
rect 16672 4208 16724 4214
rect 16672 4150 16724 4156
rect 16764 4140 16816 4146
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16302 2952 16358 2961
rect 16302 2887 16358 2896
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 15304 88 15424 116
rect 15842 128 15898 480
rect 16500 134 16528 4126
rect 16764 4082 16816 4088
rect 16578 3496 16634 3505
rect 16578 3431 16634 3440
rect 16592 3398 16620 3431
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16592 3058 16620 3334
rect 16776 3194 16804 4082
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16868 3126 16896 6190
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 17144 5030 17172 5782
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17236 5098 17264 5646
rect 17224 5092 17276 5098
rect 17224 5034 17276 5040
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17144 4758 17172 4966
rect 17132 4752 17184 4758
rect 17132 4694 17184 4700
rect 17328 4690 17356 6938
rect 17420 6866 17448 7346
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17512 6798 17540 7686
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17328 4282 17356 4626
rect 17040 4276 17092 4282
rect 17316 4276 17368 4282
rect 17092 4236 17172 4264
rect 17040 4218 17092 4224
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 15304 82 15332 88
rect 14922 54 15332 82
rect 15842 76 15844 128
rect 15896 76 15898 128
rect 14922 0 14978 54
rect 15842 0 15898 76
rect 16488 128 16540 134
rect 16488 70 16540 76
rect 16776 82 16804 2314
rect 16868 2310 16896 2450
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16868 1737 16896 2246
rect 17144 2009 17172 4236
rect 17316 4218 17368 4224
rect 17130 2000 17186 2009
rect 17130 1935 17186 1944
rect 16854 1728 16910 1737
rect 16854 1663 16910 1672
rect 16854 82 16910 480
rect 16776 54 16910 82
rect 17420 82 17448 6598
rect 17512 6458 17540 6734
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17604 6390 17632 8486
rect 17788 8362 17816 9318
rect 18156 8838 18184 9386
rect 18708 9382 18736 10406
rect 18786 9616 18842 9625
rect 18786 9551 18842 9560
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 17776 8356 17828 8362
rect 17776 8298 17828 8304
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17788 7206 17816 7890
rect 18156 7342 18184 8774
rect 18616 7750 18644 8910
rect 18708 8362 18736 9318
rect 18800 8430 18828 9551
rect 18788 8424 18840 8430
rect 18788 8366 18840 8372
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18800 8090 18828 8366
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18616 7410 18644 7686
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17592 6384 17644 6390
rect 17592 6326 17644 6332
rect 17788 5817 17816 7142
rect 18156 6866 18184 7278
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18800 6390 18828 6598
rect 18984 6458 19012 6734
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 17774 5808 17830 5817
rect 17774 5743 17830 5752
rect 18880 5636 18932 5642
rect 18880 5578 18932 5584
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18708 5302 18736 5510
rect 18696 5296 18748 5302
rect 18696 5238 18748 5244
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18708 5030 18736 5102
rect 18788 5092 18840 5098
rect 18788 5034 18840 5040
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17788 3641 17816 4422
rect 18524 4282 18552 4762
rect 18800 4758 18828 5034
rect 18892 4826 18920 5578
rect 18984 5545 19012 6394
rect 18970 5536 19026 5545
rect 18970 5471 19026 5480
rect 19076 5273 19104 10639
rect 19260 10266 19288 11154
rect 19352 10538 19380 11290
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 19996 10810 20024 10950
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19340 10532 19392 10538
rect 19340 10474 19392 10480
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19996 10266 20024 10610
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19168 9674 19196 10066
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19168 9646 19288 9674
rect 19062 5264 19118 5273
rect 19062 5199 19118 5208
rect 19156 5092 19208 5098
rect 19156 5034 19208 5040
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18788 4752 18840 4758
rect 18788 4694 18840 4700
rect 18878 4720 18934 4729
rect 19062 4720 19118 4729
rect 18934 4678 19012 4706
rect 18878 4655 18934 4664
rect 18984 4622 19012 4678
rect 19062 4655 19118 4664
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18880 4616 18932 4622
rect 18880 4558 18932 4564
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18420 4004 18472 4010
rect 18420 3946 18472 3952
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17972 3738 18000 3878
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17774 3632 17830 3641
rect 17774 3567 17830 3576
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17604 2650 17632 3470
rect 17788 2922 17816 3567
rect 17972 3194 18000 3674
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18432 3058 18460 3946
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18524 3194 18552 3334
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 18524 2854 18552 3130
rect 18512 2848 18564 2854
rect 18512 2790 18564 2796
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 17774 82 17830 480
rect 17420 54 17830 82
rect 18616 82 18644 4422
rect 18708 4146 18736 4558
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18708 4049 18736 4082
rect 18694 4040 18750 4049
rect 18694 3975 18750 3984
rect 18800 2650 18828 4218
rect 18892 4010 18920 4558
rect 19076 4146 19104 4655
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 19076 3738 19104 4082
rect 19168 4010 19196 5034
rect 19260 4282 19288 9646
rect 19444 9178 19472 9998
rect 20272 9994 20300 12786
rect 20364 12442 20392 12786
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20456 11694 20484 12650
rect 20640 12102 20668 13262
rect 20824 12782 20852 13398
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20640 11898 20668 12038
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20824 11694 20852 12718
rect 21100 12458 21128 12922
rect 20916 12430 21128 12458
rect 20916 11898 20944 12430
rect 21100 12374 21128 12430
rect 20996 12368 21048 12374
rect 20996 12310 21048 12316
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 21008 11898 21036 12310
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 21100 11150 21128 11698
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 20732 10266 20760 11086
rect 21192 10810 21220 11222
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 20904 10668 20956 10674
rect 21284 10656 21312 13806
rect 21376 11558 21404 14554
rect 21916 14476 21968 14482
rect 21916 14418 21968 14424
rect 21928 13802 21956 14418
rect 21916 13796 21968 13802
rect 21916 13738 21968 13744
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21744 12714 21772 13262
rect 21928 12889 21956 13738
rect 21914 12880 21970 12889
rect 21914 12815 21970 12824
rect 21732 12708 21784 12714
rect 21732 12650 21784 12656
rect 21744 12238 21772 12650
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21824 11280 21876 11286
rect 21824 11222 21876 11228
rect 21836 10742 21864 11222
rect 21824 10736 21876 10742
rect 21824 10678 21876 10684
rect 22020 10674 22048 22374
rect 22098 20360 22154 20369
rect 22098 20295 22154 20304
rect 22112 18834 22140 20295
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 22480 18426 22508 27474
rect 23032 27443 23060 27474
rect 23294 25256 23350 25265
rect 23294 25191 23350 25200
rect 23308 24274 23336 25191
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 22928 24064 22980 24070
rect 22928 24006 22980 24012
rect 22836 23588 22888 23594
rect 22756 23548 22836 23576
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22480 18222 22508 18362
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 22664 17814 22692 18566
rect 22652 17808 22704 17814
rect 22652 17750 22704 17756
rect 22376 17672 22428 17678
rect 22376 17614 22428 17620
rect 22388 16590 22416 17614
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22480 17134 22508 17478
rect 22664 17338 22692 17750
rect 22756 17610 22784 23548
rect 22836 23530 22888 23536
rect 22940 23474 22968 24006
rect 23308 23866 23336 24210
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 24228 23798 24256 27526
rect 24398 27520 24454 27526
rect 24860 27532 24912 27538
rect 25778 27532 25834 28000
rect 25778 27520 25780 27532
rect 24860 27474 24912 27480
rect 25832 27520 25834 27532
rect 26240 27532 26292 27538
rect 25780 27474 25832 27480
rect 27158 27532 27214 28000
rect 27158 27520 27160 27532
rect 26240 27474 26292 27480
rect 27212 27520 27214 27532
rect 27160 27474 27212 27480
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24216 23792 24268 23798
rect 24216 23734 24268 23740
rect 22848 23446 22968 23474
rect 22744 17604 22796 17610
rect 22744 17546 22796 17552
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 22468 17128 22520 17134
rect 22468 17070 22520 17076
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22572 16726 22600 16934
rect 22560 16720 22612 16726
rect 22560 16662 22612 16668
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22204 16250 22232 16526
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 22388 15162 22416 16526
rect 22572 15706 22600 16662
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22284 15088 22336 15094
rect 22284 15030 22336 15036
rect 22296 14550 22324 15030
rect 22284 14544 22336 14550
rect 22284 14486 22336 14492
rect 22296 14074 22324 14486
rect 22466 14376 22522 14385
rect 22466 14311 22522 14320
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 12850 22140 13670
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22388 12753 22416 12786
rect 22374 12744 22430 12753
rect 22284 12708 22336 12714
rect 22374 12679 22430 12688
rect 22284 12650 22336 12656
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 22100 11620 22152 11626
rect 22100 11562 22152 11568
rect 22112 11014 22140 11562
rect 22100 11008 22152 11014
rect 22100 10950 22152 10956
rect 22008 10668 22060 10674
rect 21284 10628 21496 10656
rect 20904 10610 20956 10616
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20260 9988 20312 9994
rect 20260 9930 20312 9936
rect 20824 9382 20852 9998
rect 20916 9586 20944 10610
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21284 10266 21312 10474
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 20996 10192 21048 10198
rect 20996 10134 21048 10140
rect 21008 9722 21036 10134
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 21008 9450 21036 9658
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 20996 9444 21048 9450
rect 20996 9386 21048 9392
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19352 8022 19380 8774
rect 19444 8498 19472 9114
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 20628 9104 20680 9110
rect 20628 9046 20680 9052
rect 19628 8838 19656 9046
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19628 8362 19656 8774
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19616 8356 19668 8362
rect 19616 8298 19668 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19996 8022 20024 8434
rect 20640 8294 20668 9046
rect 20824 8634 20852 9318
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 21008 8634 21036 8910
rect 21192 8906 21220 9522
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 21192 8362 21220 8842
rect 21284 8362 21312 9590
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 8022 20668 8230
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19984 8016 20036 8022
rect 19984 7958 20036 7964
rect 20628 8016 20680 8022
rect 20628 7958 20680 7964
rect 19352 7546 19380 7958
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19444 6934 19472 7142
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19996 6934 20024 7822
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 19432 6928 19484 6934
rect 19432 6870 19484 6876
rect 19984 6928 20036 6934
rect 19984 6870 20036 6876
rect 19444 6458 19472 6870
rect 20364 6662 20392 7346
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 20260 6180 20312 6186
rect 20260 6122 20312 6128
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19432 5840 19484 5846
rect 19432 5782 19484 5788
rect 19444 5030 19472 5782
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19536 4826 19564 5850
rect 20272 5642 20300 6122
rect 20260 5636 20312 5642
rect 20260 5578 20312 5584
rect 19892 5568 19944 5574
rect 19892 5510 19944 5516
rect 19904 5370 19932 5510
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 19524 4208 19576 4214
rect 19524 4150 19576 4156
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19156 4004 19208 4010
rect 19156 3946 19208 3952
rect 19260 3777 19288 4082
rect 19246 3768 19302 3777
rect 19064 3732 19116 3738
rect 19246 3703 19302 3712
rect 19064 3674 19116 3680
rect 19536 3670 19564 4150
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19524 3664 19576 3670
rect 19524 3606 19576 3612
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 18800 2446 18828 2586
rect 19260 2446 19288 2994
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 18786 82 18842 480
rect 18616 54 18842 82
rect 19536 66 19564 3334
rect 19996 3194 20024 3878
rect 20364 3466 20392 6598
rect 20444 6180 20496 6186
rect 20444 6122 20496 6128
rect 20456 5234 20484 6122
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20456 4826 20484 5170
rect 20548 5098 20576 5306
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20536 5092 20588 5098
rect 20536 5034 20588 5040
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20640 3942 20668 5170
rect 20732 4826 20760 5646
rect 20824 5574 20852 6734
rect 20916 6633 20944 6802
rect 21008 6730 21036 7822
rect 21192 7478 21220 8298
rect 21364 8016 21416 8022
rect 21364 7958 21416 7964
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 21284 7410 21312 7686
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 21376 7274 21404 7958
rect 21364 7268 21416 7274
rect 21364 7210 21416 7216
rect 21376 7002 21404 7210
rect 21364 6996 21416 7002
rect 21364 6938 21416 6944
rect 20996 6724 21048 6730
rect 20996 6666 21048 6672
rect 20902 6624 20958 6633
rect 20902 6559 20958 6568
rect 20916 6458 20944 6559
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 21364 6180 21416 6186
rect 21364 6122 21416 6128
rect 21088 5840 21140 5846
rect 21088 5782 21140 5788
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20824 4622 20852 5510
rect 21100 5030 21128 5782
rect 21376 5574 21404 6122
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21272 5092 21324 5098
rect 21272 5034 21324 5040
rect 21088 5024 21140 5030
rect 21088 4966 21140 4972
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20916 4282 20944 4626
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19996 2854 20024 3130
rect 20640 3126 20668 3878
rect 21008 3670 21036 4490
rect 21100 4154 21128 4966
rect 21100 4126 21220 4154
rect 21192 3670 21220 4126
rect 20996 3664 21048 3670
rect 20996 3606 21048 3612
rect 21180 3664 21232 3670
rect 21180 3606 21232 3612
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 21088 3120 21140 3126
rect 21088 3062 21140 3068
rect 20168 2916 20220 2922
rect 20168 2858 20220 2864
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20180 2650 20208 2858
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 20548 2582 20576 2790
rect 20536 2576 20588 2582
rect 20536 2518 20588 2524
rect 19984 2372 20036 2378
rect 19984 2314 20036 2320
rect 19706 82 19762 480
rect 19996 82 20024 2314
rect 16854 0 16910 54
rect 17774 0 17830 54
rect 18786 0 18842 54
rect 19524 60 19576 66
rect 19524 2 19576 8
rect 19706 54 20024 82
rect 20718 82 20774 480
rect 21100 82 21128 3062
rect 21192 2854 21220 3606
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21284 2582 21312 5034
rect 21376 3641 21404 5510
rect 21468 4690 21496 10628
rect 22008 10610 22060 10616
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21560 7410 21588 9930
rect 22112 9722 22140 10950
rect 22204 10810 22232 12582
rect 22296 11626 22324 12650
rect 22284 11620 22336 11626
rect 22284 11562 22336 11568
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22296 10470 22324 11086
rect 22388 10606 22416 12679
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22190 9752 22246 9761
rect 22100 9716 22152 9722
rect 22190 9687 22246 9696
rect 22100 9658 22152 9664
rect 22204 9654 22232 9687
rect 22192 9648 22244 9654
rect 22192 9590 22244 9596
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 22112 8945 22140 9454
rect 22098 8936 22154 8945
rect 22098 8871 22154 8880
rect 21914 8528 21970 8537
rect 21914 8463 21970 8472
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 21560 6934 21588 7346
rect 21548 6928 21600 6934
rect 21548 6870 21600 6876
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21652 5846 21680 6122
rect 21640 5840 21692 5846
rect 21640 5782 21692 5788
rect 21548 5636 21600 5642
rect 21548 5578 21600 5584
rect 21456 4684 21508 4690
rect 21456 4626 21508 4632
rect 21456 4140 21508 4146
rect 21456 4082 21508 4088
rect 21362 3632 21418 3641
rect 21362 3567 21418 3576
rect 21376 2582 21404 3567
rect 21468 3534 21496 4082
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21560 3194 21588 5578
rect 21928 5166 21956 8463
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 22112 6390 22140 6666
rect 22100 6384 22152 6390
rect 22100 6326 22152 6332
rect 22100 6180 22152 6186
rect 22100 6122 22152 6128
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 21732 5024 21784 5030
rect 21732 4966 21784 4972
rect 21744 4622 21772 4966
rect 21928 4826 21956 5102
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 21744 4282 21772 4558
rect 21732 4276 21784 4282
rect 21732 4218 21784 4224
rect 22112 4154 22140 6122
rect 22204 5778 22232 9590
rect 22192 5772 22244 5778
rect 22192 5714 22244 5720
rect 22204 4826 22232 5714
rect 22192 4820 22244 4826
rect 22192 4762 22244 4768
rect 22020 4126 22140 4154
rect 21732 3664 21784 3670
rect 21732 3606 21784 3612
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 21560 2854 21588 3130
rect 21744 3058 21772 3606
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 21836 3058 21864 3470
rect 21732 3052 21784 3058
rect 21732 2994 21784 3000
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 21836 2650 21864 2994
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 21272 2576 21324 2582
rect 21272 2518 21324 2524
rect 21364 2576 21416 2582
rect 21364 2518 21416 2524
rect 21454 2544 21510 2553
rect 21376 2446 21404 2518
rect 21454 2479 21510 2488
rect 21468 2446 21496 2479
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 21836 2378 21864 2586
rect 21824 2372 21876 2378
rect 21824 2314 21876 2320
rect 20718 54 21128 82
rect 21638 82 21694 480
rect 22020 82 22048 4126
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22204 3738 22232 3878
rect 22296 3738 22324 10406
rect 22376 8084 22428 8090
rect 22376 8026 22428 8032
rect 22388 6866 22416 8026
rect 22480 7954 22508 14311
rect 22848 13462 22876 23446
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24674 21992 24730 22001
rect 24674 21927 24730 21936
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21010 24716 21927
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20602 24716 20946
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24766 18864 24822 18873
rect 24766 18799 24822 18808
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24780 17882 24808 18799
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 23112 17808 23164 17814
rect 23112 17750 23164 17756
rect 23124 17270 23152 17750
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 23112 17264 23164 17270
rect 22926 17232 22982 17241
rect 23112 17206 23164 17212
rect 22926 17167 22982 17176
rect 22940 16250 22968 17167
rect 23848 17128 23900 17134
rect 23848 17070 23900 17076
rect 23204 16720 23256 16726
rect 23204 16662 23256 16668
rect 23216 16250 23244 16662
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 22940 16046 22968 16186
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 22940 14074 22968 15982
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 22928 14068 22980 14074
rect 22928 14010 22980 14016
rect 22940 13870 22968 14010
rect 22928 13864 22980 13870
rect 22928 13806 22980 13812
rect 23296 13796 23348 13802
rect 23296 13738 23348 13744
rect 22836 13456 22888 13462
rect 22836 13398 22888 13404
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22664 12374 22692 13126
rect 22940 12986 22968 13398
rect 22928 12980 22980 12986
rect 22980 12940 23060 12968
rect 22928 12922 22980 12928
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 22940 12374 22968 12582
rect 23032 12442 23060 12940
rect 23020 12436 23072 12442
rect 23020 12378 23072 12384
rect 22652 12368 22704 12374
rect 22652 12310 22704 12316
rect 22928 12368 22980 12374
rect 22928 12310 22980 12316
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 22572 11354 22600 12174
rect 22664 11898 22692 12310
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22848 11286 22876 12174
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23124 11626 23152 12038
rect 23112 11620 23164 11626
rect 23112 11562 23164 11568
rect 23124 11286 23152 11562
rect 22836 11280 22888 11286
rect 22836 11222 22888 11228
rect 23112 11280 23164 11286
rect 23112 11222 23164 11228
rect 23204 11280 23256 11286
rect 23204 11222 23256 11228
rect 23124 10810 23152 11222
rect 23112 10804 23164 10810
rect 23112 10746 23164 10752
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22480 7546 22508 7890
rect 22468 7540 22520 7546
rect 22468 7482 22520 7488
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22388 6458 22416 6802
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 22480 6254 22508 7482
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22664 6322 22692 6734
rect 22652 6316 22704 6322
rect 22652 6258 22704 6264
rect 22468 6248 22520 6254
rect 22468 6190 22520 6196
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22572 5710 22600 6054
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 22388 5030 22416 5102
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 22376 4480 22428 4486
rect 22376 4422 22428 4428
rect 22388 4049 22416 4422
rect 22572 4146 22600 4762
rect 22756 4154 22784 10542
rect 23216 10266 23244 11222
rect 23308 10470 23336 13738
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23676 13530 23704 13670
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23676 12918 23704 13466
rect 23664 12912 23716 12918
rect 23664 12854 23716 12860
rect 23572 11824 23624 11830
rect 23572 11766 23624 11772
rect 23480 11552 23532 11558
rect 23584 11540 23612 11766
rect 23532 11512 23612 11540
rect 23480 11494 23532 11500
rect 23768 11098 23796 14214
rect 23676 11070 23796 11098
rect 23296 10464 23348 10470
rect 23296 10406 23348 10412
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 23308 10198 23336 10406
rect 23296 10192 23348 10198
rect 23296 10134 23348 10140
rect 22928 10124 22980 10130
rect 22928 10066 22980 10072
rect 22940 9654 22968 10066
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 22928 9648 22980 9654
rect 22928 9590 22980 9596
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22940 5030 22968 5714
rect 22928 5024 22980 5030
rect 22928 4966 22980 4972
rect 22940 4690 22968 4966
rect 22836 4684 22888 4690
rect 22836 4626 22888 4632
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 22848 4282 22876 4626
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 22560 4140 22612 4146
rect 22756 4126 22876 4154
rect 22560 4082 22612 4088
rect 22848 4049 22876 4126
rect 22374 4040 22430 4049
rect 22374 3975 22430 3984
rect 22834 4040 22890 4049
rect 22834 3975 22890 3984
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22284 3732 22336 3738
rect 22284 3674 22336 3680
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 22480 3126 22508 3538
rect 23216 3194 23244 9862
rect 23308 9722 23336 10134
rect 23386 10024 23442 10033
rect 23386 9959 23442 9968
rect 23400 9926 23428 9959
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 23400 9602 23428 9862
rect 23308 9574 23428 9602
rect 23308 4758 23336 9574
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23400 5778 23428 8774
rect 23676 6934 23704 11070
rect 23754 10976 23810 10985
rect 23754 10911 23810 10920
rect 23768 10470 23796 10911
rect 23756 10464 23808 10470
rect 23756 10406 23808 10412
rect 23860 8430 23888 17070
rect 24228 16998 24256 17682
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24216 16992 24268 16998
rect 24216 16934 24268 16940
rect 24228 16017 24256 16934
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24214 16008 24270 16017
rect 24214 15943 24270 15952
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24032 14884 24084 14890
rect 24032 14826 24084 14832
rect 24044 14482 24072 14826
rect 24032 14476 24084 14482
rect 24032 14418 24084 14424
rect 24044 13802 24072 14418
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24872 14074 24900 27474
rect 25792 27443 25820 27474
rect 25134 26616 25190 26625
rect 25134 26551 25190 26560
rect 25148 23866 25176 26551
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25148 23662 25176 23802
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 25134 23488 25190 23497
rect 25134 23423 25190 23432
rect 25148 22778 25176 23423
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 25148 22574 25176 22714
rect 25136 22568 25188 22574
rect 25136 22510 25188 22516
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24032 13796 24084 13802
rect 24032 13738 24084 13744
rect 26252 13394 26280 27474
rect 27172 27443 27200 27474
rect 24768 13388 24820 13394
rect 24768 13330 24820 13336
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 24044 12850 24072 13262
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24780 12986 24808 13330
rect 27618 13152 27674 13161
rect 27618 13087 27674 13096
rect 27632 12986 27660 13087
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 27620 12980 27672 12986
rect 27620 12922 27672 12928
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 24044 11286 24072 12786
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 24216 12232 24268 12238
rect 24216 12174 24268 12180
rect 24136 11354 24164 12174
rect 24228 11830 24256 12174
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24780 11898 24808 12310
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24216 11824 24268 11830
rect 24216 11766 24268 11772
rect 24400 11824 24452 11830
rect 24400 11766 24452 11772
rect 24412 11354 24440 11766
rect 24124 11348 24176 11354
rect 24124 11290 24176 11296
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24032 11280 24084 11286
rect 24032 11222 24084 11228
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10810 24716 11154
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24136 10266 24164 10542
rect 24124 10260 24176 10266
rect 24124 10202 24176 10208
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24766 8800 24822 8809
rect 24289 8732 24585 8752
rect 24766 8735 24822 8744
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24780 8634 24808 8735
rect 24768 8628 24820 8634
rect 24768 8570 24820 8576
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 23664 6928 23716 6934
rect 23664 6870 23716 6876
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23388 5772 23440 5778
rect 23388 5714 23440 5720
rect 23400 5370 23428 5714
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23296 4752 23348 4758
rect 23296 4694 23348 4700
rect 23492 3505 23520 4966
rect 23478 3496 23534 3505
rect 23478 3431 23534 3440
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 22468 3120 22520 3126
rect 22374 3088 22430 3097
rect 22468 3062 22520 3068
rect 22374 3023 22430 3032
rect 22388 2990 22416 3023
rect 22376 2984 22428 2990
rect 22376 2926 22428 2932
rect 23572 2848 23624 2854
rect 23572 2790 23624 2796
rect 23584 2650 23612 2790
rect 23768 2650 23796 6598
rect 24044 6118 24072 6802
rect 24214 6760 24270 6769
rect 24214 6695 24270 6704
rect 24228 6322 24256 6695
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24872 6361 24900 12718
rect 25044 11212 25096 11218
rect 25044 11154 25096 11160
rect 25056 10470 25084 11154
rect 25410 11112 25466 11121
rect 25410 11047 25466 11056
rect 25424 10810 25452 11047
rect 25412 10804 25464 10810
rect 25412 10746 25464 10752
rect 25228 10600 25280 10606
rect 25228 10542 25280 10548
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 25056 8537 25084 10406
rect 25240 9518 25268 10542
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25042 8528 25098 8537
rect 25042 8463 25098 8472
rect 27620 6996 27672 7002
rect 27620 6938 27672 6944
rect 27632 6905 27660 6938
rect 27618 6896 27674 6905
rect 25504 6860 25556 6866
rect 27618 6831 27674 6840
rect 25504 6802 25556 6808
rect 25516 6458 25544 6802
rect 25504 6452 25556 6458
rect 25504 6394 25556 6400
rect 24858 6352 24914 6361
rect 24216 6316 24268 6322
rect 24858 6287 24914 6296
rect 24216 6258 24268 6264
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 24044 5545 24072 6054
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24030 5536 24086 5545
rect 24030 5471 24086 5480
rect 24030 5264 24086 5273
rect 23848 5228 23900 5234
rect 24030 5199 24086 5208
rect 23848 5170 23900 5176
rect 23572 2644 23624 2650
rect 23572 2586 23624 2592
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 22836 2372 22888 2378
rect 22836 2314 22888 2320
rect 21638 54 22048 82
rect 22650 82 22706 480
rect 22848 82 22876 2314
rect 22650 54 22876 82
rect 23570 82 23626 480
rect 23860 82 23888 5170
rect 23940 5160 23992 5166
rect 23940 5102 23992 5108
rect 23952 4185 23980 5102
rect 24044 4690 24072 5199
rect 24136 4729 24164 5850
rect 24216 5704 24268 5710
rect 24216 5646 24268 5652
rect 24228 5370 24256 5646
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24122 4720 24178 4729
rect 24032 4684 24084 4690
rect 24122 4655 24178 4664
rect 24032 4626 24084 4632
rect 24044 4282 24072 4626
rect 24872 4622 24900 6287
rect 27618 6216 27674 6225
rect 27618 6151 27674 6160
rect 25134 4856 25190 4865
rect 25134 4791 25190 4800
rect 24124 4616 24176 4622
rect 24124 4558 24176 4564
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24032 4276 24084 4282
rect 24032 4218 24084 4224
rect 23938 4176 23994 4185
rect 23938 4111 23994 4120
rect 24136 3602 24164 4558
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 25148 4282 25176 4791
rect 25504 4684 25556 4690
rect 25504 4626 25556 4632
rect 25136 4276 25188 4282
rect 25136 4218 25188 4224
rect 25148 4078 25176 4218
rect 25516 4146 25544 4626
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 27068 4140 27120 4146
rect 27068 4082 27120 4088
rect 25136 4072 25188 4078
rect 25136 4014 25188 4020
rect 25872 4072 25924 4078
rect 25872 4014 25924 4020
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25516 3670 25544 3878
rect 25504 3664 25556 3670
rect 25504 3606 25556 3612
rect 24124 3596 24176 3602
rect 24124 3538 24176 3544
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 24136 3126 24164 3538
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 24688 2854 24716 3538
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 24676 2848 24728 2854
rect 24676 2790 24728 2796
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 24044 2009 24072 2450
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24030 2000 24086 2009
rect 24030 1935 24086 1944
rect 23570 54 23888 82
rect 24582 82 24638 480
rect 24872 82 24900 2926
rect 24582 54 24900 82
rect 25502 82 25558 480
rect 25884 82 25912 4014
rect 26148 2848 26200 2854
rect 26148 2790 26200 2796
rect 25502 54 25912 82
rect 26160 82 26188 2790
rect 26514 82 26570 480
rect 26160 54 26570 82
rect 27080 82 27108 4082
rect 27632 2281 27660 6151
rect 27618 2272 27674 2281
rect 27618 2207 27674 2216
rect 27434 82 27490 480
rect 27080 54 27490 82
rect 19706 0 19762 54
rect 20718 0 20774 54
rect 21638 0 21694 54
rect 22650 0 22706 54
rect 23570 0 23626 54
rect 24582 0 24638 54
rect 25502 0 25558 54
rect 26514 0 26570 54
rect 27434 0 27490 54
<< via2 >>
rect 1214 24792 1270 24848
rect 110 23568 166 23624
rect 110 21800 166 21856
rect 110 19216 166 19272
rect 1582 15952 1638 16008
rect 110 13096 166 13152
rect 1582 14320 1638 14376
rect 2042 11192 2098 11248
rect 4710 26560 4766 26616
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 3422 17720 3478 17776
rect 1950 9696 2006 9752
rect 3974 10784 4030 10840
rect 3422 9560 3478 9616
rect 4158 9696 4214 9752
rect 1398 9016 1454 9072
rect 1398 7792 1454 7848
rect 1582 7520 1638 7576
rect 1490 6568 1546 6624
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5262 13776 5318 13832
rect 5170 10648 5226 10704
rect 5170 9696 5226 9752
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 9034 24792 9090 24848
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 8574 19760 8630 19816
rect 11334 19216 11390 19272
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 8114 13388 8170 13424
rect 8114 13368 8116 13388
rect 8116 13368 8168 13388
rect 8168 13368 8170 13388
rect 8206 13232 8262 13288
rect 8390 12824 8446 12880
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5538 7248 5594 7304
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5906 2352 5962 2408
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 8758 13096 8814 13152
rect 8758 11600 8814 11656
rect 8666 8880 8722 8936
rect 6826 4120 6882 4176
rect 6918 3984 6974 4040
rect 6550 3576 6606 3632
rect 6182 2896 6238 2952
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 9632 13772 9688 13828
rect 9494 13368 9550 13424
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15934 24792 15990 24848
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 10782 13232 10838 13288
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 11978 12688 12034 12744
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 7562 4392 7618 4448
rect 7746 3440 7802 3496
rect 7470 1672 7526 1728
rect 8022 1400 8078 1456
rect 8942 5752 8998 5808
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10690 6160 10746 6216
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10414 4528 10470 4584
rect 10138 4120 10194 4176
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 12438 13368 12494 13424
rect 13358 17720 13414 17776
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 12622 13232 12678 13288
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14278 13096 14334 13152
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15382 12824 15438 12880
rect 16578 12824 16634 12880
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 13542 8744 13598 8800
rect 12254 6704 12310 6760
rect 11978 4120 12034 4176
rect 11978 3596 12034 3632
rect 11978 3576 11980 3596
rect 11980 3576 12032 3596
rect 12032 3576 12034 3596
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14002 8880 14058 8936
rect 14186 9424 14242 9480
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15934 9968 15990 10024
rect 13634 6296 13690 6352
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14094 7792 14150 7848
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 16762 11192 16818 11248
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15382 6568 15438 6624
rect 12438 3440 12494 3496
rect 11334 584 11390 640
rect 11978 40 12034 96
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14738 4664 14794 4720
rect 14922 4528 14978 4584
rect 14738 4392 14794 4448
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14462 3032 14518 3088
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15290 2488 15346 2544
rect 14646 2352 14702 2408
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 13450 1944 13506 2000
rect 16394 7248 16450 7304
rect 15474 3712 15530 3768
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 18602 17720 18658 17776
rect 17222 9968 17278 10024
rect 18234 15952 18290 16008
rect 17682 11600 17738 11656
rect 18694 15408 18750 15464
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 18694 10920 18750 10976
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19062 10648 19118 10704
rect 17314 9696 17370 9752
rect 17498 8472 17554 8528
rect 16302 2896 16358 2952
rect 16578 3440 16634 3496
rect 17130 1944 17186 2000
rect 16854 1672 16910 1728
rect 18786 9560 18842 9616
rect 17774 5752 17830 5808
rect 18970 5480 19026 5536
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19062 5208 19118 5264
rect 18878 4664 18934 4720
rect 19062 4664 19118 4720
rect 17774 3576 17830 3632
rect 18694 3984 18750 4040
rect 21914 12824 21970 12880
rect 22098 20304 22154 20360
rect 23294 25200 23350 25256
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 22466 14320 22522 14376
rect 22374 12688 22430 12744
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19246 3712 19302 3768
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20902 6568 20958 6624
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 22190 9696 22246 9752
rect 22098 8880 22154 8936
rect 21914 8472 21970 8528
rect 21362 3576 21418 3632
rect 21454 2488 21510 2544
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24674 21936 24730 21992
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24766 18808 24822 18864
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 22926 17176 22982 17232
rect 22374 3984 22430 4040
rect 22834 3984 22890 4040
rect 23386 9968 23442 10024
rect 23754 10920 23810 10976
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24214 15952 24270 16008
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 25134 26560 25190 26616
rect 25134 23432 25190 23488
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 27618 13096 27674 13152
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24766 8744 24822 8800
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 23478 3440 23534 3496
rect 22374 3032 22430 3088
rect 24214 6704 24270 6760
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 25410 11056 25466 11112
rect 25042 8472 25098 8528
rect 27618 6840 27674 6896
rect 24858 6296 24914 6352
rect 24030 5480 24086 5536
rect 24030 5208 24086 5264
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24122 4664 24178 4720
rect 27618 6160 27674 6216
rect 25134 4800 25190 4856
rect 23938 4120 23994 4176
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24030 1944 24086 2000
rect 27618 2216 27674 2272
<< metal3 >>
rect 0 27072 480 27192
rect 27520 27072 28000 27192
rect 62 26618 122 27072
rect 4705 26618 4771 26621
rect 62 26616 4771 26618
rect 62 26560 4710 26616
rect 4766 26560 4771 26616
rect 62 26558 4771 26560
rect 4705 26555 4771 26558
rect 25129 26618 25195 26621
rect 27662 26618 27722 27072
rect 25129 26616 27722 26618
rect 25129 26560 25134 26616
rect 25190 26560 27722 26616
rect 25129 26558 27722 26560
rect 25129 26555 25195 26558
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 27520 25576 28000 25696
rect 19610 25535 19930 25536
rect 0 25304 480 25424
rect 62 24850 122 25304
rect 23289 25258 23355 25261
rect 27662 25258 27722 25576
rect 23289 25256 27722 25258
rect 23289 25200 23294 25256
rect 23350 25200 27722 25256
rect 23289 25198 27722 25200
rect 23289 25195 23355 25198
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 1209 24850 1275 24853
rect 62 24848 1275 24850
rect 62 24792 1214 24848
rect 1270 24792 1275 24848
rect 62 24790 1275 24792
rect 1209 24787 1275 24790
rect 9029 24850 9095 24853
rect 15929 24850 15995 24853
rect 9029 24848 15995 24850
rect 9029 24792 9034 24848
rect 9090 24792 15934 24848
rect 15990 24792 15995 24848
rect 9029 24790 15995 24792
rect 9029 24787 9095 24790
rect 15929 24787 15995 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 27520 23944 28000 24064
rect 24277 23903 24597 23904
rect 0 23624 480 23656
rect 0 23568 110 23624
rect 166 23568 480 23624
rect 0 23536 480 23568
rect 25129 23490 25195 23493
rect 27662 23490 27722 23944
rect 25129 23488 27722 23490
rect 25129 23432 25134 23488
rect 25190 23432 27722 23488
rect 25129 23430 27722 23432
rect 25129 23427 25195 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 27520 22448 28000 22568
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 24669 21994 24735 21997
rect 27662 21994 27722 22448
rect 24669 21992 27722 21994
rect 24669 21936 24674 21992
rect 24730 21936 27722 21992
rect 24669 21934 27722 21936
rect 24669 21931 24735 21934
rect 0 21856 480 21888
rect 0 21800 110 21856
rect 166 21800 480 21856
rect 0 21768 480 21800
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 27520 20816 28000 20936
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 22093 20362 22159 20365
rect 27662 20362 27722 20816
rect 22093 20360 27722 20362
rect 22093 20304 22098 20360
rect 22154 20304 27722 20360
rect 22093 20302 27722 20304
rect 22093 20299 22159 20302
rect 10277 20160 10597 20161
rect 0 20000 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 62 19818 122 20000
rect 8569 19818 8635 19821
rect 62 19816 8635 19818
rect 62 19760 8574 19816
rect 8630 19760 8635 19816
rect 62 19758 8635 19760
rect 8569 19755 8635 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 27520 19320 28000 19440
rect 105 19274 171 19277
rect 11329 19274 11395 19277
rect 105 19272 11395 19274
rect 105 19216 110 19272
rect 166 19216 11334 19272
rect 11390 19216 11395 19272
rect 105 19214 11395 19216
rect 105 19211 171 19214
rect 11329 19211 11395 19214
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 24761 18866 24827 18869
rect 27662 18866 27722 19320
rect 24761 18864 27722 18866
rect 24761 18808 24766 18864
rect 24822 18808 27722 18864
rect 24761 18806 27722 18808
rect 24761 18803 24827 18806
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 0 18232 480 18352
rect 62 17778 122 18232
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 3417 17778 3483 17781
rect 62 17776 3483 17778
rect 62 17720 3422 17776
rect 3478 17720 3483 17776
rect 62 17718 3483 17720
rect 3417 17715 3483 17718
rect 13353 17778 13419 17781
rect 18597 17778 18663 17781
rect 13353 17776 18663 17778
rect 13353 17720 13358 17776
rect 13414 17720 18602 17776
rect 18658 17720 18663 17776
rect 13353 17718 18663 17720
rect 13353 17715 13419 17718
rect 18597 17715 18663 17718
rect 27520 17688 28000 17808
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 22921 17234 22987 17237
rect 27662 17234 27722 17688
rect 22921 17232 27722 17234
rect 22921 17176 22926 17232
rect 22982 17176 27722 17232
rect 22921 17174 27722 17176
rect 22921 17171 22987 17174
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 0 16464 480 16584
rect 62 16010 122 16464
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 27520 16192 28000 16312
rect 1577 16010 1643 16013
rect 62 16008 1643 16010
rect 62 15952 1582 16008
rect 1638 15952 1643 16008
rect 62 15950 1643 15952
rect 1577 15947 1643 15950
rect 18229 16010 18295 16013
rect 24209 16010 24275 16013
rect 18229 16008 24275 16010
rect 18229 15952 18234 16008
rect 18290 15952 24214 16008
rect 24270 15952 24275 16008
rect 18229 15950 24275 15952
rect 18229 15947 18295 15950
rect 24209 15947 24275 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 18689 15466 18755 15469
rect 27662 15466 27722 16192
rect 18689 15464 27722 15466
rect 18689 15408 18694 15464
rect 18750 15408 27722 15464
rect 18689 15406 27722 15408
rect 18689 15403 18755 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 0 14832 480 14952
rect 62 14378 122 14832
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 27520 14696 28000 14816
rect 19610 14655 19930 14656
rect 1577 14378 1643 14381
rect 62 14376 1643 14378
rect 62 14320 1582 14376
rect 1638 14320 1643 14376
rect 62 14318 1643 14320
rect 1577 14315 1643 14318
rect 22461 14378 22527 14381
rect 27662 14378 27722 14696
rect 22461 14376 27722 14378
rect 22461 14320 22466 14376
rect 22522 14320 27722 14376
rect 22461 14318 27722 14320
rect 22461 14315 22527 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 5257 13834 5323 13837
rect 5257 13833 9690 13834
rect 5257 13832 9693 13833
rect 5257 13776 5262 13832
rect 5318 13828 9693 13832
rect 5318 13776 9632 13828
rect 5257 13774 9632 13776
rect 5257 13771 5323 13774
rect 9627 13772 9632 13774
rect 9688 13772 9693 13828
rect 9627 13767 9693 13772
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 8109 13426 8175 13429
rect 9489 13426 9555 13429
rect 12433 13426 12499 13429
rect 8109 13424 12499 13426
rect 8109 13368 8114 13424
rect 8170 13368 9494 13424
rect 9550 13368 12438 13424
rect 12494 13368 12499 13424
rect 8109 13366 12499 13368
rect 8109 13363 8175 13366
rect 9489 13363 9555 13366
rect 12433 13363 12499 13366
rect 8201 13290 8267 13293
rect 10777 13290 10843 13293
rect 12617 13290 12683 13293
rect 8201 13288 12683 13290
rect 8201 13232 8206 13288
rect 8262 13232 10782 13288
rect 10838 13232 12622 13288
rect 12678 13232 12683 13288
rect 8201 13230 12683 13232
rect 8201 13227 8267 13230
rect 10777 13227 10843 13230
rect 12617 13227 12683 13230
rect 0 13152 480 13184
rect 0 13096 110 13152
rect 166 13096 480 13152
rect 0 13064 480 13096
rect 8753 13154 8819 13157
rect 14273 13154 14339 13157
rect 8753 13152 14339 13154
rect 8753 13096 8758 13152
rect 8814 13096 14278 13152
rect 14334 13096 14339 13152
rect 8753 13094 14339 13096
rect 8753 13091 8819 13094
rect 14273 13091 14339 13094
rect 27520 13152 28000 13184
rect 27520 13096 27618 13152
rect 27674 13096 28000 13152
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13096
rect 24277 13023 24597 13024
rect 8385 12882 8451 12885
rect 15377 12882 15443 12885
rect 8385 12880 15443 12882
rect 8385 12824 8390 12880
rect 8446 12824 15382 12880
rect 15438 12824 15443 12880
rect 8385 12822 15443 12824
rect 8385 12819 8451 12822
rect 15377 12819 15443 12822
rect 16573 12882 16639 12885
rect 21909 12882 21975 12885
rect 16573 12880 21975 12882
rect 16573 12824 16578 12880
rect 16634 12824 21914 12880
rect 21970 12824 21975 12880
rect 16573 12822 21975 12824
rect 16573 12819 16639 12822
rect 21909 12819 21975 12822
rect 11973 12746 12039 12749
rect 22369 12746 22435 12749
rect 11973 12744 22435 12746
rect 11973 12688 11978 12744
rect 12034 12688 22374 12744
rect 22430 12688 22435 12744
rect 11973 12686 22435 12688
rect 11973 12683 12039 12686
rect 22369 12683 22435 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 8753 11658 8819 11661
rect 17677 11658 17743 11661
rect 8753 11656 17743 11658
rect 8753 11600 8758 11656
rect 8814 11600 17682 11656
rect 17738 11600 17743 11656
rect 8753 11598 17743 11600
rect 8753 11595 8819 11598
rect 17677 11595 17743 11598
rect 27520 11568 28000 11688
rect 10277 11456 10597 11457
rect 0 11296 480 11416
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 62 10842 122 11296
rect 2037 11250 2103 11253
rect 16757 11250 16823 11253
rect 2037 11248 16823 11250
rect 2037 11192 2042 11248
rect 2098 11192 16762 11248
rect 16818 11192 16823 11248
rect 2037 11190 16823 11192
rect 2037 11187 2103 11190
rect 16757 11187 16823 11190
rect 25405 11114 25471 11117
rect 27662 11114 27722 11568
rect 25405 11112 27722 11114
rect 25405 11056 25410 11112
rect 25466 11056 27722 11112
rect 25405 11054 27722 11056
rect 25405 11051 25471 11054
rect 18689 10978 18755 10981
rect 23749 10978 23815 10981
rect 18689 10976 23815 10978
rect 18689 10920 18694 10976
rect 18750 10920 23754 10976
rect 23810 10920 23815 10976
rect 18689 10918 23815 10920
rect 18689 10915 18755 10918
rect 23749 10915 23815 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 3969 10842 4035 10845
rect 62 10840 4035 10842
rect 62 10784 3974 10840
rect 4030 10784 4035 10840
rect 62 10782 4035 10784
rect 3969 10779 4035 10782
rect 5165 10706 5231 10709
rect 19057 10706 19123 10709
rect 5165 10704 19123 10706
rect 5165 10648 5170 10704
rect 5226 10648 19062 10704
rect 19118 10648 19123 10704
rect 5165 10646 19123 10648
rect 5165 10643 5231 10646
rect 19057 10643 19123 10646
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 15929 10026 15995 10029
rect 17217 10026 17283 10029
rect 23381 10026 23447 10029
rect 15929 10024 23447 10026
rect 15929 9968 15934 10024
rect 15990 9968 17222 10024
rect 17278 9968 23386 10024
rect 23442 9968 23447 10024
rect 15929 9966 23447 9968
rect 15929 9963 15995 9966
rect 17217 9963 17283 9966
rect 23381 9963 23447 9966
rect 27520 9936 28000 10056
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 1945 9754 2011 9757
rect 4153 9754 4219 9757
rect 5165 9754 5231 9757
rect 1945 9752 5231 9754
rect 1945 9696 1950 9752
rect 2006 9696 4158 9752
rect 4214 9696 5170 9752
rect 5226 9696 5231 9752
rect 1945 9694 5231 9696
rect 1945 9691 2011 9694
rect 4153 9691 4219 9694
rect 5165 9691 5231 9694
rect 17309 9754 17375 9757
rect 22185 9754 22251 9757
rect 17309 9752 22251 9754
rect 17309 9696 17314 9752
rect 17370 9696 22190 9752
rect 22246 9696 22251 9752
rect 17309 9694 22251 9696
rect 17309 9691 17375 9694
rect 22185 9691 22251 9694
rect 0 9528 480 9648
rect 3417 9618 3483 9621
rect 18781 9618 18847 9621
rect 3417 9616 18847 9618
rect 3417 9560 3422 9616
rect 3478 9560 18786 9616
rect 18842 9560 18847 9616
rect 3417 9558 18847 9560
rect 3417 9555 3483 9558
rect 18781 9555 18847 9558
rect 62 9074 122 9528
rect 14181 9482 14247 9485
rect 27662 9482 27722 9936
rect 14181 9480 27722 9482
rect 14181 9424 14186 9480
rect 14242 9424 27722 9480
rect 14181 9422 27722 9424
rect 14181 9419 14247 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 1393 9074 1459 9077
rect 62 9072 1459 9074
rect 62 9016 1398 9072
rect 1454 9016 1459 9072
rect 62 9014 1459 9016
rect 1393 9011 1459 9014
rect 8661 8938 8727 8941
rect 9438 8938 9444 8940
rect 8661 8936 9444 8938
rect 8661 8880 8666 8936
rect 8722 8880 9444 8936
rect 8661 8878 9444 8880
rect 8661 8875 8727 8878
rect 9438 8876 9444 8878
rect 9508 8938 9514 8940
rect 13997 8938 14063 8941
rect 22093 8938 22159 8941
rect 9508 8936 14063 8938
rect 9508 8880 14002 8936
rect 14058 8880 14063 8936
rect 9508 8878 14063 8880
rect 9508 8876 9514 8878
rect 13997 8875 14063 8878
rect 14782 8936 22159 8938
rect 14782 8880 22098 8936
rect 22154 8880 22159 8936
rect 14782 8878 22159 8880
rect 13537 8802 13603 8805
rect 14782 8802 14842 8878
rect 22093 8875 22159 8878
rect 13537 8800 14842 8802
rect 13537 8744 13542 8800
rect 13598 8744 14842 8800
rect 13537 8742 14842 8744
rect 24761 8802 24827 8805
rect 27654 8802 27660 8804
rect 24761 8800 27660 8802
rect 24761 8744 24766 8800
rect 24822 8744 27660 8800
rect 24761 8742 27660 8744
rect 13537 8739 13603 8742
rect 24761 8739 24827 8742
rect 27654 8740 27660 8742
rect 27724 8740 27730 8804
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 17493 8530 17559 8533
rect 21909 8530 21975 8533
rect 25037 8530 25103 8533
rect 17493 8528 25103 8530
rect 17493 8472 17498 8528
rect 17554 8472 21914 8528
rect 21970 8472 25042 8528
rect 25098 8472 25103 8528
rect 17493 8470 25103 8472
rect 17493 8467 17559 8470
rect 21909 8467 21975 8470
rect 25037 8467 25103 8470
rect 27520 8532 28000 8560
rect 27520 8468 27660 8532
rect 27724 8468 28000 8532
rect 27520 8440 28000 8468
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 0 7760 480 7880
rect 1393 7850 1459 7853
rect 14089 7850 14155 7853
rect 1393 7848 14155 7850
rect 1393 7792 1398 7848
rect 1454 7792 14094 7848
rect 14150 7792 14155 7848
rect 1393 7790 14155 7792
rect 1393 7787 1459 7790
rect 14089 7787 14155 7790
rect 62 7578 122 7760
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 1577 7578 1643 7581
rect 62 7576 1643 7578
rect 62 7520 1582 7576
rect 1638 7520 1643 7576
rect 62 7518 1643 7520
rect 1577 7515 1643 7518
rect 5533 7306 5599 7309
rect 16389 7306 16455 7309
rect 5533 7304 16455 7306
rect 5533 7248 5538 7304
rect 5594 7248 16394 7304
rect 16450 7248 16455 7304
rect 5533 7246 16455 7248
rect 5533 7243 5599 7246
rect 16389 7243 16455 7246
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 27520 6896 28000 6928
rect 27520 6840 27618 6896
rect 27674 6840 28000 6896
rect 27520 6808 28000 6840
rect 12249 6762 12315 6765
rect 24209 6762 24275 6765
rect 12249 6760 24275 6762
rect 12249 6704 12254 6760
rect 12310 6704 24214 6760
rect 24270 6704 24275 6760
rect 12249 6702 24275 6704
rect 12249 6699 12315 6702
rect 24209 6699 24275 6702
rect 1485 6626 1551 6629
rect 62 6624 1551 6626
rect 62 6568 1490 6624
rect 1546 6568 1551 6624
rect 62 6566 1551 6568
rect 62 6112 122 6566
rect 1485 6563 1551 6566
rect 15377 6626 15443 6629
rect 20897 6626 20963 6629
rect 15377 6624 20963 6626
rect 15377 6568 15382 6624
rect 15438 6568 20902 6624
rect 20958 6568 20963 6624
rect 15377 6566 20963 6568
rect 15377 6563 15443 6566
rect 20897 6563 20963 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 238 6292 244 6356
rect 308 6354 314 6356
rect 13629 6354 13695 6357
rect 24853 6354 24919 6357
rect 308 6352 24919 6354
rect 308 6296 13634 6352
rect 13690 6296 24858 6352
rect 24914 6296 24919 6352
rect 308 6294 24919 6296
rect 308 6292 314 6294
rect 13629 6291 13695 6294
rect 24853 6291 24919 6294
rect 10685 6218 10751 6221
rect 27613 6218 27679 6221
rect 10685 6216 27679 6218
rect 10685 6160 10690 6216
rect 10746 6160 27618 6216
rect 27674 6160 27679 6216
rect 10685 6158 27679 6160
rect 10685 6155 10751 6158
rect 27613 6155 27679 6158
rect 0 5992 480 6112
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 8937 5810 9003 5813
rect 17769 5810 17835 5813
rect 8937 5808 17835 5810
rect 8937 5752 8942 5808
rect 8998 5752 17774 5808
rect 17830 5752 17835 5808
rect 8937 5750 17835 5752
rect 8937 5747 9003 5750
rect 17769 5747 17835 5750
rect 18965 5538 19031 5541
rect 24025 5538 24091 5541
rect 18965 5536 24091 5538
rect 18965 5480 18970 5536
rect 19026 5480 24030 5536
rect 24086 5480 24091 5536
rect 18965 5478 24091 5480
rect 18965 5475 19031 5478
rect 24025 5475 24091 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 27520 5312 28000 5432
rect 19057 5266 19123 5269
rect 24025 5266 24091 5269
rect 19057 5264 24091 5266
rect 19057 5208 19062 5264
rect 19118 5208 24030 5264
rect 24086 5208 24091 5264
rect 19057 5206 24091 5208
rect 19057 5203 19123 5206
rect 24025 5203 24091 5206
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 25129 4858 25195 4861
rect 27662 4858 27722 5312
rect 25129 4856 27722 4858
rect 25129 4800 25134 4856
rect 25190 4800 27722 4856
rect 25129 4798 27722 4800
rect 25129 4795 25195 4798
rect 14733 4722 14799 4725
rect 18873 4722 18939 4725
rect 14733 4720 18939 4722
rect 14733 4664 14738 4720
rect 14794 4664 18878 4720
rect 18934 4664 18939 4720
rect 14733 4662 18939 4664
rect 14733 4659 14799 4662
rect 18873 4659 18939 4662
rect 19057 4722 19123 4725
rect 24117 4722 24183 4725
rect 19057 4720 24183 4722
rect 19057 4664 19062 4720
rect 19118 4664 24122 4720
rect 24178 4664 24183 4720
rect 19057 4662 24183 4664
rect 19057 4659 19123 4662
rect 24117 4659 24183 4662
rect 10409 4586 10475 4589
rect 14917 4586 14983 4589
rect 10409 4584 14983 4586
rect 10409 4528 10414 4584
rect 10470 4528 14922 4584
rect 14978 4528 14983 4584
rect 10409 4526 14983 4528
rect 10409 4523 10475 4526
rect 14917 4523 14983 4526
rect 7557 4450 7623 4453
rect 14733 4450 14799 4453
rect 7557 4448 14799 4450
rect 7557 4392 7562 4448
rect 7618 4392 14738 4448
rect 14794 4392 14799 4448
rect 7557 4390 14799 4392
rect 7557 4387 7623 4390
rect 14733 4387 14799 4390
rect 5610 4384 5930 4385
rect 0 4316 480 4344
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 0 4252 60 4316
rect 124 4252 480 4316
rect 0 4224 480 4252
rect 6821 4178 6887 4181
rect 10133 4178 10199 4181
rect 6821 4176 10199 4178
rect 6821 4120 6826 4176
rect 6882 4120 10138 4176
rect 10194 4120 10199 4176
rect 6821 4118 10199 4120
rect 6821 4115 6887 4118
rect 10133 4115 10199 4118
rect 11973 4178 12039 4181
rect 23933 4178 23999 4181
rect 11973 4176 23999 4178
rect 11973 4120 11978 4176
rect 12034 4120 23938 4176
rect 23994 4120 23999 4176
rect 11973 4118 23999 4120
rect 11973 4115 12039 4118
rect 23933 4115 23999 4118
rect 6913 4042 6979 4045
rect 9438 4042 9444 4044
rect 6913 4040 9444 4042
rect 6913 3984 6918 4040
rect 6974 3984 9444 4040
rect 6913 3982 9444 3984
rect 6913 3979 6979 3982
rect 9438 3980 9444 3982
rect 9508 3980 9514 4044
rect 18689 4042 18755 4045
rect 22369 4042 22435 4045
rect 18689 4040 22435 4042
rect 18689 3984 18694 4040
rect 18750 3984 22374 4040
rect 22430 3984 22435 4040
rect 18689 3982 22435 3984
rect 18689 3979 18755 3982
rect 22369 3979 22435 3982
rect 22829 4042 22895 4045
rect 22829 4040 27722 4042
rect 22829 3984 22834 4040
rect 22890 3984 27722 4040
rect 22829 3982 27722 3984
rect 22829 3979 22895 3982
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 27662 3800 27722 3982
rect 19610 3775 19930 3776
rect 15469 3770 15535 3773
rect 19241 3770 19307 3773
rect 15469 3768 19307 3770
rect 15469 3712 15474 3768
rect 15530 3712 19246 3768
rect 19302 3712 19307 3768
rect 15469 3710 19307 3712
rect 15469 3707 15535 3710
rect 19241 3707 19307 3710
rect 27520 3680 28000 3800
rect 6545 3634 6611 3637
rect 11973 3634 12039 3637
rect 6545 3632 12039 3634
rect 6545 3576 6550 3632
rect 6606 3576 11978 3632
rect 12034 3576 12039 3632
rect 6545 3574 12039 3576
rect 6545 3571 6611 3574
rect 11973 3571 12039 3574
rect 17769 3634 17835 3637
rect 21357 3634 21423 3637
rect 17769 3632 21423 3634
rect 17769 3576 17774 3632
rect 17830 3576 21362 3632
rect 21418 3576 21423 3632
rect 17769 3574 21423 3576
rect 17769 3571 17835 3574
rect 21357 3571 21423 3574
rect 7741 3498 7807 3501
rect 12433 3498 12499 3501
rect 7741 3496 12499 3498
rect 7741 3440 7746 3496
rect 7802 3440 12438 3496
rect 12494 3440 12499 3496
rect 7741 3438 12499 3440
rect 7741 3435 7807 3438
rect 12433 3435 12499 3438
rect 16573 3498 16639 3501
rect 23473 3498 23539 3501
rect 16573 3496 23539 3498
rect 16573 3440 16578 3496
rect 16634 3440 23478 3496
rect 23534 3440 23539 3496
rect 16573 3438 23539 3440
rect 16573 3435 16639 3438
rect 23473 3435 23539 3438
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 14457 3090 14523 3093
rect 22369 3090 22435 3093
rect 14457 3088 22435 3090
rect 14457 3032 14462 3088
rect 14518 3032 22374 3088
rect 22430 3032 22435 3088
rect 14457 3030 22435 3032
rect 14457 3027 14523 3030
rect 22369 3027 22435 3030
rect 6177 2954 6243 2957
rect 16297 2954 16363 2957
rect 6177 2952 16363 2954
rect 6177 2896 6182 2952
rect 6238 2896 16302 2952
rect 16358 2896 16363 2952
rect 6177 2894 16363 2896
rect 6177 2891 6243 2894
rect 16297 2891 16363 2894
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 0 2456 480 2576
rect 15285 2546 15351 2549
rect 21449 2546 21515 2549
rect 15285 2544 21515 2546
rect 15285 2488 15290 2544
rect 15346 2488 21454 2544
rect 21510 2488 21515 2544
rect 15285 2486 21515 2488
rect 15285 2483 15351 2486
rect 21449 2483 21515 2486
rect 62 2002 122 2456
rect 5901 2410 5967 2413
rect 14641 2410 14707 2413
rect 5901 2408 14707 2410
rect 5901 2352 5906 2408
rect 5962 2352 14646 2408
rect 14702 2352 14707 2408
rect 5901 2350 14707 2352
rect 5901 2347 5967 2350
rect 14641 2347 14707 2350
rect 27520 2272 28000 2304
rect 27520 2216 27618 2272
rect 27674 2216 28000 2272
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 27520 2184 28000 2216
rect 24277 2143 24597 2144
rect 13445 2002 13511 2005
rect 62 2000 13511 2002
rect 62 1944 13450 2000
rect 13506 1944 13511 2000
rect 62 1942 13511 1944
rect 13445 1939 13511 1942
rect 17125 2002 17191 2005
rect 24025 2002 24091 2005
rect 17125 2000 24091 2002
rect 17125 1944 17130 2000
rect 17186 1944 24030 2000
rect 24086 1944 24091 2000
rect 17125 1942 24091 1944
rect 17125 1939 17191 1942
rect 24025 1939 24091 1942
rect 7465 1730 7531 1733
rect 16849 1730 16915 1733
rect 7465 1728 16915 1730
rect 7465 1672 7470 1728
rect 7526 1672 16854 1728
rect 16910 1672 16915 1728
rect 7465 1670 16915 1672
rect 7465 1667 7531 1670
rect 16849 1667 16915 1670
rect 8017 1458 8083 1461
rect 62 1456 8083 1458
rect 62 1400 8022 1456
rect 8078 1400 8083 1456
rect 62 1398 8083 1400
rect 62 944 122 1398
rect 8017 1395 8083 1398
rect 0 824 480 944
rect 27520 780 28000 808
rect 27520 716 27660 780
rect 27724 716 28000 780
rect 27520 688 28000 716
rect 11329 642 11395 645
rect 11329 640 19350 642
rect 11329 584 11334 640
rect 11390 584 19350 640
rect 11329 582 19350 584
rect 11329 579 11395 582
rect 19290 506 19350 582
rect 27654 506 27660 508
rect 19290 446 27660 506
rect 27654 444 27660 446
rect 27724 444 27730 508
rect 9622 36 9628 100
rect 9692 98 9698 100
rect 11973 98 12039 101
rect 9692 96 12039 98
rect 9692 40 11978 96
rect 12034 40 12039 96
rect 9692 38 12039 40
rect 9692 36 9698 38
rect 11973 35 12039 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 9444 8876 9508 8940
rect 27660 8740 27724 8804
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 27660 8468 27724 8532
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 244 6292 308 6356
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 60 4252 124 4316
rect 9444 3980 9508 4044
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 27660 716 27724 780
rect 27660 444 27724 508
rect 9628 36 9692 100
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 9443 8940 9509 8941
rect 9443 8876 9444 8940
rect 9508 8876 9509 8940
rect 9443 8875 9509 8876
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 243 6356 309 6357
rect 243 6292 244 6356
rect 308 6292 309 6356
rect 243 6291 309 6292
rect 246 5130 306 6291
rect 62 5070 306 5130
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 62 4317 122 5070
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 59 4316 125 4317
rect 59 4252 60 4316
rect 124 4252 125 4316
rect 59 4251 125 4252
rect 5610 3296 5931 4320
rect 9446 4170 9506 8875
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 9446 4110 9690 4170
rect 9446 4045 9506 4110
rect 9443 4044 9509 4045
rect 9443 3980 9444 4044
rect 9508 3980 9509 4044
rect 9443 3979 9509 3980
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 9630 101 9690 4110
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 27659 8804 27725 8805
rect 27659 8740 27660 8804
rect 27724 8740 27725 8804
rect 27659 8739 27725 8740
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 27662 8533 27722 8739
rect 27659 8532 27725 8533
rect 27659 8468 27660 8532
rect 27724 8468 27725 8532
rect 27659 8467 27725 8468
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 27659 780 27725 781
rect 27659 716 27660 780
rect 27724 716 27725 780
rect 27659 715 27725 716
rect 27662 509 27722 715
rect 27659 508 27725 509
rect 27659 444 27660 508
rect 27724 444 27725 508
rect 27659 443 27725 444
rect 9627 100 9693 101
rect 9627 36 9628 100
rect 9692 36 9693 100
rect 9627 35 9693 36
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_0_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_conb_1  _132_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_43 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_47
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_42
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _142_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 7544 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_85
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_81
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use scs8hd_nor4_4  _115_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 1602 592
use scs8hd_inv_8  _044_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _043_
timestamp 1586364061
transform 1 0 7728 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_91
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_106
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_115
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_111
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__D
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__C
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_120
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_119
timestamp 1586364061
transform 1 0 12052 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_140
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_134
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_148
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_144
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_158
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_154
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_152 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15088 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_162
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_177
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _161_
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_181
timestamp 1586364061
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_181
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_202
timestamp 1586364061
transform 1 0 19688 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_198
timestamp 1586364061
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_202
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_215
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_219
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_236 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _154_
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_243
timestamp 1586364061
transform 1 0 23460 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_239
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_248
timestamp 1586364061
transform 1 0 23920 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_252
timestamp 1586364061
transform 1 0 24288 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_256
timestamp 1586364061
transform 1 0 24656 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_252
timestamp 1586364061
transform 1 0 24288 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_259
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_267
timestamp 1586364061
transform 1 0 25668 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_263
timestamp 1586364061
transform 1 0 25300 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_275
timestamp 1586364061
transform 1 0 26404 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_conb_1  _135_
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _141_
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__064__C
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_55
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_4  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_2  _139_
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__C
timestamp 1586364061
transform 1 0 8924 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_73
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_81
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_87
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _116_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_2  _151_
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_110
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_114
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_130
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_172
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 17572 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_196
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _149_
timestamp 1586364061
transform 1 0 19320 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_235
timestamp 1586364061
transform 1 0 22724 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_246
timestamp 1586364061
transform 1 0 23736 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24472 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_257
timestamp 1586364061
transform 1 0 24748 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_269
timestamp 1586364061
transform 1 0 25852 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_70
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _049_
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__D
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_83
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_87
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _117_
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 1602 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__C
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__D
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_108
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_149
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_153
timestamp 1586364061
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_166
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18952 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18768 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_190
timestamp 1586364061
transform 1 0 18584 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _046_
timestamp 1586364061
transform 1 0 20700 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_205
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_209
timestamp 1586364061
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_222
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_226
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_233
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_237
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_241
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_251
timestamp 1586364061
transform 1 0 24196 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_262
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_273
timestamp 1586364061
transform 1 0 26220 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_6  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 590 592
use scs8hd_or3_4  _064_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_89
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use scs8hd_nor4_4  _114_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_127
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 314 592
use scs8hd_buf_2  _155_
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_148
timestamp 1586364061
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_162
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_181
timestamp 1586364061
transform 1 0 17756 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19504 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_198
timestamp 1586364061
transform 1 0 19320 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _073_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _069_
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_241
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_252
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_56
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__C
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 866 592
use scs8hd_or3_4  _058_
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__058__C
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_79
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_83
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _048_
timestamp 1586364061
transform 1 0 10672 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__060__B
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_96
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_100
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11868 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_5_119
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_141
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_145
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_158
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_162
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18584 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20332 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_201
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_205
timestamp 1586364061
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 21896 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_218
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_222
timestamp 1586364061
transform 1 0 21528 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 22908 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_235
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_239
timestamp 1586364061
transform 1 0 23092 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_248
timestamp 1586364061
transform 1 0 23920 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_252
timestamp 1586364061
transform 1 0 24288 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_259
timestamp 1586364061
transform 1 0 24932 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_263
timestamp 1586364061
transform 1 0 25300 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_275
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_or3_4  _062_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_46
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_50
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_3  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_67
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_or3_4  _068_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_or3_4  _066_
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 866 592
use scs8hd_or3_4  _054_
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_nor4_4  _112_
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__D
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__C
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_96
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__C
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_100
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_107
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use scs8hd_or3_4  _060_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_111
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_128
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_134
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_128
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_160
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_164
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_165
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_173
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_192
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18952 0 -1 5984
box -38 -48 1050 592
use scs8hd_inv_8  _045_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_7_201
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_211
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_209
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19688 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_228
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_228
timestamp 1586364061
transform 1 0 22080 0 1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_7_238
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_234
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_248
timestamp 1586364061
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_241
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use scs8hd_nor2_4  _071_
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 24012 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_252
timestamp 1586364061
transform 1 0 24288 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_267
timestamp 1586364061
transform 1 0 25668 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_263
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_259
timestamp 1586364061
transform 1 0 24932 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_258
timestamp 1586364061
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_270
timestamp 1586364061
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _144_
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_52
timestamp 1586364061
transform 1 0 5888 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_71
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__112__C
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_85
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_103
timestamp 1586364061
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_118
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_122
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_1  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_135
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_2  _158_
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_161
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_189
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _074_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_228
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_235
timestamp 1586364061
transform 1 0 22724 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_8  FILLER_8_246
timestamp 1586364061
transform 1 0 23736 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_2  _140_
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_254
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_259
timestamp 1586364061
transform 1 0 24932 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _143_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 590 592
use scs8hd_inv_8  _041_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__041__A
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_41
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 406 592
use scs8hd_inv_8  _053_
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_104
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_139
timestamp 1586364061
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_152
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_172
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_176
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_214
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_227
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_231
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_234
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_242
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_54
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_8  _052_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use scs8hd_or3_4  _118_
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_97
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_101
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_111
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_115
timestamp 1586364061
transform 1 0 11684 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_118
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_158
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16192 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_175
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17940 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_194
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_228
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_235
timestamp 1586364061
transform 1 0 22724 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_259
timestamp 1586364061
transform 1 0 24932 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_271
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use scs8hd_nor4_4  _113_
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__113__D
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__C
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_77
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__D
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_102
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_106
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 314 592
use scs8hd_conb_1  _133_
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_161
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_165
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_172
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_176
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_190
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_194
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_209
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_226
timestamp 1586364061
transform 1 0 21896 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_230
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_242
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 774 592
use scs8hd_buf_2  _138_
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_253
timestamp 1586364061
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_259
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_263
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_275
timestamp 1586364061
transform 1 0 26404 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use scs8hd_conb_1  _134_
timestamp 1586364061
transform 1 0 4508 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_40
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _042_
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__055__C
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_63
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__D
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_76
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_or4_4  _083_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__D
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__C
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 11316 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_120
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_124
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_128
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_138
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_142
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_6  FILLER_12_176
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 17940 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_185
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_207
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_228
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 406 592
use scs8hd_conb_1  _125_
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_235
timestamp 1586364061
transform 1 0 22724 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_247
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_259
timestamp 1586364061
transform 1 0 24932 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_271
timestamp 1586364061
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_35
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_66
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_54
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use scs8hd_nand3_4  _055_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 1326 592
use scs8hd_inv_8  _050_
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 866 592
use scs8hd_or4_4  _097_
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__B
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__D
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_76
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_80
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__C
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_106
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_or4_4  _090_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_or3_4  _056_
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_110
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__C
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_116
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_121
timestamp 1586364061
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _137_
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_128
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_132
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_144
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_152
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_165
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_169
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_167
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_179
timestamp 1586364061
transform 1 0 17572 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_196
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_192
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 1050 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 17940 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_203
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_198
timestamp 1586364061
transform 1 0 19320 0 1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use scs8hd_conb_1  _130_
timestamp 1586364061
transform 1 0 19504 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_207
timestamp 1586364061
transform 1 0 20148 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_206
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__061__B
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_223
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_228
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_238
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_234
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_241
timestamp 1586364061
transform 1 0 23276 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_242
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__B
timestamp 1586364061
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_nor2_4  _061_
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_271
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_or2_4  _104_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _105_
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_73
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_90
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_94
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_107
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13340 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_131
timestamp 1586364061
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_150
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_167
timestamp 1586364061
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_176
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _131_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_180
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_187
timestamp 1586364061
transform 1 0 18308 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_210
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_227
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _065_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_233
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_237
timestamp 1586364061
transform 1 0 22908 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_241
timestamp 1586364061
transform 1 0 23276 0 1 10336
box -38 -48 130 592
use scs8hd_buf_2  _152_
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_258
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_266
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_270
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _051_
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__C
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_81
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_85
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 9752 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_103
timestamp 1586364061
transform 1 0 10580 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_107
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 590 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_165
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_169
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_177
timestamp 1586364061
transform 1 0 17388 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_16_187
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_225
timestamp 1586364061
transform 1 0 21804 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_229
timestamp 1586364061
transform 1 0 22172 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22724 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_234
timestamp 1586364061
transform 1 0 22632 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_244
timestamp 1586364061
transform 1 0 23552 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_248
timestamp 1586364061
transform 1 0 23920 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _063_
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 866 592
use scs8hd_fill_1  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_261
timestamp 1586364061
transform 1 0 25116 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_273
timestamp 1586364061
transform 1 0 26220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_or2_4  _082_
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 130 592
use scs8hd_or3_4  _075_
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_78
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_99
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_151
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_155
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_168
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_188
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_192
timestamp 1586364061
transform 1 0 18768 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_211
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_221
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _128_
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_17_265
timestamp 1586364061
transform 1 0 25484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10304 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_134
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_151
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_175
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17664 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_18_191
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19504 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 -1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23644 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_241
timestamp 1586364061
transform 1 0 23276 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_247
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_258
timestamp 1586364061
transform 1 0 24840 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_270
timestamp 1586364061
transform 1 0 25944 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_274
timestamp 1586364061
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_2  _153_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_35
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_47
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_73
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_85
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_90
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_101
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_119
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_128
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_141
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 590 592
use scs8hd_decap_4  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_140
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_158
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _057_
timestamp 1586364061
transform 1 0 15732 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _059_
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 17296 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_162
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_185
timestamp 1586364061
transform 1 0 18124 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_189
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_204
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_208
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_210
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_206
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_225
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_229
timestamp 1586364061
transform 1 0 22172 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_232
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22540 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_248
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_244
timestamp 1586364061
transform 1 0 23552 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23736 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22724 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use scs8hd_buf_2  _150_
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_258
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_266
timestamp 1586364061
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_254
timestamp 1586364061
transform 1 0 24472 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_258
timestamp 1586364061
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_270
timestamp 1586364061
transform 1 0 25944 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_276
timestamp 1586364061
transform 1 0 26496 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_270
timestamp 1586364061
transform 1 0 25944 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  _147_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_23
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_47
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _077_
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_67
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_80
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_84
timestamp 1586364061
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_104
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_140
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_154
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_158
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_162
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_187
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 20792 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 20424 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_212
timestamp 1586364061
transform 1 0 20608 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _091_
timestamp 1586364061
transform 1 0 20976 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 21988 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_225
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_229
timestamp 1586364061
transform 1 0 22172 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_248
timestamp 1586364061
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_252
timestamp 1586364061
transform 1 0 24288 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_256
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_268
timestamp 1586364061
transform 1 0 25760 0 1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_21_276
timestamp 1586364061
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 590 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_74
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_90
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_97
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_101
timestamp 1586364061
transform 1 0 10396 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_113
timestamp 1586364061
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 17020 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_165
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_182
timestamp 1586364061
transform 1 0 17848 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_192
timestamp 1586364061
transform 1 0 18768 0 -1 14688
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _067_
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_241
timestamp 1586364061
transform 1 0 23276 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_252
timestamp 1586364061
transform 1 0 24288 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_264
timestamp 1586364061
transform 1 0 25392 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_272
timestamp 1586364061
transform 1 0 26128 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_19
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_31
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_43
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_23_55
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 590 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_85
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_100
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_104
timestamp 1586364061
transform 1 0 10672 0 1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _081_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_108
timestamp 1586364061
transform 1 0 11040 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_137
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_187
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_191
timestamp 1586364061
transform 1 0 18676 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_206
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_210
timestamp 1586364061
transform 1 0 20424 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_225
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_229
timestamp 1586364061
transform 1 0 22172 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_233
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_237
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_243
timestamp 1586364061
transform 1 0 23460 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_buf_2  _146_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_76
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_110
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_120
timestamp 1586364061
transform 1 0 12144 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_128
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_132
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use scs8hd_conb_1  _129_
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_167
timestamp 1586364061
transform 1 0 16468 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_174
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19136 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_182
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_194
timestamp 1586364061
transform 1 0 18952 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_198
timestamp 1586364061
transform 1 0 19320 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_6  FILLER_24_205
timestamp 1586364061
transform 1 0 19964 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_211
timestamp 1586364061
transform 1 0 20516 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_224
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_234
timestamp 1586364061
transform 1 0 22632 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_246
timestamp 1586364061
transform 1 0 23736 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_258
timestamp 1586364061
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_270
timestamp 1586364061
transform 1 0 25944 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_274
timestamp 1586364061
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 6440 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_60
timestamp 1586364061
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_66
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_70
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 8280 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_73
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_87
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_91
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_104
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_108
timestamp 1586364061
transform 1 0 11040 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_112
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_141
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_152
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_165
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_169
timestamp 1586364061
transform 1 0 16652 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_195
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_199
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_206
timestamp 1586364061
transform 1 0 20056 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_210
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22356 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_223
timestamp 1586364061
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_227
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_234
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_238
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_242
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_67
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 1050 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_104
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_93
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_99
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_112
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_108
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_122
timestamp 1586364061
transform 1 0 12328 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14076 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_126
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_134
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_152
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 17020 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_165
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_169
timestamp 1586364061
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_173
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_178
timestamp 1586364061
transform 1 0 17480 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_187
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_182
timestamp 1586364061
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_186
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_182
timestamp 1586364061
transform 1 0 17848 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_191
timestamp 1586364061
transform 1 0 18676 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18952 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18952 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20700 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_205
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_205
timestamp 1586364061
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_209
timestamp 1586364061
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22264 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_222
timestamp 1586364061
transform 1 0 21528 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_226
timestamp 1586364061
transform 1 0 21896 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_237
timestamp 1586364061
transform 1 0 22908 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_233
timestamp 1586364061
transform 1 0 22540 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23092 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_248
timestamp 1586364061
transform 1 0 23920 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_241
timestamp 1586364061
transform 1 0 23276 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_conb_1  _127_
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_241
timestamp 1586364061
transform 1 0 23276 0 -1 16864
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_253
timestamp 1586364061
transform 1 0 24380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_265
timestamp 1586364061
transform 1 0 25484 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_252
timestamp 1586364061
transform 1 0 24288 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_273
timestamp 1586364061
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_74
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11684 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_28_124
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_128
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_149
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_167
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 1142 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_179
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_189
timestamp 1586364061
transform 1 0 18492 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_212
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_1  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_225
timestamp 1586364061
transform 1 0 21804 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22540 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_242
timestamp 1586364061
transform 1 0 23368 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _162_
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_254
timestamp 1586364061
transform 1 0 24472 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_259
timestamp 1586364061
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_73
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_79
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_93
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 12604 0 1 17952
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_134
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_138
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_151
timestamp 1586364061
transform 1 0 14996 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_157
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_168
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_172
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_176
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_182
timestamp 1586364061
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_202
timestamp 1586364061
transform 1 0 19688 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_206
timestamp 1586364061
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_219
timestamp 1586364061
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_223
timestamp 1586364061
transform 1 0 21620 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_230
timestamp 1586364061
transform 1 0 22264 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_234
timestamp 1586364061
transform 1 0 22632 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_242
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use scs8hd_conb_1  _126_
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_113
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_121
timestamp 1586364061
transform 1 0 12236 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_133
timestamp 1586364061
transform 1 0 13340 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_164
timestamp 1586364061
transform 1 0 16192 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_176
timestamp 1586364061
transform 1 0 17296 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_188
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_200
timestamp 1586364061
transform 1 0 19504 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_30_212
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21436 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_236
timestamp 1586364061
transform 1 0 22816 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_248
timestamp 1586364061
transform 1 0 23920 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_260
timestamp 1586364061
transform 1 0 25024 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_272
timestamp 1586364061
transform 1 0 26128 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_109
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_113
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_117
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_120
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_127
timestamp 1586364061
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_131
timestamp 1586364061
transform 1 0 13156 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_158
timestamp 1586364061
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_162
timestamp 1586364061
transform 1 0 16008 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_174
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_182
timestamp 1586364061
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11960 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_121
timestamp 1586364061
transform 1 0 12236 0 -1 20128
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 13800 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_133
timestamp 1586364061
transform 1 0 13340 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_137
timestamp 1586364061
transform 1 0 13708 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_140
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_258
timestamp 1586364061
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_270
timestamp 1586364061
transform 1 0 25944 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_19
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_43
timestamp 1586364061
transform 1 0 5060 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_37_55
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_258
timestamp 1586364061
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_262
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_274
timestamp 1586364061
transform 1 0 26312 0 1 22304
box -38 -48 314 592
use scs8hd_buf_2  _156_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_37
timestamp 1586364061
transform 1 0 4508 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_41
timestamp 1586364061
transform 1 0 4876 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _136_
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_66
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_70
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_82
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_94
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_106
timestamp 1586364061
transform 1 0 10856 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _148_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _145_
timestamp 1586364061
transform 1 0 14076 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 12972 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_127
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_131
timestamp 1586364061
transform 1 0 13156 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_139
timestamp 1586364061
transform 1 0 13892 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_145
timestamp 1586364061
transform 1 0 14444 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_149
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _160_
timestamp 1586364061
transform 1 0 15916 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 16468 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_165
timestamp 1586364061
transform 1 0 16284 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_169
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_177
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_181
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _159_
timestamp 1586364061
transform 1 0 17572 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_192
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 18952 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _157_
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_195
timestamp 1586364061
transform 1 0 19044 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_183
timestamp 1586364061
transform 1 0 17940 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_40_207
timestamp 1586364061
transform 1 0 20148 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_213
timestamp 1586364061
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_228
timestamp 1586364061
transform 1 0 22080 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_240
timestamp 1586364061
transform 1 0 23184 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_236
timestamp 1586364061
transform 1 0 22816 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23276 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23276 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_244
timestamp 1586364061
transform 1 0 23552 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_258
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_262
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_256
timestamp 1586364061
transform 1 0 24656 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_40_268
timestamp 1586364061
transform 1 0 25760 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_274
timestamp 1586364061
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 662 27520 718 28000 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 824 480 944 6 address[1]
port 1 nsew default input
rlabel metal3 s 27520 688 28000 808 6 address[2]
port 2 nsew default input
rlabel metal2 s 2318 0 2374 480 6 address[3]
port 3 nsew default input
rlabel metal3 s 27520 2184 28000 2304 6 address[4]
port 4 nsew default input
rlabel metal2 s 2042 27520 2098 28000 6 address[5]
port 5 nsew default input
rlabel metal2 s 3422 27520 3478 28000 6 address[6]
port 6 nsew default input
rlabel metal3 s 0 2456 480 2576 6 chanx_left_in[0]
port 7 nsew default input
rlabel metal2 s 3330 0 3386 480 6 chanx_left_in[1]
port 8 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[2]
port 9 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[3]
port 10 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 chanx_left_in[4]
port 11 nsew default input
rlabel metal2 s 4250 0 4306 480 6 chanx_left_in[5]
port 12 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chanx_left_in[6]
port 13 nsew default input
rlabel metal2 s 4802 27520 4858 28000 6 chanx_left_in[7]
port 14 nsew default input
rlabel metal3 s 27520 5312 28000 5432 6 chanx_left_in[8]
port 15 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chanx_left_out[0]
port 16 nsew default tristate
rlabel metal3 s 0 7760 480 7880 6 chanx_left_out[1]
port 17 nsew default tristate
rlabel metal2 s 7194 0 7250 480 6 chanx_left_out[2]
port 18 nsew default tristate
rlabel metal2 s 8114 0 8170 480 6 chanx_left_out[3]
port 19 nsew default tristate
rlabel metal3 s 27520 6808 28000 6928 6 chanx_left_out[4]
port 20 nsew default tristate
rlabel metal2 s 9126 0 9182 480 6 chanx_left_out[5]
port 21 nsew default tristate
rlabel metal3 s 27520 8440 28000 8560 6 chanx_left_out[6]
port 22 nsew default tristate
rlabel metal3 s 27520 9936 28000 10056 6 chanx_left_out[7]
port 23 nsew default tristate
rlabel metal2 s 6182 27520 6238 28000 6 chanx_left_out[8]
port 24 nsew default tristate
rlabel metal3 s 0 9528 480 9648 6 chanx_right_in[0]
port 25 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chanx_right_in[1]
port 26 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chanx_right_in[2]
port 27 nsew default input
rlabel metal2 s 11058 0 11114 480 6 chanx_right_in[3]
port 28 nsew default input
rlabel metal2 s 9034 27520 9090 28000 6 chanx_right_in[4]
port 29 nsew default input
rlabel metal2 s 10414 27520 10470 28000 6 chanx_right_in[5]
port 30 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chanx_right_in[6]
port 31 nsew default input
rlabel metal2 s 11794 27520 11850 28000 6 chanx_right_in[7]
port 32 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_right_in[8]
port 33 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_right_out[0]
port 34 nsew default tristate
rlabel metal3 s 27520 11568 28000 11688 6 chanx_right_out[1]
port 35 nsew default tristate
rlabel metal2 s 12990 0 13046 480 6 chanx_right_out[2]
port 36 nsew default tristate
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_out[3]
port 37 nsew default tristate
rlabel metal2 s 13910 0 13966 480 6 chanx_right_out[4]
port 38 nsew default tristate
rlabel metal2 s 13174 27520 13230 28000 6 chanx_right_out[5]
port 39 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_right_out[6]
port 40 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_right_out[7]
port 41 nsew default tristate
rlabel metal2 s 14646 27520 14702 28000 6 chanx_right_out[8]
port 42 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chany_top_in[0]
port 43 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chany_top_in[1]
port 44 nsew default input
rlabel metal2 s 16026 27520 16082 28000 6 chany_top_in[2]
port 45 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_top_in[3]
port 46 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chany_top_in[4]
port 47 nsew default input
rlabel metal2 s 15842 0 15898 480 6 chany_top_in[5]
port 48 nsew default input
rlabel metal3 s 27520 14696 28000 14816 6 chany_top_in[6]
port 49 nsew default input
rlabel metal3 s 27520 16192 28000 16312 6 chany_top_in[7]
port 50 nsew default input
rlabel metal3 s 27520 17688 28000 17808 6 chany_top_in[8]
port 51 nsew default input
rlabel metal3 s 27520 19320 28000 19440 6 chany_top_out[0]
port 52 nsew default tristate
rlabel metal2 s 16854 0 16910 480 6 chany_top_out[1]
port 53 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[2]
port 54 nsew default tristate
rlabel metal2 s 18786 27520 18842 28000 6 chany_top_out[3]
port 55 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_top_out[4]
port 56 nsew default tristate
rlabel metal2 s 20166 27520 20222 28000 6 chany_top_out[5]
port 57 nsew default tristate
rlabel metal3 s 0 23536 480 23656 6 chany_top_out[6]
port 58 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 chany_top_out[7]
port 59 nsew default tristate
rlabel metal2 s 19706 0 19762 480 6 chany_top_out[8]
port 60 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 data_in
port 61 nsew default input
rlabel metal2 s 478 0 534 480 6 enable
port 62 nsew default input
rlabel metal2 s 20718 0 20774 480 6 left_bottom_grid_pin_11_
port 63 nsew default input
rlabel metal2 s 23018 27520 23074 28000 6 left_bottom_grid_pin_13_
port 64 nsew default input
rlabel metal2 s 21638 0 21694 480 6 left_bottom_grid_pin_15_
port 65 nsew default input
rlabel metal3 s 27520 20816 28000 20936 6 left_bottom_grid_pin_1_
port 66 nsew default input
rlabel metal3 s 27520 22448 28000 22568 6 left_bottom_grid_pin_3_
port 67 nsew default input
rlabel metal3 s 27520 23944 28000 24064 6 left_bottom_grid_pin_5_
port 68 nsew default input
rlabel metal2 s 21638 27520 21694 28000 6 left_bottom_grid_pin_7_
port 69 nsew default input
rlabel metal3 s 0 25304 480 25424 6 left_bottom_grid_pin_9_
port 70 nsew default input
rlabel metal2 s 22650 0 22706 480 6 left_top_grid_pin_10_
port 71 nsew default input
rlabel metal2 s 26514 0 26570 480 6 right_bottom_grid_pin_11_
port 72 nsew default input
rlabel metal2 s 27434 0 27490 480 6 right_bottom_grid_pin_13_
port 73 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 right_bottom_grid_pin_15_
port 74 nsew default input
rlabel metal2 s 23570 0 23626 480 6 right_bottom_grid_pin_1_
port 75 nsew default input
rlabel metal2 s 24582 0 24638 480 6 right_bottom_grid_pin_3_
port 76 nsew default input
rlabel metal3 s 27520 25576 28000 25696 6 right_bottom_grid_pin_5_
port 77 nsew default input
rlabel metal2 s 25502 0 25558 480 6 right_bottom_grid_pin_7_
port 78 nsew default input
rlabel metal2 s 24398 27520 24454 28000 6 right_bottom_grid_pin_9_
port 79 nsew default input
rlabel metal2 s 25778 27520 25834 28000 6 right_top_grid_pin_10_
port 80 nsew default input
rlabel metal2 s 27158 27520 27214 28000 6 top_left_grid_pin_13_
port 81 nsew default input
rlabel metal3 s 0 27072 480 27192 6 top_right_grid_pin_11_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
